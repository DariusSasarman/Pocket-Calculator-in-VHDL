library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity Eight_bit_twos_complement_to_seven_seg_display is
    Port ( number : in STD_LOGIC_VECTOR (7 downto 0);
           display : out STD_LOGIC_VECTOR (31 downto 0));
end Eight_bit_twos_complement_to_seven_seg_display;

architecture Behavioral of Eight_bit_twos_complement_to_seven_seg_display is
type rom_type is array (integer range -128 to 127) of std_logic_vector(31 downto 0);
constant ROM : rom_type := (
  -128 => x"BFF9A480",
  -127 => x"BFF9A4F8",
  -126 => x"BFF9A482",
  -125 => x"BFF9A492",
  -124 => x"BFF9A499",
  -123 => x"BFF9A4B0",
  -122 => x"BFF9A4A4",
  -121 => x"BFF9A4F9",
  -120 => x"BFF9A4C0",
  -119 => x"BFF9F990",
  -118 => x"BFF9F980",
  -117 => x"BFF9F9F8",
  -116 => x"BFF9F982",
  -115 => x"BFF9F992",
  -114 => x"BFF9F999",
  -113 => x"BFF9F9B0",
  -112 => x"BFF9F9A4",
  -111 => x"BFF9F9F9",
  -110 => x"BFF9F9C0",
  -109 => x"BFF9C090",
  -108 => x"BFF9C080",
  -107 => x"BFF9C0F8",
  -106 => x"BFF9C082",
  -105 => x"BFF9C092",
  -104 => x"BFF9C099",
  -103 => x"BFF9C0B0",
  -102 => x"BFF9C0A4",
  -101 => x"BFF9C0F9",
  -100 => x"BFF9C0C0",
   -99 => x"C0BF9090",
   -98 => x"C0BF9080",
   -97 => x"C0BF90F8",
   -96 => x"C0BF9082",
   -95 => x"C0BF9092",
   -94 => x"C0BF9099",
   -93 => x"C0BF90B0",
   -92 => x"C0BF90A4",
   -91 => x"C0BF90F9",
   -90 => x"C0BF90C0",
   -89 => x"C0BF8090",
   -88 => x"C0BF8080",
   -87 => x"C0BF80F8",
   -86 => x"C0BF8082",
   -85 => x"C0BF8092",
   -84 => x"C0BF8099",
   -83 => x"C0BF80B0",
   -82 => x"C0BF80A4",
   -81 => x"C0BF80F9",
   -80 => x"C0BF80C0",
   -79 => x"C0BFF890",
   -78 => x"C0BFF880",
   -77 => x"C0BFF8F8",
   -76 => x"C0BFF882",
   -75 => x"C0BFF892",
   -74 => x"C0BFF899",
   -73 => x"C0BFF8B0",
   -72 => x"C0BFF8A4",
   -71 => x"C0BFF8F9",
   -70 => x"C0BFF8C0",
   -69 => x"C0BF8290",
   -68 => x"C0BF8280",
   -67 => x"C0BF82F8",
   -66 => x"C0BF8282",
   -65 => x"C0BF8292",
   -64 => x"C0BF8299",
   -63 => x"C0BF82B0",
   -62 => x"C0BF82A4",
   -61 => x"C0BF82F9",
   -60 => x"C0BF82C0",
   -59 => x"C0BF9290",
   -58 => x"C0BF9280",
   -57 => x"C0BF92F8",
   -56 => x"C0BF9282",
   -55 => x"C0BF9292",
   -54 => x"C0BF9299",
   -53 => x"C0BF92B0",
   -52 => x"C0BF92A4",
   -51 => x"C0BF92F9",
   -50 => x"C0BF92C0",
   -49 => x"C0BF9990",
   -48 => x"C0BF9980",
   -47 => x"C0BF99F8",
   -46 => x"C0BF9982",
   -45 => x"C0BF9992",
   -44 => x"C0BF9999",
   -43 => x"C0BF99B0",
   -42 => x"C0BF99A4",
   -41 => x"C0BF99F9",
   -40 => x"C0BF99C0",
   -39 => x"C0BFB090",
   -38 => x"C0BFB080",
   -37 => x"C0BFB0F8",
   -36 => x"C0BFB082",
   -35 => x"C0BFB092",
   -34 => x"C0BFB099",
   -33 => x"C0BFB0B0",
   -32 => x"C0BFB0A4",
   -31 => x"C0BFB0F9",
   -30 => x"C0BFB0C0",
   -29 => x"C0BFA490",
   -28 => x"C0BFA480",
   -27 => x"C0BFA4F8",
   -26 => x"C0BFA482",
   -25 => x"C0BFA492",
   -24 => x"C0BFA499",
   -23 => x"C0BFA4B0",
   -22 => x"C0BFA4A4",
   -21 => x"C0BFA4F9",
   -20 => x"C0BFA4C0",
   -19 => x"C0BFF990",
   -18 => x"C0BFF980",
   -17 => x"C0BFF9F8",
   -16 => x"C0BFF982",
   -15 => x"C0BFF992",
   -14 => x"C0BFF999",
   -13 => x"C0BFF9B0",
   -12 => x"C0BFF9A4",
   -11 => x"C0BFF9F9",
   -10 => x"C0BFF9C0",
    -9 => x"C0C0BF90",
    -8 => x"C0C0BF80",
    -7 => x"C0C0BFF8",
    -6 => x"C0C0BF82",
    -5 => x"C0C0BF92",
    -4 => x"C0C0BF99",
    -3 => x"C0C0BFB0",
    -2 => x"C0C0BFA4",
    -1 => x"C0C0BFF9",
     0 => x"C0C0C0C0",
     1 => x"C0C0C0F9",
     2 => x"C0C0C0A4",
     3 => x"C0C0C0B0",
     4 => x"C0C0C099",
     5 => x"C0C0C092",
     6 => x"C0C0C082",
     7 => x"C0C0C0F8",
     8 => x"C0C0C080",
     9 => x"C0C0C090",
    10 => x"C0C0F9C0",
    11 => x"C0C0F9F9",
    12 => x"C0C0F9A4",
    13 => x"C0C0F9B0",
    14 => x"C0C0F999",
    15 => x"C0C0F992",
    16 => x"C0C0F982",
    17 => x"C0C0F9F8",
    18 => x"C0C0F980",
    19 => x"C0C0F990",
    20 => x"C0C0A4C0",
    21 => x"C0C0A4F9",
    22 => x"C0C0A4A4",
    23 => x"C0C0A4B0",
    24 => x"C0C0A499",
    25 => x"C0C0A492",
    26 => x"C0C0A482",
    27 => x"C0C0A4F8",
    28 => x"C0C0A480",
    29 => x"C0C0A490",
    30 => x"C0C0B0C0",
    31 => x"C0C0B0F9",
    32 => x"C0C0B0A4",
    33 => x"C0C0B0B0",
    34 => x"C0C0B099",
    35 => x"C0C0B092",
    36 => x"C0C0B082",
    37 => x"C0C0B0F8",
    38 => x"C0C0B080",
    39 => x"C0C0B090",
    40 => x"C0C099C0",
    41 => x"C0C099F9",
    42 => x"C0C099A4",
    43 => x"C0C099B0",
    44 => x"C0C09999",
    45 => x"C0C09992",
    46 => x"C0C09982",
    47 => x"C0C099F8",
    48 => x"C0C09980",
    49 => x"C0C09990",
    50 => x"C0C092C0",
    51 => x"C0C092F9",
    52 => x"C0C092A4",
    53 => x"C0C092B0",
    54 => x"C0C09299",
    55 => x"C0C09292",
    56 => x"C0C09282",
    57 => x"C0C092F8",
    58 => x"C0C09280",
    59 => x"C0C09290",
    60 => x"C0C082C0",
    61 => x"C0C082F9",
    62 => x"C0C082A4",
    63 => x"C0C082B0",
    64 => x"C0C08299",
    65 => x"C0C08292",
    66 => x"C0C08282",
    67 => x"C0C082F8",
    68 => x"C0C08280",
    69 => x"C0C08290",
    70 => x"C0C0F8C0",
    71 => x"C0C0F8F9",
    72 => x"C0C0F8A4",
    73 => x"C0C0F8B0",
    74 => x"C0C0F899",
    75 => x"C0C0F892",
    76 => x"C0C0F882",
    77 => x"C0C0F8F8",
    78 => x"C0C0F880",
    79 => x"C0C0F890",
    80 => x"C0C080C0",
    81 => x"C0C080F9",
    82 => x"C0C080A4",
    83 => x"C0C080B0",
    84 => x"C0C08099",
    85 => x"C0C08092",
    86 => x"C0C08082",
    87 => x"C0C080F8",
    88 => x"C0C08080",
    89 => x"C0C08090",
    90 => x"C0C090C0",
    91 => x"C0C090F9",
    92 => x"C0C090A4",
    93 => x"C0C090B0",
    94 => x"C0C09099",
    95 => x"C0C09092",
    96 => x"C0C09082",
    97 => x"C0C090F8",
    98 => x"C0C09080",
    99 => x"C0C09090",
   100 => x"C0F9C0C0",
   101 => x"C0F9C0F9",
   102 => x"C0F9C0A4",
   103 => x"C0F9C0B0",
   104 => x"C0F9C099",
   105 => x"C0F9C092",
   106 => x"C0F9C082",
   107 => x"C0F9C0F8",
   108 => x"C0F9C080",
   109 => x"C0F9C090",
   110 => x"C0F9F9C0",
   111 => x"C0F9F9F9",
   112 => x"C0F9F9A4",
   113 => x"C0F9F9B0",
   114 => x"C0F9F999",
   115 => x"C0F9F992",
   116 => x"C0F9F982",
   117 => x"C0F9F9F8",
   118 => x"C0F9F980",
   119 => x"C0F9F990",
   120 => x"C0F9A4C0",
   121 => x"C0F9A4F9",
   122 => x"C0F9A4A4",
   123 => x"C0F9A4B0",
   124 => x"C0F9A499",
   125 => x"C0F9A492",
   126 => x"C0F9A482",
   127 => x"C0F9A4F8"
);
    
begin

display <= ROM(to_integer(signed(number)));

end Behavioral;
