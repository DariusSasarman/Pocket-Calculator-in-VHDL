library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity subtraction_output_processor is
   Port(
       inp : in std_logic_vector ( 8 downto 0);
       outp: out std_logic_vector( 63 downto 0)
       );
end subtraction_output_processor;

architecture Behavioral of subtraction_output_processor is

type rom_type is array (integer range -256 to 255) of std_logic_vector(31 downto 0);
constant ROM : rom_type := (
  -256 => x"BFA49282",
  -255 => x"BFA49292",
  -254 => x"BFA49299",
  -253 => x"BFA492B0",
  -252 => x"BFA492A4",
  -251 => x"BFA492F9",
  -250 => x"BFA492C0",
  -249 => x"BFA49990",
  -248 => x"BFA49980",
  -247 => x"BFA499F8",
  -246 => x"BFA49982",
  -245 => x"BFA49992",
  -244 => x"BFA49999",
  -243 => x"BFA499B0",
  -242 => x"BFA499A4",
  -241 => x"BFA499F9",
  -240 => x"BFA499C0",
  -239 => x"BFA4B090",
  -238 => x"BFA4B080",
  -237 => x"BFA4B0F8",
  -236 => x"BFA4B082",
  -235 => x"BFA4B092",
  -234 => x"BFA4B099",
  -233 => x"BFA4B0B0",
  -232 => x"BFA4B0A4",
  -231 => x"BFA4B0F9",
  -230 => x"BFA4B0C0",
  -229 => x"BFA4A490",
  -228 => x"BFA4A480",
  -227 => x"BFA4A4F8",
  -226 => x"BFA4A482",
  -225 => x"BFA4A492",
  -224 => x"BFA4A499",
  -223 => x"BFA4A4B0",
  -222 => x"BFA4A4A4",
  -221 => x"BFA4A4F9",
  -220 => x"BFA4A4C0",
  -219 => x"BFA4F990",
  -218 => x"BFA4F980",
  -217 => x"BFA4F9F8",
  -216 => x"BFA4F982",
  -215 => x"BFA4F992",
  -214 => x"BFA4F999",
  -213 => x"BFA4F9B0",
  -212 => x"BFA4F9A4",
  -211 => x"BFA4F9F9",
  -210 => x"BFA4F9C0",
  -209 => x"BFA4C090",
  -208 => x"BFA4C080",
  -207 => x"BFA4C0F8",
  -206 => x"BFA4C082",
  -205 => x"BFA4C092",
  -204 => x"BFA4C099",
  -203 => x"BFA4C0B0",
  -202 => x"BFA4C0A4",
  -201 => x"BFA4C0F9",
  -200 => x"BFA4C0C0",
  -199 => x"BFF99090",
  -198 => x"BFF99080",
  -197 => x"BFF990F8",
  -196 => x"BFF99082",
  -195 => x"BFF99092",
  -194 => x"BFF99099",
  -193 => x"BFF990B0",
  -192 => x"BFF990A4",
  -191 => x"BFF990F9",
  -190 => x"BFF990C0",
  -189 => x"BFF98090",
  -188 => x"BFF98080",
  -187 => x"BFF980F8",
  -186 => x"BFF98082",
  -185 => x"BFF98092",
  -184 => x"BFF98099",
  -183 => x"BFF980B0",
  -182 => x"BFF980A4",
  -181 => x"BFF980F9",
  -180 => x"BFF980C0",
  -179 => x"BFF9F890",
  -178 => x"BFF9F880",
  -177 => x"BFF9F8F8",
  -176 => x"BFF9F882",
  -175 => x"BFF9F892",
  -174 => x"BFF9F899",
  -173 => x"BFF9F8B0",
  -172 => x"BFF9F8A4",
  -171 => x"BFF9F8F9",
  -170 => x"BFF9F8C0",
  -169 => x"BFF98290",
  -168 => x"BFF98280",
  -167 => x"BFF982F8",
  -166 => x"BFF98282",
  -165 => x"BFF98292",
  -164 => x"BFF98299",
  -163 => x"BFF982B0",
  -162 => x"BFF982A4",
  -161 => x"BFF982F9",
  -160 => x"BFF982C0",
  -159 => x"BFF99290",
  -158 => x"BFF99280",
  -157 => x"BFF992F8",
  -156 => x"BFF99282",
  -155 => x"BFF99292",
  -154 => x"BFF99299",
  -153 => x"BFF992B0",
  -152 => x"BFF992A4",
  -151 => x"BFF992F9",
  -150 => x"BFF992C0",
  -149 => x"BFF99990",
  -148 => x"BFF99980",
  -147 => x"BFF999F8",
  -146 => x"BFF99982",
  -145 => x"BFF99992",
  -144 => x"BFF99999",
  -143 => x"BFF999B0",
  -142 => x"BFF999A4",
  -141 => x"BFF999F9",
  -140 => x"BFF999C0",
  -139 => x"BFF9B090",
  -138 => x"BFF9B080",
  -137 => x"BFF9B0F8",
  -136 => x"BFF9B082",
  -135 => x"BFF9B092",
  -134 => x"BFF9B099",
  -133 => x"BFF9B0B0",
  -132 => x"BFF9B0A4",
  -131 => x"BFF9B0F9",
  -130 => x"BFF9B0C0",
  -129 => x"BFF9A490",
  -128 => x"BFF9A480",
  -127 => x"BFF9A4F8",
  -126 => x"BFF9A482",
  -125 => x"BFF9A492",
  -124 => x"BFF9A499",
  -123 => x"BFF9A4B0",
  -122 => x"BFF9A4A4",
  -121 => x"BFF9A4F9",
  -120 => x"BFF9A4C0",
  -119 => x"BFF9F990",
  -118 => x"BFF9F980",
  -117 => x"BFF9F9F8",
  -116 => x"BFF9F982",
  -115 => x"BFF9F992",
  -114 => x"BFF9F999",
  -113 => x"BFF9F9B0",
  -112 => x"BFF9F9A4",
  -111 => x"BFF9F9F9",
  -110 => x"BFF9F9C0",
  -109 => x"BFF9C090",
  -108 => x"BFF9C080",
  -107 => x"BFF9C0F8",
  -106 => x"BFF9C082",
  -105 => x"BFF9C092",
  -104 => x"BFF9C099",
  -103 => x"BFF9C0B0",
  -102 => x"BFF9C0A4",
  -101 => x"BFF9C0F9",
  -100 => x"BFF9C0C0",
   -99 => x"C0BF9090",
   -98 => x"C0BF9080",
   -97 => x"C0BF90F8",
   -96 => x"C0BF9082",
   -95 => x"C0BF9092",
   -94 => x"C0BF9099",
   -93 => x"C0BF90B0",
   -92 => x"C0BF90A4",
   -91 => x"C0BF90F9",
   -90 => x"C0BF90C0",
   -89 => x"C0BF8090",
   -88 => x"C0BF8080",
   -87 => x"C0BF80F8",
   -86 => x"C0BF8082",
   -85 => x"C0BF8092",
   -84 => x"C0BF8099",
   -83 => x"C0BF80B0",
   -82 => x"C0BF80A4",
   -81 => x"C0BF80F9",
   -80 => x"C0BF80C0",
   -79 => x"C0BFF890",
   -78 => x"C0BFF880",
   -77 => x"C0BFF8F8",
   -76 => x"C0BFF882",
   -75 => x"C0BFF892",
   -74 => x"C0BFF899",
   -73 => x"C0BFF8B0",
   -72 => x"C0BFF8A4",
   -71 => x"C0BFF8F9",
   -70 => x"C0BFF8C0",
   -69 => x"C0BF8290",
   -68 => x"C0BF8280",
   -67 => x"C0BF82F8",
   -66 => x"C0BF8282",
   -65 => x"C0BF8292",
   -64 => x"C0BF8299",
   -63 => x"C0BF82B0",
   -62 => x"C0BF82A4",
   -61 => x"C0BF82F9",
   -60 => x"C0BF82C0",
   -59 => x"C0BF9290",
   -58 => x"C0BF9280",
   -57 => x"C0BF92F8",
   -56 => x"C0BF9282",
   -55 => x"C0BF9292",
   -54 => x"C0BF9299",
   -53 => x"C0BF92B0",
   -52 => x"C0BF92A4",
   -51 => x"C0BF92F9",
   -50 => x"C0BF92C0",
   -49 => x"C0BF9990",
   -48 => x"C0BF9980",
   -47 => x"C0BF99F8",
   -46 => x"C0BF9982",
   -45 => x"C0BF9992",
   -44 => x"C0BF9999",
   -43 => x"C0BF99B0",
   -42 => x"C0BF99A4",
   -41 => x"C0BF99F9",
   -40 => x"C0BF99C0",
   -39 => x"C0BFB090",
   -38 => x"C0BFB080",
   -37 => x"C0BFB0F8",
   -36 => x"C0BFB082",
   -35 => x"C0BFB092",
   -34 => x"C0BFB099",
   -33 => x"C0BFB0B0",
   -32 => x"C0BFB0A4",
   -31 => x"C0BFB0F9",
   -30 => x"C0BFB0C0",
   -29 => x"C0BFA490",
   -28 => x"C0BFA480",
   -27 => x"C0BFA4F8",
   -26 => x"C0BFA482",
   -25 => x"C0BFA492",
   -24 => x"C0BFA499",
   -23 => x"C0BFA4B0",
   -22 => x"C0BFA4A4",
   -21 => x"C0BFA4F9",
   -20 => x"C0BFA4C0",
   -19 => x"C0BFF990",
   -18 => x"C0BFF980",
   -17 => x"C0BFF9F8",
   -16 => x"C0BFF982",
   -15 => x"C0BFF992",
   -14 => x"C0BFF999",
   -13 => x"C0BFF9B0",
   -12 => x"C0BFF9A4",
   -11 => x"C0BFF9F9",
   -10 => x"C0BFF9C0",
    -9 => x"C0C0BF90",
    -8 => x"C0C0BF80",
    -7 => x"C0C0BFF8",
    -6 => x"C0C0BF82",
    -5 => x"C0C0BF92",
    -4 => x"C0C0BF99",
    -3 => x"C0C0BFB0",
    -2 => x"C0C0BFA4",
    -1 => x"C0C0BFF9",
     0 => x"C0C0C0C0",
     1 => x"C0C0C0F9",
     2 => x"C0C0C0A4",
     3 => x"C0C0C0B0",
     4 => x"C0C0C099",
     5 => x"C0C0C092",
     6 => x"C0C0C082",
     7 => x"C0C0C0F8",
     8 => x"C0C0C080",
     9 => x"C0C0C090",
    10 => x"C0C0F9C0",
    11 => x"C0C0F9F9",
    12 => x"C0C0F9A4",
    13 => x"C0C0F9B0",
    14 => x"C0C0F999",
    15 => x"C0C0F992",
    16 => x"C0C0F982",
    17 => x"C0C0F9F8",
    18 => x"C0C0F980",
    19 => x"C0C0F990",
    20 => x"C0C0A4C0",
    21 => x"C0C0A4F9",
    22 => x"C0C0A4A4",
    23 => x"C0C0A4B0",
    24 => x"C0C0A499",
    25 => x"C0C0A492",
    26 => x"C0C0A482",
    27 => x"C0C0A4F8",
    28 => x"C0C0A480",
    29 => x"C0C0A490",
    30 => x"C0C0B0C0",
    31 => x"C0C0B0F9",
    32 => x"C0C0B0A4",
    33 => x"C0C0B0B0",
    34 => x"C0C0B099",
    35 => x"C0C0B092",
    36 => x"C0C0B082",
    37 => x"C0C0B0F8",
    38 => x"C0C0B080",
    39 => x"C0C0B090",
    40 => x"C0C099C0",
    41 => x"C0C099F9",
    42 => x"C0C099A4",
    43 => x"C0C099B0",
    44 => x"C0C09999",
    45 => x"C0C09992",
    46 => x"C0C09982",
    47 => x"C0C099F8",
    48 => x"C0C09980",
    49 => x"C0C09990",
    50 => x"C0C092C0",
    51 => x"C0C092F9",
    52 => x"C0C092A4",
    53 => x"C0C092B0",
    54 => x"C0C09299",
    55 => x"C0C09292",
    56 => x"C0C09282",
    57 => x"C0C092F8",
    58 => x"C0C09280",
    59 => x"C0C09290",
    60 => x"C0C082C0",
    61 => x"C0C082F9",
    62 => x"C0C082A4",
    63 => x"C0C082B0",
    64 => x"C0C08299",
    65 => x"C0C08292",
    66 => x"C0C08282",
    67 => x"C0C082F8",
    68 => x"C0C08280",
    69 => x"C0C08290",
    70 => x"C0C0F8C0",
    71 => x"C0C0F8F9",
    72 => x"C0C0F8A4",
    73 => x"C0C0F8B0",
    74 => x"C0C0F899",
    75 => x"C0C0F892",
    76 => x"C0C0F882",
    77 => x"C0C0F8F8",
    78 => x"C0C0F880",
    79 => x"C0C0F890",
    80 => x"C0C080C0",
    81 => x"C0C080F9",
    82 => x"C0C080A4",
    83 => x"C0C080B0",
    84 => x"C0C08099",
    85 => x"C0C08092",
    86 => x"C0C08082",
    87 => x"C0C080F8",
    88 => x"C0C08080",
    89 => x"C0C08090",
    90 => x"C0C090C0",
    91 => x"C0C090F9",
    92 => x"C0C090A4",
    93 => x"C0C090B0",
    94 => x"C0C09099",
    95 => x"C0C09092",
    96 => x"C0C09082",
    97 => x"C0C090F8",
    98 => x"C0C09080",
    99 => x"C0C09090",
   100 => x"C0F9C0C0",
   101 => x"C0F9C0F9",
   102 => x"C0F9C0A4",
   103 => x"C0F9C0B0",
   104 => x"C0F9C099",
   105 => x"C0F9C092",
   106 => x"C0F9C082",
   107 => x"C0F9C0F8",
   108 => x"C0F9C080",
   109 => x"C0F9C090",
   110 => x"C0F9F9C0",
   111 => x"C0F9F9F9",
   112 => x"C0F9F9A4",
   113 => x"C0F9F9B0",
   114 => x"C0F9F999",
   115 => x"C0F9F992",
   116 => x"C0F9F982",
   117 => x"C0F9F9F8",
   118 => x"C0F9F980",
   119 => x"C0F9F990",
   120 => x"C0F9A4C0",
   121 => x"C0F9A4F9",
   122 => x"C0F9A4A4",
   123 => x"C0F9A4B0",
   124 => x"C0F9A499",
   125 => x"C0F9A492",
   126 => x"C0F9A482",
   127 => x"C0F9A4F8",
   128 => x"C0F9A480",
   129 => x"C0F9A490",
   130 => x"C0F9B0C0",
   131 => x"C0F9B0F9",
   132 => x"C0F9B0A4",
   133 => x"C0F9B0B0",
   134 => x"C0F9B099",
   135 => x"C0F9B092",
   136 => x"C0F9B082",
   137 => x"C0F9B0F8",
   138 => x"C0F9B080",
   139 => x"C0F9B090",
   140 => x"C0F999C0",
   141 => x"C0F999F9",
   142 => x"C0F999A4",
   143 => x"C0F999B0",
   144 => x"C0F99999",
   145 => x"C0F99992",
   146 => x"C0F99982",
   147 => x"C0F999F8",
   148 => x"C0F99980",
   149 => x"C0F99990",
   150 => x"C0F992C0",
   151 => x"C0F992F9",
   152 => x"C0F992A4",
   153 => x"C0F992B0",
   154 => x"C0F99299",
   155 => x"C0F99292",
   156 => x"C0F99282",
   157 => x"C0F992F8",
   158 => x"C0F99280",
   159 => x"C0F99290",
   160 => x"C0F982C0",
   161 => x"C0F982F9",
   162 => x"C0F982A4",
   163 => x"C0F982B0",
   164 => x"C0F98299",
   165 => x"C0F98292",
   166 => x"C0F98282",
   167 => x"C0F982F8",
   168 => x"C0F98280",
   169 => x"C0F98290",
   170 => x"C0F9F8C0",
   171 => x"C0F9F8F9",
   172 => x"C0F9F8A4",
   173 => x"C0F9F8B0",
   174 => x"C0F9F899",
   175 => x"C0F9F892",
   176 => x"C0F9F882",
   177 => x"C0F9F8F8",
   178 => x"C0F9F880",
   179 => x"C0F9F890",
   180 => x"C0F980C0",
   181 => x"C0F980F9",
   182 => x"C0F980A4",
   183 => x"C0F980B0",
   184 => x"C0F98099",
   185 => x"C0F98092",
   186 => x"C0F98082",
   187 => x"C0F980F8",
   188 => x"C0F98080",
   189 => x"C0F98090",
   190 => x"C0F990C0",
   191 => x"C0F990F9",
   192 => x"C0F990A4",
   193 => x"C0F990B0",
   194 => x"C0F99099",
   195 => x"C0F99092",
   196 => x"C0F99082",
   197 => x"C0F990F8",
   198 => x"C0F99080",
   199 => x"C0F99090",
   200 => x"C0A4C0C0",
   201 => x"C0A4C0F9",
   202 => x"C0A4C0A4",
   203 => x"C0A4C0B0",
   204 => x"C0A4C099",
   205 => x"C0A4C092",
   206 => x"C0A4C082",
   207 => x"C0A4C0F8",
   208 => x"C0A4C080",
   209 => x"C0A4C090",
   210 => x"C0A4F9C0",
   211 => x"C0A4F9F9",
   212 => x"C0A4F9A4",
   213 => x"C0A4F9B0",
   214 => x"C0A4F999",
   215 => x"C0A4F992",
   216 => x"C0A4F982",
   217 => x"C0A4F9F8",
   218 => x"C0A4F980",
   219 => x"C0A4F990",
   220 => x"C0A4A4C0",
   221 => x"C0A4A4F9",
   222 => x"C0A4A4A4",
   223 => x"C0A4A4B0",
   224 => x"C0A4A499",
   225 => x"C0A4A492",
   226 => x"C0A4A482",
   227 => x"C0A4A4F8",
   228 => x"C0A4A480",
   229 => x"C0A4A490",
   230 => x"C0A4B0C0",
   231 => x"C0A4B0F9",
   232 => x"C0A4B0A4",
   233 => x"C0A4B0B0",
   234 => x"C0A4B099",
   235 => x"C0A4B092",
   236 => x"C0A4B082",
   237 => x"C0A4B0F8",
   238 => x"C0A4B080",
   239 => x"C0A4B090",
   240 => x"C0A499C0",
   241 => x"C0A499F9",
   242 => x"C0A499A4",
   243 => x"C0A499B0",
   244 => x"C0A49999",
   245 => x"C0A49992",
   246 => x"C0A49982",
   247 => x"C0A499F8",
   248 => x"C0A49980",
   249 => x"C0A49990",
   250 => x"C0A492C0",
   251 => x"C0A492F9",
   252 => x"C0A492A4",
   253 => x"C0A492B0",
   254 => x"C0A49299",
   255 => x"C0A49292"
);
begin

outp(31 downto 0) <= ROM(to_integer(signed(inp)));
outp(63 downto 32)<= x"C0C0C0C0";

end Behavioral;
