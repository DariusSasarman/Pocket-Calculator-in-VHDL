library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity division_output_processor is
     Port (   
           quotient: in std_logic_vector (7 downto 0);
           remainder:  in std_logic_vector (7 downto 0);
           sign_bit: in std_logic;
           outp : out std_logic_vector (63 downto 0));
end division_output_processor;

architecture Behavioral of division_output_processor is
type rom_type is array (INTEGER RANGE 0 to 255) of std_logic_vector(23 downto 0);
constant ROM : rom_type := (
     0 => x"C0C0C0",
     1 => x"C0C0F9",
     2 => x"C0C0A4",
     3 => x"C0C0B0",
     4 => x"C0C099",
     5 => x"C0C092",
     6 => x"C0C082",
     7 => x"C0C0F8",
     8 => x"C0C080",
     9 => x"C0C090",
    10 => x"C0F9C0",
    11 => x"C0F9F9",
    12 => x"C0F9A4",
    13 => x"C0F9B0",
    14 => x"C0F999",
    15 => x"C0F992",
    16 => x"C0F982",
    17 => x"C0F9F8",
    18 => x"C0F980",
    19 => x"C0F990",
    20 => x"C0A4C0",
    21 => x"C0A4F9",
    22 => x"C0A4A4",
    23 => x"C0A4B0",
    24 => x"C0A499",
    25 => x"C0A492",
    26 => x"C0A482",
    27 => x"C0A4F8",
    28 => x"C0A480",
    29 => x"C0A490",
    30 => x"C0B0C0",
    31 => x"C0B0F9",
    32 => x"C0B0A4",
    33 => x"C0B0B0",
    34 => x"C0B099",
    35 => x"C0B092",
    36 => x"C0B082",
    37 => x"C0B0F8",
    38 => x"C0B080",
    39 => x"C0B090",
    40 => x"C099C0",
    41 => x"C099F9",
    42 => x"C099A4",
    43 => x"C099B0",
    44 => x"C09999",
    45 => x"C09992",
    46 => x"C09982",
    47 => x"C099F8",
    48 => x"C09980",
    49 => x"C09990",
    50 => x"C092C0",
    51 => x"C092F9",
    52 => x"C092A4",
    53 => x"C092B0",
    54 => x"C09299",
    55 => x"C09292",
    56 => x"C09282",
    57 => x"C092F8",
    58 => x"C09280",
    59 => x"C09290",
    60 => x"C082C0",
    61 => x"C082F9",
    62 => x"C082A4",
    63 => x"C082B0",
    64 => x"C08299",
    65 => x"C08292",
    66 => x"C08282",
    67 => x"C082F8",
    68 => x"C08280",
    69 => x"C08290",
    70 => x"C0F8C0",
    71 => x"C0F8F9",
    72 => x"C0F8A4",
    73 => x"C0F8B0",
    74 => x"C0F899",
    75 => x"C0F892",
    76 => x"C0F882",
    77 => x"C0F8F8",
    78 => x"C0F880",
    79 => x"C0F890",
    80 => x"C080C0",
    81 => x"C080F9",
    82 => x"C080A4",
    83 => x"C080B0",
    84 => x"C08099",
    85 => x"C08092",
    86 => x"C08082",
    87 => x"C080F8",
    88 => x"C08080",
    89 => x"C08090",
    90 => x"C090C0",
    91 => x"C090F9",
    92 => x"C090A4",
    93 => x"C090B0",
    94 => x"C09099",
    95 => x"C09092",
    96 => x"C09082",
    97 => x"C090F8",
    98 => x"C09080",
    99 => x"C09090",
   100 => x"F9C0C0",
   101 => x"F9C0F9",
   102 => x"F9C0A4",
   103 => x"F9C0B0",
   104 => x"F9C099",
   105 => x"F9C092",
   106 => x"F9C082",
   107 => x"F9C0F8",
   108 => x"F9C080",
   109 => x"F9C090",
   110 => x"F9F9C0",
   111 => x"F9F9F9",
   112 => x"F9F9A4",
   113 => x"F9F9B0",
   114 => x"F9F999",
   115 => x"F9F992",
   116 => x"F9F982",
   117 => x"F9F9F8",
   118 => x"F9F980",
   119 => x"F9F990",
   120 => x"F9A4C0",
   121 => x"F9A4F9",
   122 => x"F9A4A4",
   123 => x"F9A4B0",
   124 => x"F9A499",
   125 => x"F9A492",
   126 => x"F9A482",
   127 => x"F9A4F8",
   128 => x"F9A480",
   129 => x"F9A490",
   130 => x"F9B0C0",
   131 => x"F9B0F9",
   132 => x"F9B0A4",
   133 => x"F9B0B0",
   134 => x"F9B099",
   135 => x"F9B092",
   136 => x"F9B082",
   137 => x"F9B0F8",
   138 => x"F9B080",
   139 => x"F9B090",
   140 => x"F999C0",
   141 => x"F999F9",
   142 => x"F999A4",
   143 => x"F999B0",
   144 => x"F99999",
   145 => x"F99992",
   146 => x"F99982",
   147 => x"F999F8",
   148 => x"F99980",
   149 => x"F99990",
   150 => x"F992C0",
   151 => x"F992F9",
   152 => x"F992A4",
   153 => x"F992B0",
   154 => x"F99299",
   155 => x"F99292",
   156 => x"F99282",
   157 => x"F992F8",
   158 => x"F99280",
   159 => x"F99290",
   160 => x"F982C0",
   161 => x"F982F9",
   162 => x"F982A4",
   163 => x"F982B0",
   164 => x"F98299",
   165 => x"F98292",
   166 => x"F98282",
   167 => x"F982F8",
   168 => x"F98280",
   169 => x"F98290",
   170 => x"F9F8C0",
   171 => x"F9F8F9",
   172 => x"F9F8A4",
   173 => x"F9F8B0",
   174 => x"F9F899",
   175 => x"F9F892",
   176 => x"F9F882",
   177 => x"F9F8F8",
   178 => x"F9F880",
   179 => x"F9F890",
   180 => x"F980C0",
   181 => x"F980F9",
   182 => x"F980A4",
   183 => x"F980B0",
   184 => x"F98099",
   185 => x"F98092",
   186 => x"F98082",
   187 => x"F980F8",
   188 => x"F98080",
   189 => x"F98090",
   190 => x"F990C0",
   191 => x"F990F9",
   192 => x"F990A4",
   193 => x"F990B0",
   194 => x"F99099",
   195 => x"F99092",
   196 => x"F99082",
   197 => x"F990F8",
   198 => x"F99080",
   199 => x"F99090",
   200 => x"A4C0C0",
   201 => x"A4C0F9",
   202 => x"A4C0A4",
   203 => x"A4C0B0",
   204 => x"A4C099",
   205 => x"A4C092",
   206 => x"A4C082",
   207 => x"A4C0F8",
   208 => x"A4C080",
   209 => x"A4C090",
   210 => x"A4F9C0",
   211 => x"A4F9F9",
   212 => x"A4F9A4",
   213 => x"A4F9B0",
   214 => x"A4F999",
   215 => x"A4F992",
   216 => x"A4F982",
   217 => x"A4F9F8",
   218 => x"A4F980",
   219 => x"A4F990",
   220 => x"A4A4C0",
   221 => x"A4A4F9",
   222 => x"A4A4A4",
   223 => x"A4A4B0",
   224 => x"A4A499",
   225 => x"A4A492",
   226 => x"A4A482",
   227 => x"A4A4F8",
   228 => x"A4A480",
   229 => x"A4A490",
   230 => x"A4B0C0",
   231 => x"A4B0F9",
   232 => x"A4B0A4",
   233 => x"A4B0B0",
   234 => x"A4B099",
   235 => x"A4B092",
   236 => x"A4B082",
   237 => x"A4B0F8",
   238 => x"A4B080",
   239 => x"A4B090",
   240 => x"A499C0",
   241 => x"A499F9",
   242 => x"A499A4",
   243 => x"A499B0",
   244 => x"A49999",
   245 => x"A49992",
   246 => x"A49982",
   247 => x"A499F8",
   248 => x"A49980",
   249 => x"A49990",
   250 => x"A492C0",
   251 => x"A492F9",
   252 => x"A492A4",
   253 => x"A492B0",
   254 => x"A49299",
   255 => x"A49292"
  );

signal sign : std_logic_vector (7 downto 0);

begin

    sign <= x"C0" when sign_bit = '0' else x"BF";
    outp(63 downto 56) <= sign;                    
    outp(55 downto 32) <= ROM(to_integer(unsigned(quotient))); 
    outp(31 downto 24) <= x"AF";                  
    outp(23 downto 0)  <= ROM(to_integer(unsigned(remainder)));  
  
end Behavioral;
