library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity multiplication_output_processor is
    Port (
        inp : in std_Logic_vector (15 downto 0);
        outp: out std_logic_vector(63 downto 0)
     );
end multiplication_output_processor;

architecture Behavioral of multiplication_output_processor is
   type rom_type is array (integer range -32768 to 32767) of std_logic_vector(63 downto 0);
constant ROM : rom_type := (
    -32768 => x"C0C0BFB0A4F88280",
-32767 => x"C0C0BFB0A4F882F8",
-32766 => x"C0C0BFB0A4F88282",
-32765 => x"C0C0BFB0A4F88292",
-32764 => x"C0C0BFB0A4F88299",
-32763 => x"C0C0BFB0A4F882B0",
-32762 => x"C0C0BFB0A4F882A4",
-32761 => x"C0C0BFB0A4F882F9",
-32760 => x"C0C0BFB0A4F882C0",
-32759 => x"C0C0BFB0A4F89290",
-32758 => x"C0C0BFB0A4F89280",
-32757 => x"C0C0BFB0A4F892F8",
-32756 => x"C0C0BFB0A4F89282",
-32755 => x"C0C0BFB0A4F89292",
-32754 => x"C0C0BFB0A4F89299",
-32753 => x"C0C0BFB0A4F892B0",
-32752 => x"C0C0BFB0A4F892A4",
-32751 => x"C0C0BFB0A4F892F9",
-32750 => x"C0C0BFB0A4F892C0",
-32749 => x"C0C0BFB0A4F89990",
-32748 => x"C0C0BFB0A4F89980",
-32747 => x"C0C0BFB0A4F899F8",
-32746 => x"C0C0BFB0A4F89982",
-32745 => x"C0C0BFB0A4F89992",
-32744 => x"C0C0BFB0A4F89999",
-32743 => x"C0C0BFB0A4F899B0",
-32742 => x"C0C0BFB0A4F899A4",
-32741 => x"C0C0BFB0A4F899F9",
-32740 => x"C0C0BFB0A4F899C0",
-32739 => x"C0C0BFB0A4F8B090",
-32738 => x"C0C0BFB0A4F8B080",
-32737 => x"C0C0BFB0A4F8B0F8",
-32736 => x"C0C0BFB0A4F8B082",
-32735 => x"C0C0BFB0A4F8B092",
-32734 => x"C0C0BFB0A4F8B099",
-32733 => x"C0C0BFB0A4F8B0B0",
-32732 => x"C0C0BFB0A4F8B0A4",
-32731 => x"C0C0BFB0A4F8B0F9",
-32730 => x"C0C0BFB0A4F8B0C0",
-32729 => x"C0C0BFB0A4F8A490",
-32728 => x"C0C0BFB0A4F8A480",
-32727 => x"C0C0BFB0A4F8A4F8",
-32726 => x"C0C0BFB0A4F8A482",
-32725 => x"C0C0BFB0A4F8A492",
-32724 => x"C0C0BFB0A4F8A499",
-32723 => x"C0C0BFB0A4F8A4B0",
-32722 => x"C0C0BFB0A4F8A4A4",
-32721 => x"C0C0BFB0A4F8A4F9",
-32720 => x"C0C0BFB0A4F8A4C0",
-32719 => x"C0C0BFB0A4F8F990",
-32718 => x"C0C0BFB0A4F8F980",
-32717 => x"C0C0BFB0A4F8F9F8",
-32716 => x"C0C0BFB0A4F8F982",
-32715 => x"C0C0BFB0A4F8F992",
-32714 => x"C0C0BFB0A4F8F999",
-32713 => x"C0C0BFB0A4F8F9B0",
-32712 => x"C0C0BFB0A4F8F9A4",
-32711 => x"C0C0BFB0A4F8F9F9",
-32710 => x"C0C0BFB0A4F8F9C0",
-32709 => x"C0C0BFB0A4F8C090",
-32708 => x"C0C0BFB0A4F8C080",
-32707 => x"C0C0BFB0A4F8C0F8",
-32706 => x"C0C0BFB0A4F8C082",
-32705 => x"C0C0BFB0A4F8C092",
-32704 => x"C0C0BFB0A4F8C099",
-32703 => x"C0C0BFB0A4F8C0B0",
-32702 => x"C0C0BFB0A4F8C0A4",
-32701 => x"C0C0BFB0A4F8C0F9",
-32700 => x"C0C0BFB0A4F8C0C0",
-32699 => x"C0C0BFB0A4829090",
-32698 => x"C0C0BFB0A4829080",
-32697 => x"C0C0BFB0A48290F8",
-32696 => x"C0C0BFB0A4829082",
-32695 => x"C0C0BFB0A4829092",
-32694 => x"C0C0BFB0A4829099",
-32693 => x"C0C0BFB0A48290B0",
-32692 => x"C0C0BFB0A48290A4",
-32691 => x"C0C0BFB0A48290F9",
-32690 => x"C0C0BFB0A48290C0",
-32689 => x"C0C0BFB0A4828090",
-32688 => x"C0C0BFB0A4828080",
-32687 => x"C0C0BFB0A48280F8",
-32686 => x"C0C0BFB0A4828082",
-32685 => x"C0C0BFB0A4828092",
-32684 => x"C0C0BFB0A4828099",
-32683 => x"C0C0BFB0A48280B0",
-32682 => x"C0C0BFB0A48280A4",
-32681 => x"C0C0BFB0A48280F9",
-32680 => x"C0C0BFB0A48280C0",
-32679 => x"C0C0BFB0A482F890",
-32678 => x"C0C0BFB0A482F880",
-32677 => x"C0C0BFB0A482F8F8",
-32676 => x"C0C0BFB0A482F882",
-32675 => x"C0C0BFB0A482F892",
-32674 => x"C0C0BFB0A482F899",
-32673 => x"C0C0BFB0A482F8B0",
-32672 => x"C0C0BFB0A482F8A4",
-32671 => x"C0C0BFB0A482F8F9",
-32670 => x"C0C0BFB0A482F8C0",
-32669 => x"C0C0BFB0A4828290",
-32668 => x"C0C0BFB0A4828280",
-32667 => x"C0C0BFB0A48282F8",
-32666 => x"C0C0BFB0A4828282",
-32665 => x"C0C0BFB0A4828292",
-32664 => x"C0C0BFB0A4828299",
-32663 => x"C0C0BFB0A48282B0",
-32662 => x"C0C0BFB0A48282A4",
-32661 => x"C0C0BFB0A48282F9",
-32660 => x"C0C0BFB0A48282C0",
-32659 => x"C0C0BFB0A4829290",
-32658 => x"C0C0BFB0A4829280",
-32657 => x"C0C0BFB0A48292F8",
-32656 => x"C0C0BFB0A4829282",
-32655 => x"C0C0BFB0A4829292",
-32654 => x"C0C0BFB0A4829299",
-32653 => x"C0C0BFB0A48292B0",
-32652 => x"C0C0BFB0A48292A4",
-32651 => x"C0C0BFB0A48292F9",
-32650 => x"C0C0BFB0A48292C0",
-32649 => x"C0C0BFB0A4829990",
-32648 => x"C0C0BFB0A4829980",
-32647 => x"C0C0BFB0A48299F8",
-32646 => x"C0C0BFB0A4829982",
-32645 => x"C0C0BFB0A4829992",
-32644 => x"C0C0BFB0A4829999",
-32643 => x"C0C0BFB0A48299B0",
-32642 => x"C0C0BFB0A48299A4",
-32641 => x"C0C0BFB0A48299F9",
-32640 => x"C0C0BFB0A48299C0",
-32639 => x"C0C0BFB0A482B090",
-32638 => x"C0C0BFB0A482B080",
-32637 => x"C0C0BFB0A482B0F8",
-32636 => x"C0C0BFB0A482B082",
-32635 => x"C0C0BFB0A482B092",
-32634 => x"C0C0BFB0A482B099",
-32633 => x"C0C0BFB0A482B0B0",
-32632 => x"C0C0BFB0A482B0A4",
-32631 => x"C0C0BFB0A482B0F9",
-32630 => x"C0C0BFB0A482B0C0",
-32629 => x"C0C0BFB0A482A490",
-32628 => x"C0C0BFB0A482A480",
-32627 => x"C0C0BFB0A482A4F8",
-32626 => x"C0C0BFB0A482A482",
-32625 => x"C0C0BFB0A482A492",
-32624 => x"C0C0BFB0A482A499",
-32623 => x"C0C0BFB0A482A4B0",
-32622 => x"C0C0BFB0A482A4A4",
-32621 => x"C0C0BFB0A482A4F9",
-32620 => x"C0C0BFB0A482A4C0",
-32619 => x"C0C0BFB0A482F990",
-32618 => x"C0C0BFB0A482F980",
-32617 => x"C0C0BFB0A482F9F8",
-32616 => x"C0C0BFB0A482F982",
-32615 => x"C0C0BFB0A482F992",
-32614 => x"C0C0BFB0A482F999",
-32613 => x"C0C0BFB0A482F9B0",
-32612 => x"C0C0BFB0A482F9A4",
-32611 => x"C0C0BFB0A482F9F9",
-32610 => x"C0C0BFB0A482F9C0",
-32609 => x"C0C0BFB0A482C090",
-32608 => x"C0C0BFB0A482C080",
-32607 => x"C0C0BFB0A482C0F8",
-32606 => x"C0C0BFB0A482C082",
-32605 => x"C0C0BFB0A482C092",
-32604 => x"C0C0BFB0A482C099",
-32603 => x"C0C0BFB0A482C0B0",
-32602 => x"C0C0BFB0A482C0A4",
-32601 => x"C0C0BFB0A482C0F9",
-32600 => x"C0C0BFB0A482C0C0",
-32599 => x"C0C0BFB0A4929090",
-32598 => x"C0C0BFB0A4929080",
-32597 => x"C0C0BFB0A49290F8",
-32596 => x"C0C0BFB0A4929082",
-32595 => x"C0C0BFB0A4929092",
-32594 => x"C0C0BFB0A4929099",
-32593 => x"C0C0BFB0A49290B0",
-32592 => x"C0C0BFB0A49290A4",
-32591 => x"C0C0BFB0A49290F9",
-32590 => x"C0C0BFB0A49290C0",
-32589 => x"C0C0BFB0A4928090",
-32588 => x"C0C0BFB0A4928080",
-32587 => x"C0C0BFB0A49280F8",
-32586 => x"C0C0BFB0A4928082",
-32585 => x"C0C0BFB0A4928092",
-32584 => x"C0C0BFB0A4928099",
-32583 => x"C0C0BFB0A49280B0",
-32582 => x"C0C0BFB0A49280A4",
-32581 => x"C0C0BFB0A49280F9",
-32580 => x"C0C0BFB0A49280C0",
-32579 => x"C0C0BFB0A492F890",
-32578 => x"C0C0BFB0A492F880",
-32577 => x"C0C0BFB0A492F8F8",
-32576 => x"C0C0BFB0A492F882",
-32575 => x"C0C0BFB0A492F892",
-32574 => x"C0C0BFB0A492F899",
-32573 => x"C0C0BFB0A492F8B0",
-32572 => x"C0C0BFB0A492F8A4",
-32571 => x"C0C0BFB0A492F8F9",
-32570 => x"C0C0BFB0A492F8C0",
-32569 => x"C0C0BFB0A4928290",
-32568 => x"C0C0BFB0A4928280",
-32567 => x"C0C0BFB0A49282F8",
-32566 => x"C0C0BFB0A4928282",
-32565 => x"C0C0BFB0A4928292",
-32564 => x"C0C0BFB0A4928299",
-32563 => x"C0C0BFB0A49282B0",
-32562 => x"C0C0BFB0A49282A4",
-32561 => x"C0C0BFB0A49282F9",
-32560 => x"C0C0BFB0A49282C0",
-32559 => x"C0C0BFB0A4929290",
-32558 => x"C0C0BFB0A4929280",
-32557 => x"C0C0BFB0A49292F8",
-32556 => x"C0C0BFB0A4929282",
-32555 => x"C0C0BFB0A4929292",
-32554 => x"C0C0BFB0A4929299",
-32553 => x"C0C0BFB0A49292B0",
-32552 => x"C0C0BFB0A49292A4",
-32551 => x"C0C0BFB0A49292F9",
-32550 => x"C0C0BFB0A49292C0",
-32549 => x"C0C0BFB0A4929990",
-32548 => x"C0C0BFB0A4929980",
-32547 => x"C0C0BFB0A49299F8",
-32546 => x"C0C0BFB0A4929982",
-32545 => x"C0C0BFB0A4929992",
-32544 => x"C0C0BFB0A4929999",
-32543 => x"C0C0BFB0A49299B0",
-32542 => x"C0C0BFB0A49299A4",
-32541 => x"C0C0BFB0A49299F9",
-32540 => x"C0C0BFB0A49299C0",
-32539 => x"C0C0BFB0A492B090",
-32538 => x"C0C0BFB0A492B080",
-32537 => x"C0C0BFB0A492B0F8",
-32536 => x"C0C0BFB0A492B082",
-32535 => x"C0C0BFB0A492B092",
-32534 => x"C0C0BFB0A492B099",
-32533 => x"C0C0BFB0A492B0B0",
-32532 => x"C0C0BFB0A492B0A4",
-32531 => x"C0C0BFB0A492B0F9",
-32530 => x"C0C0BFB0A492B0C0",
-32529 => x"C0C0BFB0A492A490",
-32528 => x"C0C0BFB0A492A480",
-32527 => x"C0C0BFB0A492A4F8",
-32526 => x"C0C0BFB0A492A482",
-32525 => x"C0C0BFB0A492A492",
-32524 => x"C0C0BFB0A492A499",
-32523 => x"C0C0BFB0A492A4B0",
-32522 => x"C0C0BFB0A492A4A4",
-32521 => x"C0C0BFB0A492A4F9",
-32520 => x"C0C0BFB0A492A4C0",
-32519 => x"C0C0BFB0A492F990",
-32518 => x"C0C0BFB0A492F980",
-32517 => x"C0C0BFB0A492F9F8",
-32516 => x"C0C0BFB0A492F982",
-32515 => x"C0C0BFB0A492F992",
-32514 => x"C0C0BFB0A492F999",
-32513 => x"C0C0BFB0A492F9B0",
-32512 => x"C0C0BFB0A492F9A4",
-32511 => x"C0C0BFB0A492F9F9",
-32510 => x"C0C0BFB0A492F9C0",
-32509 => x"C0C0BFB0A492C090",
-32508 => x"C0C0BFB0A492C080",
-32507 => x"C0C0BFB0A492C0F8",
-32506 => x"C0C0BFB0A492C082",
-32505 => x"C0C0BFB0A492C092",
-32504 => x"C0C0BFB0A492C099",
-32503 => x"C0C0BFB0A492C0B0",
-32502 => x"C0C0BFB0A492C0A4",
-32501 => x"C0C0BFB0A492C0F9",
-32500 => x"C0C0BFB0A492C0C0",
-32499 => x"C0C0BFB0A4999090",
-32498 => x"C0C0BFB0A4999080",
-32497 => x"C0C0BFB0A49990F8",
-32496 => x"C0C0BFB0A4999082",
-32495 => x"C0C0BFB0A4999092",
-32494 => x"C0C0BFB0A4999099",
-32493 => x"C0C0BFB0A49990B0",
-32492 => x"C0C0BFB0A49990A4",
-32491 => x"C0C0BFB0A49990F9",
-32490 => x"C0C0BFB0A49990C0",
-32489 => x"C0C0BFB0A4998090",
-32488 => x"C0C0BFB0A4998080",
-32487 => x"C0C0BFB0A49980F8",
-32486 => x"C0C0BFB0A4998082",
-32485 => x"C0C0BFB0A4998092",
-32484 => x"C0C0BFB0A4998099",
-32483 => x"C0C0BFB0A49980B0",
-32482 => x"C0C0BFB0A49980A4",
-32481 => x"C0C0BFB0A49980F9",
-32480 => x"C0C0BFB0A49980C0",
-32479 => x"C0C0BFB0A499F890",
-32478 => x"C0C0BFB0A499F880",
-32477 => x"C0C0BFB0A499F8F8",
-32476 => x"C0C0BFB0A499F882",
-32475 => x"C0C0BFB0A499F892",
-32474 => x"C0C0BFB0A499F899",
-32473 => x"C0C0BFB0A499F8B0",
-32472 => x"C0C0BFB0A499F8A4",
-32471 => x"C0C0BFB0A499F8F9",
-32470 => x"C0C0BFB0A499F8C0",
-32469 => x"C0C0BFB0A4998290",
-32468 => x"C0C0BFB0A4998280",
-32467 => x"C0C0BFB0A49982F8",
-32466 => x"C0C0BFB0A4998282",
-32465 => x"C0C0BFB0A4998292",
-32464 => x"C0C0BFB0A4998299",
-32463 => x"C0C0BFB0A49982B0",
-32462 => x"C0C0BFB0A49982A4",
-32461 => x"C0C0BFB0A49982F9",
-32460 => x"C0C0BFB0A49982C0",
-32459 => x"C0C0BFB0A4999290",
-32458 => x"C0C0BFB0A4999280",
-32457 => x"C0C0BFB0A49992F8",
-32456 => x"C0C0BFB0A4999282",
-32455 => x"C0C0BFB0A4999292",
-32454 => x"C0C0BFB0A4999299",
-32453 => x"C0C0BFB0A49992B0",
-32452 => x"C0C0BFB0A49992A4",
-32451 => x"C0C0BFB0A49992F9",
-32450 => x"C0C0BFB0A49992C0",
-32449 => x"C0C0BFB0A4999990",
-32448 => x"C0C0BFB0A4999980",
-32447 => x"C0C0BFB0A49999F8",
-32446 => x"C0C0BFB0A4999982",
-32445 => x"C0C0BFB0A4999992",
-32444 => x"C0C0BFB0A4999999",
-32443 => x"C0C0BFB0A49999B0",
-32442 => x"C0C0BFB0A49999A4",
-32441 => x"C0C0BFB0A49999F9",
-32440 => x"C0C0BFB0A49999C0",
-32439 => x"C0C0BFB0A499B090",
-32438 => x"C0C0BFB0A499B080",
-32437 => x"C0C0BFB0A499B0F8",
-32436 => x"C0C0BFB0A499B082",
-32435 => x"C0C0BFB0A499B092",
-32434 => x"C0C0BFB0A499B099",
-32433 => x"C0C0BFB0A499B0B0",
-32432 => x"C0C0BFB0A499B0A4",
-32431 => x"C0C0BFB0A499B0F9",
-32430 => x"C0C0BFB0A499B0C0",
-32429 => x"C0C0BFB0A499A490",
-32428 => x"C0C0BFB0A499A480",
-32427 => x"C0C0BFB0A499A4F8",
-32426 => x"C0C0BFB0A499A482",
-32425 => x"C0C0BFB0A499A492",
-32424 => x"C0C0BFB0A499A499",
-32423 => x"C0C0BFB0A499A4B0",
-32422 => x"C0C0BFB0A499A4A4",
-32421 => x"C0C0BFB0A499A4F9",
-32420 => x"C0C0BFB0A499A4C0",
-32419 => x"C0C0BFB0A499F990",
-32418 => x"C0C0BFB0A499F980",
-32417 => x"C0C0BFB0A499F9F8",
-32416 => x"C0C0BFB0A499F982",
-32415 => x"C0C0BFB0A499F992",
-32414 => x"C0C0BFB0A499F999",
-32413 => x"C0C0BFB0A499F9B0",
-32412 => x"C0C0BFB0A499F9A4",
-32411 => x"C0C0BFB0A499F9F9",
-32410 => x"C0C0BFB0A499F9C0",
-32409 => x"C0C0BFB0A499C090",
-32408 => x"C0C0BFB0A499C080",
-32407 => x"C0C0BFB0A499C0F8",
-32406 => x"C0C0BFB0A499C082",
-32405 => x"C0C0BFB0A499C092",
-32404 => x"C0C0BFB0A499C099",
-32403 => x"C0C0BFB0A499C0B0",
-32402 => x"C0C0BFB0A499C0A4",
-32401 => x"C0C0BFB0A499C0F9",
-32400 => x"C0C0BFB0A499C0C0",
-32399 => x"C0C0BFB0A4B09090",
-32398 => x"C0C0BFB0A4B09080",
-32397 => x"C0C0BFB0A4B090F8",
-32396 => x"C0C0BFB0A4B09082",
-32395 => x"C0C0BFB0A4B09092",
-32394 => x"C0C0BFB0A4B09099",
-32393 => x"C0C0BFB0A4B090B0",
-32392 => x"C0C0BFB0A4B090A4",
-32391 => x"C0C0BFB0A4B090F9",
-32390 => x"C0C0BFB0A4B090C0",
-32389 => x"C0C0BFB0A4B08090",
-32388 => x"C0C0BFB0A4B08080",
-32387 => x"C0C0BFB0A4B080F8",
-32386 => x"C0C0BFB0A4B08082",
-32385 => x"C0C0BFB0A4B08092",
-32384 => x"C0C0BFB0A4B08099",
-32383 => x"C0C0BFB0A4B080B0",
-32382 => x"C0C0BFB0A4B080A4",
-32381 => x"C0C0BFB0A4B080F9",
-32380 => x"C0C0BFB0A4B080C0",
-32379 => x"C0C0BFB0A4B0F890",
-32378 => x"C0C0BFB0A4B0F880",
-32377 => x"C0C0BFB0A4B0F8F8",
-32376 => x"C0C0BFB0A4B0F882",
-32375 => x"C0C0BFB0A4B0F892",
-32374 => x"C0C0BFB0A4B0F899",
-32373 => x"C0C0BFB0A4B0F8B0",
-32372 => x"C0C0BFB0A4B0F8A4",
-32371 => x"C0C0BFB0A4B0F8F9",
-32370 => x"C0C0BFB0A4B0F8C0",
-32369 => x"C0C0BFB0A4B08290",
-32368 => x"C0C0BFB0A4B08280",
-32367 => x"C0C0BFB0A4B082F8",
-32366 => x"C0C0BFB0A4B08282",
-32365 => x"C0C0BFB0A4B08292",
-32364 => x"C0C0BFB0A4B08299",
-32363 => x"C0C0BFB0A4B082B0",
-32362 => x"C0C0BFB0A4B082A4",
-32361 => x"C0C0BFB0A4B082F9",
-32360 => x"C0C0BFB0A4B082C0",
-32359 => x"C0C0BFB0A4B09290",
-32358 => x"C0C0BFB0A4B09280",
-32357 => x"C0C0BFB0A4B092F8",
-32356 => x"C0C0BFB0A4B09282",
-32355 => x"C0C0BFB0A4B09292",
-32354 => x"C0C0BFB0A4B09299",
-32353 => x"C0C0BFB0A4B092B0",
-32352 => x"C0C0BFB0A4B092A4",
-32351 => x"C0C0BFB0A4B092F9",
-32350 => x"C0C0BFB0A4B092C0",
-32349 => x"C0C0BFB0A4B09990",
-32348 => x"C0C0BFB0A4B09980",
-32347 => x"C0C0BFB0A4B099F8",
-32346 => x"C0C0BFB0A4B09982",
-32345 => x"C0C0BFB0A4B09992",
-32344 => x"C0C0BFB0A4B09999",
-32343 => x"C0C0BFB0A4B099B0",
-32342 => x"C0C0BFB0A4B099A4",
-32341 => x"C0C0BFB0A4B099F9",
-32340 => x"C0C0BFB0A4B099C0",
-32339 => x"C0C0BFB0A4B0B090",
-32338 => x"C0C0BFB0A4B0B080",
-32337 => x"C0C0BFB0A4B0B0F8",
-32336 => x"C0C0BFB0A4B0B082",
-32335 => x"C0C0BFB0A4B0B092",
-32334 => x"C0C0BFB0A4B0B099",
-32333 => x"C0C0BFB0A4B0B0B0",
-32332 => x"C0C0BFB0A4B0B0A4",
-32331 => x"C0C0BFB0A4B0B0F9",
-32330 => x"C0C0BFB0A4B0B0C0",
-32329 => x"C0C0BFB0A4B0A490",
-32328 => x"C0C0BFB0A4B0A480",
-32327 => x"C0C0BFB0A4B0A4F8",
-32326 => x"C0C0BFB0A4B0A482",
-32325 => x"C0C0BFB0A4B0A492",
-32324 => x"C0C0BFB0A4B0A499",
-32323 => x"C0C0BFB0A4B0A4B0",
-32322 => x"C0C0BFB0A4B0A4A4",
-32321 => x"C0C0BFB0A4B0A4F9",
-32320 => x"C0C0BFB0A4B0A4C0",
-32319 => x"C0C0BFB0A4B0F990",
-32318 => x"C0C0BFB0A4B0F980",
-32317 => x"C0C0BFB0A4B0F9F8",
-32316 => x"C0C0BFB0A4B0F982",
-32315 => x"C0C0BFB0A4B0F992",
-32314 => x"C0C0BFB0A4B0F999",
-32313 => x"C0C0BFB0A4B0F9B0",
-32312 => x"C0C0BFB0A4B0F9A4",
-32311 => x"C0C0BFB0A4B0F9F9",
-32310 => x"C0C0BFB0A4B0F9C0",
-32309 => x"C0C0BFB0A4B0C090",
-32308 => x"C0C0BFB0A4B0C080",
-32307 => x"C0C0BFB0A4B0C0F8",
-32306 => x"C0C0BFB0A4B0C082",
-32305 => x"C0C0BFB0A4B0C092",
-32304 => x"C0C0BFB0A4B0C099",
-32303 => x"C0C0BFB0A4B0C0B0",
-32302 => x"C0C0BFB0A4B0C0A4",
-32301 => x"C0C0BFB0A4B0C0F9",
-32300 => x"C0C0BFB0A4B0C0C0",
-32299 => x"C0C0BFB0A4A49090",
-32298 => x"C0C0BFB0A4A49080",
-32297 => x"C0C0BFB0A4A490F8",
-32296 => x"C0C0BFB0A4A49082",
-32295 => x"C0C0BFB0A4A49092",
-32294 => x"C0C0BFB0A4A49099",
-32293 => x"C0C0BFB0A4A490B0",
-32292 => x"C0C0BFB0A4A490A4",
-32291 => x"C0C0BFB0A4A490F9",
-32290 => x"C0C0BFB0A4A490C0",
-32289 => x"C0C0BFB0A4A48090",
-32288 => x"C0C0BFB0A4A48080",
-32287 => x"C0C0BFB0A4A480F8",
-32286 => x"C0C0BFB0A4A48082",
-32285 => x"C0C0BFB0A4A48092",
-32284 => x"C0C0BFB0A4A48099",
-32283 => x"C0C0BFB0A4A480B0",
-32282 => x"C0C0BFB0A4A480A4",
-32281 => x"C0C0BFB0A4A480F9",
-32280 => x"C0C0BFB0A4A480C0",
-32279 => x"C0C0BFB0A4A4F890",
-32278 => x"C0C0BFB0A4A4F880",
-32277 => x"C0C0BFB0A4A4F8F8",
-32276 => x"C0C0BFB0A4A4F882",
-32275 => x"C0C0BFB0A4A4F892",
-32274 => x"C0C0BFB0A4A4F899",
-32273 => x"C0C0BFB0A4A4F8B0",
-32272 => x"C0C0BFB0A4A4F8A4",
-32271 => x"C0C0BFB0A4A4F8F9",
-32270 => x"C0C0BFB0A4A4F8C0",
-32269 => x"C0C0BFB0A4A48290",
-32268 => x"C0C0BFB0A4A48280",
-32267 => x"C0C0BFB0A4A482F8",
-32266 => x"C0C0BFB0A4A48282",
-32265 => x"C0C0BFB0A4A48292",
-32264 => x"C0C0BFB0A4A48299",
-32263 => x"C0C0BFB0A4A482B0",
-32262 => x"C0C0BFB0A4A482A4",
-32261 => x"C0C0BFB0A4A482F9",
-32260 => x"C0C0BFB0A4A482C0",
-32259 => x"C0C0BFB0A4A49290",
-32258 => x"C0C0BFB0A4A49280",
-32257 => x"C0C0BFB0A4A492F8",
-32256 => x"C0C0BFB0A4A49282",
-32255 => x"C0C0BFB0A4A49292",
-32254 => x"C0C0BFB0A4A49299",
-32253 => x"C0C0BFB0A4A492B0",
-32252 => x"C0C0BFB0A4A492A4",
-32251 => x"C0C0BFB0A4A492F9",
-32250 => x"C0C0BFB0A4A492C0",
-32249 => x"C0C0BFB0A4A49990",
-32248 => x"C0C0BFB0A4A49980",
-32247 => x"C0C0BFB0A4A499F8",
-32246 => x"C0C0BFB0A4A49982",
-32245 => x"C0C0BFB0A4A49992",
-32244 => x"C0C0BFB0A4A49999",
-32243 => x"C0C0BFB0A4A499B0",
-32242 => x"C0C0BFB0A4A499A4",
-32241 => x"C0C0BFB0A4A499F9",
-32240 => x"C0C0BFB0A4A499C0",
-32239 => x"C0C0BFB0A4A4B090",
-32238 => x"C0C0BFB0A4A4B080",
-32237 => x"C0C0BFB0A4A4B0F8",
-32236 => x"C0C0BFB0A4A4B082",
-32235 => x"C0C0BFB0A4A4B092",
-32234 => x"C0C0BFB0A4A4B099",
-32233 => x"C0C0BFB0A4A4B0B0",
-32232 => x"C0C0BFB0A4A4B0A4",
-32231 => x"C0C0BFB0A4A4B0F9",
-32230 => x"C0C0BFB0A4A4B0C0",
-32229 => x"C0C0BFB0A4A4A490",
-32228 => x"C0C0BFB0A4A4A480",
-32227 => x"C0C0BFB0A4A4A4F8",
-32226 => x"C0C0BFB0A4A4A482",
-32225 => x"C0C0BFB0A4A4A492",
-32224 => x"C0C0BFB0A4A4A499",
-32223 => x"C0C0BFB0A4A4A4B0",
-32222 => x"C0C0BFB0A4A4A4A4",
-32221 => x"C0C0BFB0A4A4A4F9",
-32220 => x"C0C0BFB0A4A4A4C0",
-32219 => x"C0C0BFB0A4A4F990",
-32218 => x"C0C0BFB0A4A4F980",
-32217 => x"C0C0BFB0A4A4F9F8",
-32216 => x"C0C0BFB0A4A4F982",
-32215 => x"C0C0BFB0A4A4F992",
-32214 => x"C0C0BFB0A4A4F999",
-32213 => x"C0C0BFB0A4A4F9B0",
-32212 => x"C0C0BFB0A4A4F9A4",
-32211 => x"C0C0BFB0A4A4F9F9",
-32210 => x"C0C0BFB0A4A4F9C0",
-32209 => x"C0C0BFB0A4A4C090",
-32208 => x"C0C0BFB0A4A4C080",
-32207 => x"C0C0BFB0A4A4C0F8",
-32206 => x"C0C0BFB0A4A4C082",
-32205 => x"C0C0BFB0A4A4C092",
-32204 => x"C0C0BFB0A4A4C099",
-32203 => x"C0C0BFB0A4A4C0B0",
-32202 => x"C0C0BFB0A4A4C0A4",
-32201 => x"C0C0BFB0A4A4C0F9",
-32200 => x"C0C0BFB0A4A4C0C0",
-32199 => x"C0C0BFB0A4F99090",
-32198 => x"C0C0BFB0A4F99080",
-32197 => x"C0C0BFB0A4F990F8",
-32196 => x"C0C0BFB0A4F99082",
-32195 => x"C0C0BFB0A4F99092",
-32194 => x"C0C0BFB0A4F99099",
-32193 => x"C0C0BFB0A4F990B0",
-32192 => x"C0C0BFB0A4F990A4",
-32191 => x"C0C0BFB0A4F990F9",
-32190 => x"C0C0BFB0A4F990C0",
-32189 => x"C0C0BFB0A4F98090",
-32188 => x"C0C0BFB0A4F98080",
-32187 => x"C0C0BFB0A4F980F8",
-32186 => x"C0C0BFB0A4F98082",
-32185 => x"C0C0BFB0A4F98092",
-32184 => x"C0C0BFB0A4F98099",
-32183 => x"C0C0BFB0A4F980B0",
-32182 => x"C0C0BFB0A4F980A4",
-32181 => x"C0C0BFB0A4F980F9",
-32180 => x"C0C0BFB0A4F980C0",
-32179 => x"C0C0BFB0A4F9F890",
-32178 => x"C0C0BFB0A4F9F880",
-32177 => x"C0C0BFB0A4F9F8F8",
-32176 => x"C0C0BFB0A4F9F882",
-32175 => x"C0C0BFB0A4F9F892",
-32174 => x"C0C0BFB0A4F9F899",
-32173 => x"C0C0BFB0A4F9F8B0",
-32172 => x"C0C0BFB0A4F9F8A4",
-32171 => x"C0C0BFB0A4F9F8F9",
-32170 => x"C0C0BFB0A4F9F8C0",
-32169 => x"C0C0BFB0A4F98290",
-32168 => x"C0C0BFB0A4F98280",
-32167 => x"C0C0BFB0A4F982F8",
-32166 => x"C0C0BFB0A4F98282",
-32165 => x"C0C0BFB0A4F98292",
-32164 => x"C0C0BFB0A4F98299",
-32163 => x"C0C0BFB0A4F982B0",
-32162 => x"C0C0BFB0A4F982A4",
-32161 => x"C0C0BFB0A4F982F9",
-32160 => x"C0C0BFB0A4F982C0",
-32159 => x"C0C0BFB0A4F99290",
-32158 => x"C0C0BFB0A4F99280",
-32157 => x"C0C0BFB0A4F992F8",
-32156 => x"C0C0BFB0A4F99282",
-32155 => x"C0C0BFB0A4F99292",
-32154 => x"C0C0BFB0A4F99299",
-32153 => x"C0C0BFB0A4F992B0",
-32152 => x"C0C0BFB0A4F992A4",
-32151 => x"C0C0BFB0A4F992F9",
-32150 => x"C0C0BFB0A4F992C0",
-32149 => x"C0C0BFB0A4F99990",
-32148 => x"C0C0BFB0A4F99980",
-32147 => x"C0C0BFB0A4F999F8",
-32146 => x"C0C0BFB0A4F99982",
-32145 => x"C0C0BFB0A4F99992",
-32144 => x"C0C0BFB0A4F99999",
-32143 => x"C0C0BFB0A4F999B0",
-32142 => x"C0C0BFB0A4F999A4",
-32141 => x"C0C0BFB0A4F999F9",
-32140 => x"C0C0BFB0A4F999C0",
-32139 => x"C0C0BFB0A4F9B090",
-32138 => x"C0C0BFB0A4F9B080",
-32137 => x"C0C0BFB0A4F9B0F8",
-32136 => x"C0C0BFB0A4F9B082",
-32135 => x"C0C0BFB0A4F9B092",
-32134 => x"C0C0BFB0A4F9B099",
-32133 => x"C0C0BFB0A4F9B0B0",
-32132 => x"C0C0BFB0A4F9B0A4",
-32131 => x"C0C0BFB0A4F9B0F9",
-32130 => x"C0C0BFB0A4F9B0C0",
-32129 => x"C0C0BFB0A4F9A490",
-32128 => x"C0C0BFB0A4F9A480",
-32127 => x"C0C0BFB0A4F9A4F8",
-32126 => x"C0C0BFB0A4F9A482",
-32125 => x"C0C0BFB0A4F9A492",
-32124 => x"C0C0BFB0A4F9A499",
-32123 => x"C0C0BFB0A4F9A4B0",
-32122 => x"C0C0BFB0A4F9A4A4",
-32121 => x"C0C0BFB0A4F9A4F9",
-32120 => x"C0C0BFB0A4F9A4C0",
-32119 => x"C0C0BFB0A4F9F990",
-32118 => x"C0C0BFB0A4F9F980",
-32117 => x"C0C0BFB0A4F9F9F8",
-32116 => x"C0C0BFB0A4F9F982",
-32115 => x"C0C0BFB0A4F9F992",
-32114 => x"C0C0BFB0A4F9F999",
-32113 => x"C0C0BFB0A4F9F9B0",
-32112 => x"C0C0BFB0A4F9F9A4",
-32111 => x"C0C0BFB0A4F9F9F9",
-32110 => x"C0C0BFB0A4F9F9C0",
-32109 => x"C0C0BFB0A4F9C090",
-32108 => x"C0C0BFB0A4F9C080",
-32107 => x"C0C0BFB0A4F9C0F8",
-32106 => x"C0C0BFB0A4F9C082",
-32105 => x"C0C0BFB0A4F9C092",
-32104 => x"C0C0BFB0A4F9C099",
-32103 => x"C0C0BFB0A4F9C0B0",
-32102 => x"C0C0BFB0A4F9C0A4",
-32101 => x"C0C0BFB0A4F9C0F9",
-32100 => x"C0C0BFB0A4F9C0C0",
-32099 => x"C0C0BFB0A4C09090",
-32098 => x"C0C0BFB0A4C09080",
-32097 => x"C0C0BFB0A4C090F8",
-32096 => x"C0C0BFB0A4C09082",
-32095 => x"C0C0BFB0A4C09092",
-32094 => x"C0C0BFB0A4C09099",
-32093 => x"C0C0BFB0A4C090B0",
-32092 => x"C0C0BFB0A4C090A4",
-32091 => x"C0C0BFB0A4C090F9",
-32090 => x"C0C0BFB0A4C090C0",
-32089 => x"C0C0BFB0A4C08090",
-32088 => x"C0C0BFB0A4C08080",
-32087 => x"C0C0BFB0A4C080F8",
-32086 => x"C0C0BFB0A4C08082",
-32085 => x"C0C0BFB0A4C08092",
-32084 => x"C0C0BFB0A4C08099",
-32083 => x"C0C0BFB0A4C080B0",
-32082 => x"C0C0BFB0A4C080A4",
-32081 => x"C0C0BFB0A4C080F9",
-32080 => x"C0C0BFB0A4C080C0",
-32079 => x"C0C0BFB0A4C0F890",
-32078 => x"C0C0BFB0A4C0F880",
-32077 => x"C0C0BFB0A4C0F8F8",
-32076 => x"C0C0BFB0A4C0F882",
-32075 => x"C0C0BFB0A4C0F892",
-32074 => x"C0C0BFB0A4C0F899",
-32073 => x"C0C0BFB0A4C0F8B0",
-32072 => x"C0C0BFB0A4C0F8A4",
-32071 => x"C0C0BFB0A4C0F8F9",
-32070 => x"C0C0BFB0A4C0F8C0",
-32069 => x"C0C0BFB0A4C08290",
-32068 => x"C0C0BFB0A4C08280",
-32067 => x"C0C0BFB0A4C082F8",
-32066 => x"C0C0BFB0A4C08282",
-32065 => x"C0C0BFB0A4C08292",
-32064 => x"C0C0BFB0A4C08299",
-32063 => x"C0C0BFB0A4C082B0",
-32062 => x"C0C0BFB0A4C082A4",
-32061 => x"C0C0BFB0A4C082F9",
-32060 => x"C0C0BFB0A4C082C0",
-32059 => x"C0C0BFB0A4C09290",
-32058 => x"C0C0BFB0A4C09280",
-32057 => x"C0C0BFB0A4C092F8",
-32056 => x"C0C0BFB0A4C09282",
-32055 => x"C0C0BFB0A4C09292",
-32054 => x"C0C0BFB0A4C09299",
-32053 => x"C0C0BFB0A4C092B0",
-32052 => x"C0C0BFB0A4C092A4",
-32051 => x"C0C0BFB0A4C092F9",
-32050 => x"C0C0BFB0A4C092C0",
-32049 => x"C0C0BFB0A4C09990",
-32048 => x"C0C0BFB0A4C09980",
-32047 => x"C0C0BFB0A4C099F8",
-32046 => x"C0C0BFB0A4C09982",
-32045 => x"C0C0BFB0A4C09992",
-32044 => x"C0C0BFB0A4C09999",
-32043 => x"C0C0BFB0A4C099B0",
-32042 => x"C0C0BFB0A4C099A4",
-32041 => x"C0C0BFB0A4C099F9",
-32040 => x"C0C0BFB0A4C099C0",
-32039 => x"C0C0BFB0A4C0B090",
-32038 => x"C0C0BFB0A4C0B080",
-32037 => x"C0C0BFB0A4C0B0F8",
-32036 => x"C0C0BFB0A4C0B082",
-32035 => x"C0C0BFB0A4C0B092",
-32034 => x"C0C0BFB0A4C0B099",
-32033 => x"C0C0BFB0A4C0B0B0",
-32032 => x"C0C0BFB0A4C0B0A4",
-32031 => x"C0C0BFB0A4C0B0F9",
-32030 => x"C0C0BFB0A4C0B0C0",
-32029 => x"C0C0BFB0A4C0A490",
-32028 => x"C0C0BFB0A4C0A480",
-32027 => x"C0C0BFB0A4C0A4F8",
-32026 => x"C0C0BFB0A4C0A482",
-32025 => x"C0C0BFB0A4C0A492",
-32024 => x"C0C0BFB0A4C0A499",
-32023 => x"C0C0BFB0A4C0A4B0",
-32022 => x"C0C0BFB0A4C0A4A4",
-32021 => x"C0C0BFB0A4C0A4F9",
-32020 => x"C0C0BFB0A4C0A4C0",
-32019 => x"C0C0BFB0A4C0F990",
-32018 => x"C0C0BFB0A4C0F980",
-32017 => x"C0C0BFB0A4C0F9F8",
-32016 => x"C0C0BFB0A4C0F982",
-32015 => x"C0C0BFB0A4C0F992",
-32014 => x"C0C0BFB0A4C0F999",
-32013 => x"C0C0BFB0A4C0F9B0",
-32012 => x"C0C0BFB0A4C0F9A4",
-32011 => x"C0C0BFB0A4C0F9F9",
-32010 => x"C0C0BFB0A4C0F9C0",
-32009 => x"C0C0BFB0A4C0C090",
-32008 => x"C0C0BFB0A4C0C080",
-32007 => x"C0C0BFB0A4C0C0F8",
-32006 => x"C0C0BFB0A4C0C082",
-32005 => x"C0C0BFB0A4C0C092",
-32004 => x"C0C0BFB0A4C0C099",
-32003 => x"C0C0BFB0A4C0C0B0",
-32002 => x"C0C0BFB0A4C0C0A4",
-32001 => x"C0C0BFB0A4C0C0F9",
-32000 => x"C0C0BFB0A4C0C0C0",
-31999 => x"C0C0BFB0F9909090",
-31998 => x"C0C0BFB0F9909080",
-31997 => x"C0C0BFB0F99090F8",
-31996 => x"C0C0BFB0F9909082",
-31995 => x"C0C0BFB0F9909092",
-31994 => x"C0C0BFB0F9909099",
-31993 => x"C0C0BFB0F99090B0",
-31992 => x"C0C0BFB0F99090A4",
-31991 => x"C0C0BFB0F99090F9",
-31990 => x"C0C0BFB0F99090C0",
-31989 => x"C0C0BFB0F9908090",
-31988 => x"C0C0BFB0F9908080",
-31987 => x"C0C0BFB0F99080F8",
-31986 => x"C0C0BFB0F9908082",
-31985 => x"C0C0BFB0F9908092",
-31984 => x"C0C0BFB0F9908099",
-31983 => x"C0C0BFB0F99080B0",
-31982 => x"C0C0BFB0F99080A4",
-31981 => x"C0C0BFB0F99080F9",
-31980 => x"C0C0BFB0F99080C0",
-31979 => x"C0C0BFB0F990F890",
-31978 => x"C0C0BFB0F990F880",
-31977 => x"C0C0BFB0F990F8F8",
-31976 => x"C0C0BFB0F990F882",
-31975 => x"C0C0BFB0F990F892",
-31974 => x"C0C0BFB0F990F899",
-31973 => x"C0C0BFB0F990F8B0",
-31972 => x"C0C0BFB0F990F8A4",
-31971 => x"C0C0BFB0F990F8F9",
-31970 => x"C0C0BFB0F990F8C0",
-31969 => x"C0C0BFB0F9908290",
-31968 => x"C0C0BFB0F9908280",
-31967 => x"C0C0BFB0F99082F8",
-31966 => x"C0C0BFB0F9908282",
-31965 => x"C0C0BFB0F9908292",
-31964 => x"C0C0BFB0F9908299",
-31963 => x"C0C0BFB0F99082B0",
-31962 => x"C0C0BFB0F99082A4",
-31961 => x"C0C0BFB0F99082F9",
-31960 => x"C0C0BFB0F99082C0",
-31959 => x"C0C0BFB0F9909290",
-31958 => x"C0C0BFB0F9909280",
-31957 => x"C0C0BFB0F99092F8",
-31956 => x"C0C0BFB0F9909282",
-31955 => x"C0C0BFB0F9909292",
-31954 => x"C0C0BFB0F9909299",
-31953 => x"C0C0BFB0F99092B0",
-31952 => x"C0C0BFB0F99092A4",
-31951 => x"C0C0BFB0F99092F9",
-31950 => x"C0C0BFB0F99092C0",
-31949 => x"C0C0BFB0F9909990",
-31948 => x"C0C0BFB0F9909980",
-31947 => x"C0C0BFB0F99099F8",
-31946 => x"C0C0BFB0F9909982",
-31945 => x"C0C0BFB0F9909992",
-31944 => x"C0C0BFB0F9909999",
-31943 => x"C0C0BFB0F99099B0",
-31942 => x"C0C0BFB0F99099A4",
-31941 => x"C0C0BFB0F99099F9",
-31940 => x"C0C0BFB0F99099C0",
-31939 => x"C0C0BFB0F990B090",
-31938 => x"C0C0BFB0F990B080",
-31937 => x"C0C0BFB0F990B0F8",
-31936 => x"C0C0BFB0F990B082",
-31935 => x"C0C0BFB0F990B092",
-31934 => x"C0C0BFB0F990B099",
-31933 => x"C0C0BFB0F990B0B0",
-31932 => x"C0C0BFB0F990B0A4",
-31931 => x"C0C0BFB0F990B0F9",
-31930 => x"C0C0BFB0F990B0C0",
-31929 => x"C0C0BFB0F990A490",
-31928 => x"C0C0BFB0F990A480",
-31927 => x"C0C0BFB0F990A4F8",
-31926 => x"C0C0BFB0F990A482",
-31925 => x"C0C0BFB0F990A492",
-31924 => x"C0C0BFB0F990A499",
-31923 => x"C0C0BFB0F990A4B0",
-31922 => x"C0C0BFB0F990A4A4",
-31921 => x"C0C0BFB0F990A4F9",
-31920 => x"C0C0BFB0F990A4C0",
-31919 => x"C0C0BFB0F990F990",
-31918 => x"C0C0BFB0F990F980",
-31917 => x"C0C0BFB0F990F9F8",
-31916 => x"C0C0BFB0F990F982",
-31915 => x"C0C0BFB0F990F992",
-31914 => x"C0C0BFB0F990F999",
-31913 => x"C0C0BFB0F990F9B0",
-31912 => x"C0C0BFB0F990F9A4",
-31911 => x"C0C0BFB0F990F9F9",
-31910 => x"C0C0BFB0F990F9C0",
-31909 => x"C0C0BFB0F990C090",
-31908 => x"C0C0BFB0F990C080",
-31907 => x"C0C0BFB0F990C0F8",
-31906 => x"C0C0BFB0F990C082",
-31905 => x"C0C0BFB0F990C092",
-31904 => x"C0C0BFB0F990C099",
-31903 => x"C0C0BFB0F990C0B0",
-31902 => x"C0C0BFB0F990C0A4",
-31901 => x"C0C0BFB0F990C0F9",
-31900 => x"C0C0BFB0F990C0C0",
-31899 => x"C0C0BFB0F9809090",
-31898 => x"C0C0BFB0F9809080",
-31897 => x"C0C0BFB0F98090F8",
-31896 => x"C0C0BFB0F9809082",
-31895 => x"C0C0BFB0F9809092",
-31894 => x"C0C0BFB0F9809099",
-31893 => x"C0C0BFB0F98090B0",
-31892 => x"C0C0BFB0F98090A4",
-31891 => x"C0C0BFB0F98090F9",
-31890 => x"C0C0BFB0F98090C0",
-31889 => x"C0C0BFB0F9808090",
-31888 => x"C0C0BFB0F9808080",
-31887 => x"C0C0BFB0F98080F8",
-31886 => x"C0C0BFB0F9808082",
-31885 => x"C0C0BFB0F9808092",
-31884 => x"C0C0BFB0F9808099",
-31883 => x"C0C0BFB0F98080B0",
-31882 => x"C0C0BFB0F98080A4",
-31881 => x"C0C0BFB0F98080F9",
-31880 => x"C0C0BFB0F98080C0",
-31879 => x"C0C0BFB0F980F890",
-31878 => x"C0C0BFB0F980F880",
-31877 => x"C0C0BFB0F980F8F8",
-31876 => x"C0C0BFB0F980F882",
-31875 => x"C0C0BFB0F980F892",
-31874 => x"C0C0BFB0F980F899",
-31873 => x"C0C0BFB0F980F8B0",
-31872 => x"C0C0BFB0F980F8A4",
-31871 => x"C0C0BFB0F980F8F9",
-31870 => x"C0C0BFB0F980F8C0",
-31869 => x"C0C0BFB0F9808290",
-31868 => x"C0C0BFB0F9808280",
-31867 => x"C0C0BFB0F98082F8",
-31866 => x"C0C0BFB0F9808282",
-31865 => x"C0C0BFB0F9808292",
-31864 => x"C0C0BFB0F9808299",
-31863 => x"C0C0BFB0F98082B0",
-31862 => x"C0C0BFB0F98082A4",
-31861 => x"C0C0BFB0F98082F9",
-31860 => x"C0C0BFB0F98082C0",
-31859 => x"C0C0BFB0F9809290",
-31858 => x"C0C0BFB0F9809280",
-31857 => x"C0C0BFB0F98092F8",
-31856 => x"C0C0BFB0F9809282",
-31855 => x"C0C0BFB0F9809292",
-31854 => x"C0C0BFB0F9809299",
-31853 => x"C0C0BFB0F98092B0",
-31852 => x"C0C0BFB0F98092A4",
-31851 => x"C0C0BFB0F98092F9",
-31850 => x"C0C0BFB0F98092C0",
-31849 => x"C0C0BFB0F9809990",
-31848 => x"C0C0BFB0F9809980",
-31847 => x"C0C0BFB0F98099F8",
-31846 => x"C0C0BFB0F9809982",
-31845 => x"C0C0BFB0F9809992",
-31844 => x"C0C0BFB0F9809999",
-31843 => x"C0C0BFB0F98099B0",
-31842 => x"C0C0BFB0F98099A4",
-31841 => x"C0C0BFB0F98099F9",
-31840 => x"C0C0BFB0F98099C0",
-31839 => x"C0C0BFB0F980B090",
-31838 => x"C0C0BFB0F980B080",
-31837 => x"C0C0BFB0F980B0F8",
-31836 => x"C0C0BFB0F980B082",
-31835 => x"C0C0BFB0F980B092",
-31834 => x"C0C0BFB0F980B099",
-31833 => x"C0C0BFB0F980B0B0",
-31832 => x"C0C0BFB0F980B0A4",
-31831 => x"C0C0BFB0F980B0F9",
-31830 => x"C0C0BFB0F980B0C0",
-31829 => x"C0C0BFB0F980A490",
-31828 => x"C0C0BFB0F980A480",
-31827 => x"C0C0BFB0F980A4F8",
-31826 => x"C0C0BFB0F980A482",
-31825 => x"C0C0BFB0F980A492",
-31824 => x"C0C0BFB0F980A499",
-31823 => x"C0C0BFB0F980A4B0",
-31822 => x"C0C0BFB0F980A4A4",
-31821 => x"C0C0BFB0F980A4F9",
-31820 => x"C0C0BFB0F980A4C0",
-31819 => x"C0C0BFB0F980F990",
-31818 => x"C0C0BFB0F980F980",
-31817 => x"C0C0BFB0F980F9F8",
-31816 => x"C0C0BFB0F980F982",
-31815 => x"C0C0BFB0F980F992",
-31814 => x"C0C0BFB0F980F999",
-31813 => x"C0C0BFB0F980F9B0",
-31812 => x"C0C0BFB0F980F9A4",
-31811 => x"C0C0BFB0F980F9F9",
-31810 => x"C0C0BFB0F980F9C0",
-31809 => x"C0C0BFB0F980C090",
-31808 => x"C0C0BFB0F980C080",
-31807 => x"C0C0BFB0F980C0F8",
-31806 => x"C0C0BFB0F980C082",
-31805 => x"C0C0BFB0F980C092",
-31804 => x"C0C0BFB0F980C099",
-31803 => x"C0C0BFB0F980C0B0",
-31802 => x"C0C0BFB0F980C0A4",
-31801 => x"C0C0BFB0F980C0F9",
-31800 => x"C0C0BFB0F980C0C0",
-31799 => x"C0C0BFB0F9F89090",
-31798 => x"C0C0BFB0F9F89080",
-31797 => x"C0C0BFB0F9F890F8",
-31796 => x"C0C0BFB0F9F89082",
-31795 => x"C0C0BFB0F9F89092",
-31794 => x"C0C0BFB0F9F89099",
-31793 => x"C0C0BFB0F9F890B0",
-31792 => x"C0C0BFB0F9F890A4",
-31791 => x"C0C0BFB0F9F890F9",
-31790 => x"C0C0BFB0F9F890C0",
-31789 => x"C0C0BFB0F9F88090",
-31788 => x"C0C0BFB0F9F88080",
-31787 => x"C0C0BFB0F9F880F8",
-31786 => x"C0C0BFB0F9F88082",
-31785 => x"C0C0BFB0F9F88092",
-31784 => x"C0C0BFB0F9F88099",
-31783 => x"C0C0BFB0F9F880B0",
-31782 => x"C0C0BFB0F9F880A4",
-31781 => x"C0C0BFB0F9F880F9",
-31780 => x"C0C0BFB0F9F880C0",
-31779 => x"C0C0BFB0F9F8F890",
-31778 => x"C0C0BFB0F9F8F880",
-31777 => x"C0C0BFB0F9F8F8F8",
-31776 => x"C0C0BFB0F9F8F882",
-31775 => x"C0C0BFB0F9F8F892",
-31774 => x"C0C0BFB0F9F8F899",
-31773 => x"C0C0BFB0F9F8F8B0",
-31772 => x"C0C0BFB0F9F8F8A4",
-31771 => x"C0C0BFB0F9F8F8F9",
-31770 => x"C0C0BFB0F9F8F8C0",
-31769 => x"C0C0BFB0F9F88290",
-31768 => x"C0C0BFB0F9F88280",
-31767 => x"C0C0BFB0F9F882F8",
-31766 => x"C0C0BFB0F9F88282",
-31765 => x"C0C0BFB0F9F88292",
-31764 => x"C0C0BFB0F9F88299",
-31763 => x"C0C0BFB0F9F882B0",
-31762 => x"C0C0BFB0F9F882A4",
-31761 => x"C0C0BFB0F9F882F9",
-31760 => x"C0C0BFB0F9F882C0",
-31759 => x"C0C0BFB0F9F89290",
-31758 => x"C0C0BFB0F9F89280",
-31757 => x"C0C0BFB0F9F892F8",
-31756 => x"C0C0BFB0F9F89282",
-31755 => x"C0C0BFB0F9F89292",
-31754 => x"C0C0BFB0F9F89299",
-31753 => x"C0C0BFB0F9F892B0",
-31752 => x"C0C0BFB0F9F892A4",
-31751 => x"C0C0BFB0F9F892F9",
-31750 => x"C0C0BFB0F9F892C0",
-31749 => x"C0C0BFB0F9F89990",
-31748 => x"C0C0BFB0F9F89980",
-31747 => x"C0C0BFB0F9F899F8",
-31746 => x"C0C0BFB0F9F89982",
-31745 => x"C0C0BFB0F9F89992",
-31744 => x"C0C0BFB0F9F89999",
-31743 => x"C0C0BFB0F9F899B0",
-31742 => x"C0C0BFB0F9F899A4",
-31741 => x"C0C0BFB0F9F899F9",
-31740 => x"C0C0BFB0F9F899C0",
-31739 => x"C0C0BFB0F9F8B090",
-31738 => x"C0C0BFB0F9F8B080",
-31737 => x"C0C0BFB0F9F8B0F8",
-31736 => x"C0C0BFB0F9F8B082",
-31735 => x"C0C0BFB0F9F8B092",
-31734 => x"C0C0BFB0F9F8B099",
-31733 => x"C0C0BFB0F9F8B0B0",
-31732 => x"C0C0BFB0F9F8B0A4",
-31731 => x"C0C0BFB0F9F8B0F9",
-31730 => x"C0C0BFB0F9F8B0C0",
-31729 => x"C0C0BFB0F9F8A490",
-31728 => x"C0C0BFB0F9F8A480",
-31727 => x"C0C0BFB0F9F8A4F8",
-31726 => x"C0C0BFB0F9F8A482",
-31725 => x"C0C0BFB0F9F8A492",
-31724 => x"C0C0BFB0F9F8A499",
-31723 => x"C0C0BFB0F9F8A4B0",
-31722 => x"C0C0BFB0F9F8A4A4",
-31721 => x"C0C0BFB0F9F8A4F9",
-31720 => x"C0C0BFB0F9F8A4C0",
-31719 => x"C0C0BFB0F9F8F990",
-31718 => x"C0C0BFB0F9F8F980",
-31717 => x"C0C0BFB0F9F8F9F8",
-31716 => x"C0C0BFB0F9F8F982",
-31715 => x"C0C0BFB0F9F8F992",
-31714 => x"C0C0BFB0F9F8F999",
-31713 => x"C0C0BFB0F9F8F9B0",
-31712 => x"C0C0BFB0F9F8F9A4",
-31711 => x"C0C0BFB0F9F8F9F9",
-31710 => x"C0C0BFB0F9F8F9C0",
-31709 => x"C0C0BFB0F9F8C090",
-31708 => x"C0C0BFB0F9F8C080",
-31707 => x"C0C0BFB0F9F8C0F8",
-31706 => x"C0C0BFB0F9F8C082",
-31705 => x"C0C0BFB0F9F8C092",
-31704 => x"C0C0BFB0F9F8C099",
-31703 => x"C0C0BFB0F9F8C0B0",
-31702 => x"C0C0BFB0F9F8C0A4",
-31701 => x"C0C0BFB0F9F8C0F9",
-31700 => x"C0C0BFB0F9F8C0C0",
-31699 => x"C0C0BFB0F9829090",
-31698 => x"C0C0BFB0F9829080",
-31697 => x"C0C0BFB0F98290F8",
-31696 => x"C0C0BFB0F9829082",
-31695 => x"C0C0BFB0F9829092",
-31694 => x"C0C0BFB0F9829099",
-31693 => x"C0C0BFB0F98290B0",
-31692 => x"C0C0BFB0F98290A4",
-31691 => x"C0C0BFB0F98290F9",
-31690 => x"C0C0BFB0F98290C0",
-31689 => x"C0C0BFB0F9828090",
-31688 => x"C0C0BFB0F9828080",
-31687 => x"C0C0BFB0F98280F8",
-31686 => x"C0C0BFB0F9828082",
-31685 => x"C0C0BFB0F9828092",
-31684 => x"C0C0BFB0F9828099",
-31683 => x"C0C0BFB0F98280B0",
-31682 => x"C0C0BFB0F98280A4",
-31681 => x"C0C0BFB0F98280F9",
-31680 => x"C0C0BFB0F98280C0",
-31679 => x"C0C0BFB0F982F890",
-31678 => x"C0C0BFB0F982F880",
-31677 => x"C0C0BFB0F982F8F8",
-31676 => x"C0C0BFB0F982F882",
-31675 => x"C0C0BFB0F982F892",
-31674 => x"C0C0BFB0F982F899",
-31673 => x"C0C0BFB0F982F8B0",
-31672 => x"C0C0BFB0F982F8A4",
-31671 => x"C0C0BFB0F982F8F9",
-31670 => x"C0C0BFB0F982F8C0",
-31669 => x"C0C0BFB0F9828290",
-31668 => x"C0C0BFB0F9828280",
-31667 => x"C0C0BFB0F98282F8",
-31666 => x"C0C0BFB0F9828282",
-31665 => x"C0C0BFB0F9828292",
-31664 => x"C0C0BFB0F9828299",
-31663 => x"C0C0BFB0F98282B0",
-31662 => x"C0C0BFB0F98282A4",
-31661 => x"C0C0BFB0F98282F9",
-31660 => x"C0C0BFB0F98282C0",
-31659 => x"C0C0BFB0F9829290",
-31658 => x"C0C0BFB0F9829280",
-31657 => x"C0C0BFB0F98292F8",
-31656 => x"C0C0BFB0F9829282",
-31655 => x"C0C0BFB0F9829292",
-31654 => x"C0C0BFB0F9829299",
-31653 => x"C0C0BFB0F98292B0",
-31652 => x"C0C0BFB0F98292A4",
-31651 => x"C0C0BFB0F98292F9",
-31650 => x"C0C0BFB0F98292C0",
-31649 => x"C0C0BFB0F9829990",
-31648 => x"C0C0BFB0F9829980",
-31647 => x"C0C0BFB0F98299F8",
-31646 => x"C0C0BFB0F9829982",
-31645 => x"C0C0BFB0F9829992",
-31644 => x"C0C0BFB0F9829999",
-31643 => x"C0C0BFB0F98299B0",
-31642 => x"C0C0BFB0F98299A4",
-31641 => x"C0C0BFB0F98299F9",
-31640 => x"C0C0BFB0F98299C0",
-31639 => x"C0C0BFB0F982B090",
-31638 => x"C0C0BFB0F982B080",
-31637 => x"C0C0BFB0F982B0F8",
-31636 => x"C0C0BFB0F982B082",
-31635 => x"C0C0BFB0F982B092",
-31634 => x"C0C0BFB0F982B099",
-31633 => x"C0C0BFB0F982B0B0",
-31632 => x"C0C0BFB0F982B0A4",
-31631 => x"C0C0BFB0F982B0F9",
-31630 => x"C0C0BFB0F982B0C0",
-31629 => x"C0C0BFB0F982A490",
-31628 => x"C0C0BFB0F982A480",
-31627 => x"C0C0BFB0F982A4F8",
-31626 => x"C0C0BFB0F982A482",
-31625 => x"C0C0BFB0F982A492",
-31624 => x"C0C0BFB0F982A499",
-31623 => x"C0C0BFB0F982A4B0",
-31622 => x"C0C0BFB0F982A4A4",
-31621 => x"C0C0BFB0F982A4F9",
-31620 => x"C0C0BFB0F982A4C0",
-31619 => x"C0C0BFB0F982F990",
-31618 => x"C0C0BFB0F982F980",
-31617 => x"C0C0BFB0F982F9F8",
-31616 => x"C0C0BFB0F982F982",
-31615 => x"C0C0BFB0F982F992",
-31614 => x"C0C0BFB0F982F999",
-31613 => x"C0C0BFB0F982F9B0",
-31612 => x"C0C0BFB0F982F9A4",
-31611 => x"C0C0BFB0F982F9F9",
-31610 => x"C0C0BFB0F982F9C0",
-31609 => x"C0C0BFB0F982C090",
-31608 => x"C0C0BFB0F982C080",
-31607 => x"C0C0BFB0F982C0F8",
-31606 => x"C0C0BFB0F982C082",
-31605 => x"C0C0BFB0F982C092",
-31604 => x"C0C0BFB0F982C099",
-31603 => x"C0C0BFB0F982C0B0",
-31602 => x"C0C0BFB0F982C0A4",
-31601 => x"C0C0BFB0F982C0F9",
-31600 => x"C0C0BFB0F982C0C0",
-31599 => x"C0C0BFB0F9929090",
-31598 => x"C0C0BFB0F9929080",
-31597 => x"C0C0BFB0F99290F8",
-31596 => x"C0C0BFB0F9929082",
-31595 => x"C0C0BFB0F9929092",
-31594 => x"C0C0BFB0F9929099",
-31593 => x"C0C0BFB0F99290B0",
-31592 => x"C0C0BFB0F99290A4",
-31591 => x"C0C0BFB0F99290F9",
-31590 => x"C0C0BFB0F99290C0",
-31589 => x"C0C0BFB0F9928090",
-31588 => x"C0C0BFB0F9928080",
-31587 => x"C0C0BFB0F99280F8",
-31586 => x"C0C0BFB0F9928082",
-31585 => x"C0C0BFB0F9928092",
-31584 => x"C0C0BFB0F9928099",
-31583 => x"C0C0BFB0F99280B0",
-31582 => x"C0C0BFB0F99280A4",
-31581 => x"C0C0BFB0F99280F9",
-31580 => x"C0C0BFB0F99280C0",
-31579 => x"C0C0BFB0F992F890",
-31578 => x"C0C0BFB0F992F880",
-31577 => x"C0C0BFB0F992F8F8",
-31576 => x"C0C0BFB0F992F882",
-31575 => x"C0C0BFB0F992F892",
-31574 => x"C0C0BFB0F992F899",
-31573 => x"C0C0BFB0F992F8B0",
-31572 => x"C0C0BFB0F992F8A4",
-31571 => x"C0C0BFB0F992F8F9",
-31570 => x"C0C0BFB0F992F8C0",
-31569 => x"C0C0BFB0F9928290",
-31568 => x"C0C0BFB0F9928280",
-31567 => x"C0C0BFB0F99282F8",
-31566 => x"C0C0BFB0F9928282",
-31565 => x"C0C0BFB0F9928292",
-31564 => x"C0C0BFB0F9928299",
-31563 => x"C0C0BFB0F99282B0",
-31562 => x"C0C0BFB0F99282A4",
-31561 => x"C0C0BFB0F99282F9",
-31560 => x"C0C0BFB0F99282C0",
-31559 => x"C0C0BFB0F9929290",
-31558 => x"C0C0BFB0F9929280",
-31557 => x"C0C0BFB0F99292F8",
-31556 => x"C0C0BFB0F9929282",
-31555 => x"C0C0BFB0F9929292",
-31554 => x"C0C0BFB0F9929299",
-31553 => x"C0C0BFB0F99292B0",
-31552 => x"C0C0BFB0F99292A4",
-31551 => x"C0C0BFB0F99292F9",
-31550 => x"C0C0BFB0F99292C0",
-31549 => x"C0C0BFB0F9929990",
-31548 => x"C0C0BFB0F9929980",
-31547 => x"C0C0BFB0F99299F8",
-31546 => x"C0C0BFB0F9929982",
-31545 => x"C0C0BFB0F9929992",
-31544 => x"C0C0BFB0F9929999",
-31543 => x"C0C0BFB0F99299B0",
-31542 => x"C0C0BFB0F99299A4",
-31541 => x"C0C0BFB0F99299F9",
-31540 => x"C0C0BFB0F99299C0",
-31539 => x"C0C0BFB0F992B090",
-31538 => x"C0C0BFB0F992B080",
-31537 => x"C0C0BFB0F992B0F8",
-31536 => x"C0C0BFB0F992B082",
-31535 => x"C0C0BFB0F992B092",
-31534 => x"C0C0BFB0F992B099",
-31533 => x"C0C0BFB0F992B0B0",
-31532 => x"C0C0BFB0F992B0A4",
-31531 => x"C0C0BFB0F992B0F9",
-31530 => x"C0C0BFB0F992B0C0",
-31529 => x"C0C0BFB0F992A490",
-31528 => x"C0C0BFB0F992A480",
-31527 => x"C0C0BFB0F992A4F8",
-31526 => x"C0C0BFB0F992A482",
-31525 => x"C0C0BFB0F992A492",
-31524 => x"C0C0BFB0F992A499",
-31523 => x"C0C0BFB0F992A4B0",
-31522 => x"C0C0BFB0F992A4A4",
-31521 => x"C0C0BFB0F992A4F9",
-31520 => x"C0C0BFB0F992A4C0",
-31519 => x"C0C0BFB0F992F990",
-31518 => x"C0C0BFB0F992F980",
-31517 => x"C0C0BFB0F992F9F8",
-31516 => x"C0C0BFB0F992F982",
-31515 => x"C0C0BFB0F992F992",
-31514 => x"C0C0BFB0F992F999",
-31513 => x"C0C0BFB0F992F9B0",
-31512 => x"C0C0BFB0F992F9A4",
-31511 => x"C0C0BFB0F992F9F9",
-31510 => x"C0C0BFB0F992F9C0",
-31509 => x"C0C0BFB0F992C090",
-31508 => x"C0C0BFB0F992C080",
-31507 => x"C0C0BFB0F992C0F8",
-31506 => x"C0C0BFB0F992C082",
-31505 => x"C0C0BFB0F992C092",
-31504 => x"C0C0BFB0F992C099",
-31503 => x"C0C0BFB0F992C0B0",
-31502 => x"C0C0BFB0F992C0A4",
-31501 => x"C0C0BFB0F992C0F9",
-31500 => x"C0C0BFB0F992C0C0",
-31499 => x"C0C0BFB0F9999090",
-31498 => x"C0C0BFB0F9999080",
-31497 => x"C0C0BFB0F99990F8",
-31496 => x"C0C0BFB0F9999082",
-31495 => x"C0C0BFB0F9999092",
-31494 => x"C0C0BFB0F9999099",
-31493 => x"C0C0BFB0F99990B0",
-31492 => x"C0C0BFB0F99990A4",
-31491 => x"C0C0BFB0F99990F9",
-31490 => x"C0C0BFB0F99990C0",
-31489 => x"C0C0BFB0F9998090",
-31488 => x"C0C0BFB0F9998080",
-31487 => x"C0C0BFB0F99980F8",
-31486 => x"C0C0BFB0F9998082",
-31485 => x"C0C0BFB0F9998092",
-31484 => x"C0C0BFB0F9998099",
-31483 => x"C0C0BFB0F99980B0",
-31482 => x"C0C0BFB0F99980A4",
-31481 => x"C0C0BFB0F99980F9",
-31480 => x"C0C0BFB0F99980C0",
-31479 => x"C0C0BFB0F999F890",
-31478 => x"C0C0BFB0F999F880",
-31477 => x"C0C0BFB0F999F8F8",
-31476 => x"C0C0BFB0F999F882",
-31475 => x"C0C0BFB0F999F892",
-31474 => x"C0C0BFB0F999F899",
-31473 => x"C0C0BFB0F999F8B0",
-31472 => x"C0C0BFB0F999F8A4",
-31471 => x"C0C0BFB0F999F8F9",
-31470 => x"C0C0BFB0F999F8C0",
-31469 => x"C0C0BFB0F9998290",
-31468 => x"C0C0BFB0F9998280",
-31467 => x"C0C0BFB0F99982F8",
-31466 => x"C0C0BFB0F9998282",
-31465 => x"C0C0BFB0F9998292",
-31464 => x"C0C0BFB0F9998299",
-31463 => x"C0C0BFB0F99982B0",
-31462 => x"C0C0BFB0F99982A4",
-31461 => x"C0C0BFB0F99982F9",
-31460 => x"C0C0BFB0F99982C0",
-31459 => x"C0C0BFB0F9999290",
-31458 => x"C0C0BFB0F9999280",
-31457 => x"C0C0BFB0F99992F8",
-31456 => x"C0C0BFB0F9999282",
-31455 => x"C0C0BFB0F9999292",
-31454 => x"C0C0BFB0F9999299",
-31453 => x"C0C0BFB0F99992B0",
-31452 => x"C0C0BFB0F99992A4",
-31451 => x"C0C0BFB0F99992F9",
-31450 => x"C0C0BFB0F99992C0",
-31449 => x"C0C0BFB0F9999990",
-31448 => x"C0C0BFB0F9999980",
-31447 => x"C0C0BFB0F99999F8",
-31446 => x"C0C0BFB0F9999982",
-31445 => x"C0C0BFB0F9999992",
-31444 => x"C0C0BFB0F9999999",
-31443 => x"C0C0BFB0F99999B0",
-31442 => x"C0C0BFB0F99999A4",
-31441 => x"C0C0BFB0F99999F9",
-31440 => x"C0C0BFB0F99999C0",
-31439 => x"C0C0BFB0F999B090",
-31438 => x"C0C0BFB0F999B080",
-31437 => x"C0C0BFB0F999B0F8",
-31436 => x"C0C0BFB0F999B082",
-31435 => x"C0C0BFB0F999B092",
-31434 => x"C0C0BFB0F999B099",
-31433 => x"C0C0BFB0F999B0B0",
-31432 => x"C0C0BFB0F999B0A4",
-31431 => x"C0C0BFB0F999B0F9",
-31430 => x"C0C0BFB0F999B0C0",
-31429 => x"C0C0BFB0F999A490",
-31428 => x"C0C0BFB0F999A480",
-31427 => x"C0C0BFB0F999A4F8",
-31426 => x"C0C0BFB0F999A482",
-31425 => x"C0C0BFB0F999A492",
-31424 => x"C0C0BFB0F999A499",
-31423 => x"C0C0BFB0F999A4B0",
-31422 => x"C0C0BFB0F999A4A4",
-31421 => x"C0C0BFB0F999A4F9",
-31420 => x"C0C0BFB0F999A4C0",
-31419 => x"C0C0BFB0F999F990",
-31418 => x"C0C0BFB0F999F980",
-31417 => x"C0C0BFB0F999F9F8",
-31416 => x"C0C0BFB0F999F982",
-31415 => x"C0C0BFB0F999F992",
-31414 => x"C0C0BFB0F999F999",
-31413 => x"C0C0BFB0F999F9B0",
-31412 => x"C0C0BFB0F999F9A4",
-31411 => x"C0C0BFB0F999F9F9",
-31410 => x"C0C0BFB0F999F9C0",
-31409 => x"C0C0BFB0F999C090",
-31408 => x"C0C0BFB0F999C080",
-31407 => x"C0C0BFB0F999C0F8",
-31406 => x"C0C0BFB0F999C082",
-31405 => x"C0C0BFB0F999C092",
-31404 => x"C0C0BFB0F999C099",
-31403 => x"C0C0BFB0F999C0B0",
-31402 => x"C0C0BFB0F999C0A4",
-31401 => x"C0C0BFB0F999C0F9",
-31400 => x"C0C0BFB0F999C0C0",
-31399 => x"C0C0BFB0F9B09090",
-31398 => x"C0C0BFB0F9B09080",
-31397 => x"C0C0BFB0F9B090F8",
-31396 => x"C0C0BFB0F9B09082",
-31395 => x"C0C0BFB0F9B09092",
-31394 => x"C0C0BFB0F9B09099",
-31393 => x"C0C0BFB0F9B090B0",
-31392 => x"C0C0BFB0F9B090A4",
-31391 => x"C0C0BFB0F9B090F9",
-31390 => x"C0C0BFB0F9B090C0",
-31389 => x"C0C0BFB0F9B08090",
-31388 => x"C0C0BFB0F9B08080",
-31387 => x"C0C0BFB0F9B080F8",
-31386 => x"C0C0BFB0F9B08082",
-31385 => x"C0C0BFB0F9B08092",
-31384 => x"C0C0BFB0F9B08099",
-31383 => x"C0C0BFB0F9B080B0",
-31382 => x"C0C0BFB0F9B080A4",
-31381 => x"C0C0BFB0F9B080F9",
-31380 => x"C0C0BFB0F9B080C0",
-31379 => x"C0C0BFB0F9B0F890",
-31378 => x"C0C0BFB0F9B0F880",
-31377 => x"C0C0BFB0F9B0F8F8",
-31376 => x"C0C0BFB0F9B0F882",
-31375 => x"C0C0BFB0F9B0F892",
-31374 => x"C0C0BFB0F9B0F899",
-31373 => x"C0C0BFB0F9B0F8B0",
-31372 => x"C0C0BFB0F9B0F8A4",
-31371 => x"C0C0BFB0F9B0F8F9",
-31370 => x"C0C0BFB0F9B0F8C0",
-31369 => x"C0C0BFB0F9B08290",
-31368 => x"C0C0BFB0F9B08280",
-31367 => x"C0C0BFB0F9B082F8",
-31366 => x"C0C0BFB0F9B08282",
-31365 => x"C0C0BFB0F9B08292",
-31364 => x"C0C0BFB0F9B08299",
-31363 => x"C0C0BFB0F9B082B0",
-31362 => x"C0C0BFB0F9B082A4",
-31361 => x"C0C0BFB0F9B082F9",
-31360 => x"C0C0BFB0F9B082C0",
-31359 => x"C0C0BFB0F9B09290",
-31358 => x"C0C0BFB0F9B09280",
-31357 => x"C0C0BFB0F9B092F8",
-31356 => x"C0C0BFB0F9B09282",
-31355 => x"C0C0BFB0F9B09292",
-31354 => x"C0C0BFB0F9B09299",
-31353 => x"C0C0BFB0F9B092B0",
-31352 => x"C0C0BFB0F9B092A4",
-31351 => x"C0C0BFB0F9B092F9",
-31350 => x"C0C0BFB0F9B092C0",
-31349 => x"C0C0BFB0F9B09990",
-31348 => x"C0C0BFB0F9B09980",
-31347 => x"C0C0BFB0F9B099F8",
-31346 => x"C0C0BFB0F9B09982",
-31345 => x"C0C0BFB0F9B09992",
-31344 => x"C0C0BFB0F9B09999",
-31343 => x"C0C0BFB0F9B099B0",
-31342 => x"C0C0BFB0F9B099A4",
-31341 => x"C0C0BFB0F9B099F9",
-31340 => x"C0C0BFB0F9B099C0",
-31339 => x"C0C0BFB0F9B0B090",
-31338 => x"C0C0BFB0F9B0B080",
-31337 => x"C0C0BFB0F9B0B0F8",
-31336 => x"C0C0BFB0F9B0B082",
-31335 => x"C0C0BFB0F9B0B092",
-31334 => x"C0C0BFB0F9B0B099",
-31333 => x"C0C0BFB0F9B0B0B0",
-31332 => x"C0C0BFB0F9B0B0A4",
-31331 => x"C0C0BFB0F9B0B0F9",
-31330 => x"C0C0BFB0F9B0B0C0",
-31329 => x"C0C0BFB0F9B0A490",
-31328 => x"C0C0BFB0F9B0A480",
-31327 => x"C0C0BFB0F9B0A4F8",
-31326 => x"C0C0BFB0F9B0A482",
-31325 => x"C0C0BFB0F9B0A492",
-31324 => x"C0C0BFB0F9B0A499",
-31323 => x"C0C0BFB0F9B0A4B0",
-31322 => x"C0C0BFB0F9B0A4A4",
-31321 => x"C0C0BFB0F9B0A4F9",
-31320 => x"C0C0BFB0F9B0A4C0",
-31319 => x"C0C0BFB0F9B0F990",
-31318 => x"C0C0BFB0F9B0F980",
-31317 => x"C0C0BFB0F9B0F9F8",
-31316 => x"C0C0BFB0F9B0F982",
-31315 => x"C0C0BFB0F9B0F992",
-31314 => x"C0C0BFB0F9B0F999",
-31313 => x"C0C0BFB0F9B0F9B0",
-31312 => x"C0C0BFB0F9B0F9A4",
-31311 => x"C0C0BFB0F9B0F9F9",
-31310 => x"C0C0BFB0F9B0F9C0",
-31309 => x"C0C0BFB0F9B0C090",
-31308 => x"C0C0BFB0F9B0C080",
-31307 => x"C0C0BFB0F9B0C0F8",
-31306 => x"C0C0BFB0F9B0C082",
-31305 => x"C0C0BFB0F9B0C092",
-31304 => x"C0C0BFB0F9B0C099",
-31303 => x"C0C0BFB0F9B0C0B0",
-31302 => x"C0C0BFB0F9B0C0A4",
-31301 => x"C0C0BFB0F9B0C0F9",
-31300 => x"C0C0BFB0F9B0C0C0",
-31299 => x"C0C0BFB0F9A49090",
-31298 => x"C0C0BFB0F9A49080",
-31297 => x"C0C0BFB0F9A490F8",
-31296 => x"C0C0BFB0F9A49082",
-31295 => x"C0C0BFB0F9A49092",
-31294 => x"C0C0BFB0F9A49099",
-31293 => x"C0C0BFB0F9A490B0",
-31292 => x"C0C0BFB0F9A490A4",
-31291 => x"C0C0BFB0F9A490F9",
-31290 => x"C0C0BFB0F9A490C0",
-31289 => x"C0C0BFB0F9A48090",
-31288 => x"C0C0BFB0F9A48080",
-31287 => x"C0C0BFB0F9A480F8",
-31286 => x"C0C0BFB0F9A48082",
-31285 => x"C0C0BFB0F9A48092",
-31284 => x"C0C0BFB0F9A48099",
-31283 => x"C0C0BFB0F9A480B0",
-31282 => x"C0C0BFB0F9A480A4",
-31281 => x"C0C0BFB0F9A480F9",
-31280 => x"C0C0BFB0F9A480C0",
-31279 => x"C0C0BFB0F9A4F890",
-31278 => x"C0C0BFB0F9A4F880",
-31277 => x"C0C0BFB0F9A4F8F8",
-31276 => x"C0C0BFB0F9A4F882",
-31275 => x"C0C0BFB0F9A4F892",
-31274 => x"C0C0BFB0F9A4F899",
-31273 => x"C0C0BFB0F9A4F8B0",
-31272 => x"C0C0BFB0F9A4F8A4",
-31271 => x"C0C0BFB0F9A4F8F9",
-31270 => x"C0C0BFB0F9A4F8C0",
-31269 => x"C0C0BFB0F9A48290",
-31268 => x"C0C0BFB0F9A48280",
-31267 => x"C0C0BFB0F9A482F8",
-31266 => x"C0C0BFB0F9A48282",
-31265 => x"C0C0BFB0F9A48292",
-31264 => x"C0C0BFB0F9A48299",
-31263 => x"C0C0BFB0F9A482B0",
-31262 => x"C0C0BFB0F9A482A4",
-31261 => x"C0C0BFB0F9A482F9",
-31260 => x"C0C0BFB0F9A482C0",
-31259 => x"C0C0BFB0F9A49290",
-31258 => x"C0C0BFB0F9A49280",
-31257 => x"C0C0BFB0F9A492F8",
-31256 => x"C0C0BFB0F9A49282",
-31255 => x"C0C0BFB0F9A49292",
-31254 => x"C0C0BFB0F9A49299",
-31253 => x"C0C0BFB0F9A492B0",
-31252 => x"C0C0BFB0F9A492A4",
-31251 => x"C0C0BFB0F9A492F9",
-31250 => x"C0C0BFB0F9A492C0",
-31249 => x"C0C0BFB0F9A49990",
-31248 => x"C0C0BFB0F9A49980",
-31247 => x"C0C0BFB0F9A499F8",
-31246 => x"C0C0BFB0F9A49982",
-31245 => x"C0C0BFB0F9A49992",
-31244 => x"C0C0BFB0F9A49999",
-31243 => x"C0C0BFB0F9A499B0",
-31242 => x"C0C0BFB0F9A499A4",
-31241 => x"C0C0BFB0F9A499F9",
-31240 => x"C0C0BFB0F9A499C0",
-31239 => x"C0C0BFB0F9A4B090",
-31238 => x"C0C0BFB0F9A4B080",
-31237 => x"C0C0BFB0F9A4B0F8",
-31236 => x"C0C0BFB0F9A4B082",
-31235 => x"C0C0BFB0F9A4B092",
-31234 => x"C0C0BFB0F9A4B099",
-31233 => x"C0C0BFB0F9A4B0B0",
-31232 => x"C0C0BFB0F9A4B0A4",
-31231 => x"C0C0BFB0F9A4B0F9",
-31230 => x"C0C0BFB0F9A4B0C0",
-31229 => x"C0C0BFB0F9A4A490",
-31228 => x"C0C0BFB0F9A4A480",
-31227 => x"C0C0BFB0F9A4A4F8",
-31226 => x"C0C0BFB0F9A4A482",
-31225 => x"C0C0BFB0F9A4A492",
-31224 => x"C0C0BFB0F9A4A499",
-31223 => x"C0C0BFB0F9A4A4B0",
-31222 => x"C0C0BFB0F9A4A4A4",
-31221 => x"C0C0BFB0F9A4A4F9",
-31220 => x"C0C0BFB0F9A4A4C0",
-31219 => x"C0C0BFB0F9A4F990",
-31218 => x"C0C0BFB0F9A4F980",
-31217 => x"C0C0BFB0F9A4F9F8",
-31216 => x"C0C0BFB0F9A4F982",
-31215 => x"C0C0BFB0F9A4F992",
-31214 => x"C0C0BFB0F9A4F999",
-31213 => x"C0C0BFB0F9A4F9B0",
-31212 => x"C0C0BFB0F9A4F9A4",
-31211 => x"C0C0BFB0F9A4F9F9",
-31210 => x"C0C0BFB0F9A4F9C0",
-31209 => x"C0C0BFB0F9A4C090",
-31208 => x"C0C0BFB0F9A4C080",
-31207 => x"C0C0BFB0F9A4C0F8",
-31206 => x"C0C0BFB0F9A4C082",
-31205 => x"C0C0BFB0F9A4C092",
-31204 => x"C0C0BFB0F9A4C099",
-31203 => x"C0C0BFB0F9A4C0B0",
-31202 => x"C0C0BFB0F9A4C0A4",
-31201 => x"C0C0BFB0F9A4C0F9",
-31200 => x"C0C0BFB0F9A4C0C0",
-31199 => x"C0C0BFB0F9F99090",
-31198 => x"C0C0BFB0F9F99080",
-31197 => x"C0C0BFB0F9F990F8",
-31196 => x"C0C0BFB0F9F99082",
-31195 => x"C0C0BFB0F9F99092",
-31194 => x"C0C0BFB0F9F99099",
-31193 => x"C0C0BFB0F9F990B0",
-31192 => x"C0C0BFB0F9F990A4",
-31191 => x"C0C0BFB0F9F990F9",
-31190 => x"C0C0BFB0F9F990C0",
-31189 => x"C0C0BFB0F9F98090",
-31188 => x"C0C0BFB0F9F98080",
-31187 => x"C0C0BFB0F9F980F8",
-31186 => x"C0C0BFB0F9F98082",
-31185 => x"C0C0BFB0F9F98092",
-31184 => x"C0C0BFB0F9F98099",
-31183 => x"C0C0BFB0F9F980B0",
-31182 => x"C0C0BFB0F9F980A4",
-31181 => x"C0C0BFB0F9F980F9",
-31180 => x"C0C0BFB0F9F980C0",
-31179 => x"C0C0BFB0F9F9F890",
-31178 => x"C0C0BFB0F9F9F880",
-31177 => x"C0C0BFB0F9F9F8F8",
-31176 => x"C0C0BFB0F9F9F882",
-31175 => x"C0C0BFB0F9F9F892",
-31174 => x"C0C0BFB0F9F9F899",
-31173 => x"C0C0BFB0F9F9F8B0",
-31172 => x"C0C0BFB0F9F9F8A4",
-31171 => x"C0C0BFB0F9F9F8F9",
-31170 => x"C0C0BFB0F9F9F8C0",
-31169 => x"C0C0BFB0F9F98290",
-31168 => x"C0C0BFB0F9F98280",
-31167 => x"C0C0BFB0F9F982F8",
-31166 => x"C0C0BFB0F9F98282",
-31165 => x"C0C0BFB0F9F98292",
-31164 => x"C0C0BFB0F9F98299",
-31163 => x"C0C0BFB0F9F982B0",
-31162 => x"C0C0BFB0F9F982A4",
-31161 => x"C0C0BFB0F9F982F9",
-31160 => x"C0C0BFB0F9F982C0",
-31159 => x"C0C0BFB0F9F99290",
-31158 => x"C0C0BFB0F9F99280",
-31157 => x"C0C0BFB0F9F992F8",
-31156 => x"C0C0BFB0F9F99282",
-31155 => x"C0C0BFB0F9F99292",
-31154 => x"C0C0BFB0F9F99299",
-31153 => x"C0C0BFB0F9F992B0",
-31152 => x"C0C0BFB0F9F992A4",
-31151 => x"C0C0BFB0F9F992F9",
-31150 => x"C0C0BFB0F9F992C0",
-31149 => x"C0C0BFB0F9F99990",
-31148 => x"C0C0BFB0F9F99980",
-31147 => x"C0C0BFB0F9F999F8",
-31146 => x"C0C0BFB0F9F99982",
-31145 => x"C0C0BFB0F9F99992",
-31144 => x"C0C0BFB0F9F99999",
-31143 => x"C0C0BFB0F9F999B0",
-31142 => x"C0C0BFB0F9F999A4",
-31141 => x"C0C0BFB0F9F999F9",
-31140 => x"C0C0BFB0F9F999C0",
-31139 => x"C0C0BFB0F9F9B090",
-31138 => x"C0C0BFB0F9F9B080",
-31137 => x"C0C0BFB0F9F9B0F8",
-31136 => x"C0C0BFB0F9F9B082",
-31135 => x"C0C0BFB0F9F9B092",
-31134 => x"C0C0BFB0F9F9B099",
-31133 => x"C0C0BFB0F9F9B0B0",
-31132 => x"C0C0BFB0F9F9B0A4",
-31131 => x"C0C0BFB0F9F9B0F9",
-31130 => x"C0C0BFB0F9F9B0C0",
-31129 => x"C0C0BFB0F9F9A490",
-31128 => x"C0C0BFB0F9F9A480",
-31127 => x"C0C0BFB0F9F9A4F8",
-31126 => x"C0C0BFB0F9F9A482",
-31125 => x"C0C0BFB0F9F9A492",
-31124 => x"C0C0BFB0F9F9A499",
-31123 => x"C0C0BFB0F9F9A4B0",
-31122 => x"C0C0BFB0F9F9A4A4",
-31121 => x"C0C0BFB0F9F9A4F9",
-31120 => x"C0C0BFB0F9F9A4C0",
-31119 => x"C0C0BFB0F9F9F990",
-31118 => x"C0C0BFB0F9F9F980",
-31117 => x"C0C0BFB0F9F9F9F8",
-31116 => x"C0C0BFB0F9F9F982",
-31115 => x"C0C0BFB0F9F9F992",
-31114 => x"C0C0BFB0F9F9F999",
-31113 => x"C0C0BFB0F9F9F9B0",
-31112 => x"C0C0BFB0F9F9F9A4",
-31111 => x"C0C0BFB0F9F9F9F9",
-31110 => x"C0C0BFB0F9F9F9C0",
-31109 => x"C0C0BFB0F9F9C090",
-31108 => x"C0C0BFB0F9F9C080",
-31107 => x"C0C0BFB0F9F9C0F8",
-31106 => x"C0C0BFB0F9F9C082",
-31105 => x"C0C0BFB0F9F9C092",
-31104 => x"C0C0BFB0F9F9C099",
-31103 => x"C0C0BFB0F9F9C0B0",
-31102 => x"C0C0BFB0F9F9C0A4",
-31101 => x"C0C0BFB0F9F9C0F9",
-31100 => x"C0C0BFB0F9F9C0C0",
-31099 => x"C0C0BFB0F9C09090",
-31098 => x"C0C0BFB0F9C09080",
-31097 => x"C0C0BFB0F9C090F8",
-31096 => x"C0C0BFB0F9C09082",
-31095 => x"C0C0BFB0F9C09092",
-31094 => x"C0C0BFB0F9C09099",
-31093 => x"C0C0BFB0F9C090B0",
-31092 => x"C0C0BFB0F9C090A4",
-31091 => x"C0C0BFB0F9C090F9",
-31090 => x"C0C0BFB0F9C090C0",
-31089 => x"C0C0BFB0F9C08090",
-31088 => x"C0C0BFB0F9C08080",
-31087 => x"C0C0BFB0F9C080F8",
-31086 => x"C0C0BFB0F9C08082",
-31085 => x"C0C0BFB0F9C08092",
-31084 => x"C0C0BFB0F9C08099",
-31083 => x"C0C0BFB0F9C080B0",
-31082 => x"C0C0BFB0F9C080A4",
-31081 => x"C0C0BFB0F9C080F9",
-31080 => x"C0C0BFB0F9C080C0",
-31079 => x"C0C0BFB0F9C0F890",
-31078 => x"C0C0BFB0F9C0F880",
-31077 => x"C0C0BFB0F9C0F8F8",
-31076 => x"C0C0BFB0F9C0F882",
-31075 => x"C0C0BFB0F9C0F892",
-31074 => x"C0C0BFB0F9C0F899",
-31073 => x"C0C0BFB0F9C0F8B0",
-31072 => x"C0C0BFB0F9C0F8A4",
-31071 => x"C0C0BFB0F9C0F8F9",
-31070 => x"C0C0BFB0F9C0F8C0",
-31069 => x"C0C0BFB0F9C08290",
-31068 => x"C0C0BFB0F9C08280",
-31067 => x"C0C0BFB0F9C082F8",
-31066 => x"C0C0BFB0F9C08282",
-31065 => x"C0C0BFB0F9C08292",
-31064 => x"C0C0BFB0F9C08299",
-31063 => x"C0C0BFB0F9C082B0",
-31062 => x"C0C0BFB0F9C082A4",
-31061 => x"C0C0BFB0F9C082F9",
-31060 => x"C0C0BFB0F9C082C0",
-31059 => x"C0C0BFB0F9C09290",
-31058 => x"C0C0BFB0F9C09280",
-31057 => x"C0C0BFB0F9C092F8",
-31056 => x"C0C0BFB0F9C09282",
-31055 => x"C0C0BFB0F9C09292",
-31054 => x"C0C0BFB0F9C09299",
-31053 => x"C0C0BFB0F9C092B0",
-31052 => x"C0C0BFB0F9C092A4",
-31051 => x"C0C0BFB0F9C092F9",
-31050 => x"C0C0BFB0F9C092C0",
-31049 => x"C0C0BFB0F9C09990",
-31048 => x"C0C0BFB0F9C09980",
-31047 => x"C0C0BFB0F9C099F8",
-31046 => x"C0C0BFB0F9C09982",
-31045 => x"C0C0BFB0F9C09992",
-31044 => x"C0C0BFB0F9C09999",
-31043 => x"C0C0BFB0F9C099B0",
-31042 => x"C0C0BFB0F9C099A4",
-31041 => x"C0C0BFB0F9C099F9",
-31040 => x"C0C0BFB0F9C099C0",
-31039 => x"C0C0BFB0F9C0B090",
-31038 => x"C0C0BFB0F9C0B080",
-31037 => x"C0C0BFB0F9C0B0F8",
-31036 => x"C0C0BFB0F9C0B082",
-31035 => x"C0C0BFB0F9C0B092",
-31034 => x"C0C0BFB0F9C0B099",
-31033 => x"C0C0BFB0F9C0B0B0",
-31032 => x"C0C0BFB0F9C0B0A4",
-31031 => x"C0C0BFB0F9C0B0F9",
-31030 => x"C0C0BFB0F9C0B0C0",
-31029 => x"C0C0BFB0F9C0A490",
-31028 => x"C0C0BFB0F9C0A480",
-31027 => x"C0C0BFB0F9C0A4F8",
-31026 => x"C0C0BFB0F9C0A482",
-31025 => x"C0C0BFB0F9C0A492",
-31024 => x"C0C0BFB0F9C0A499",
-31023 => x"C0C0BFB0F9C0A4B0",
-31022 => x"C0C0BFB0F9C0A4A4",
-31021 => x"C0C0BFB0F9C0A4F9",
-31020 => x"C0C0BFB0F9C0A4C0",
-31019 => x"C0C0BFB0F9C0F990",
-31018 => x"C0C0BFB0F9C0F980",
-31017 => x"C0C0BFB0F9C0F9F8",
-31016 => x"C0C0BFB0F9C0F982",
-31015 => x"C0C0BFB0F9C0F992",
-31014 => x"C0C0BFB0F9C0F999",
-31013 => x"C0C0BFB0F9C0F9B0",
-31012 => x"C0C0BFB0F9C0F9A4",
-31011 => x"C0C0BFB0F9C0F9F9",
-31010 => x"C0C0BFB0F9C0F9C0",
-31009 => x"C0C0BFB0F9C0C090",
-31008 => x"C0C0BFB0F9C0C080",
-31007 => x"C0C0BFB0F9C0C0F8",
-31006 => x"C0C0BFB0F9C0C082",
-31005 => x"C0C0BFB0F9C0C092",
-31004 => x"C0C0BFB0F9C0C099",
-31003 => x"C0C0BFB0F9C0C0B0",
-31002 => x"C0C0BFB0F9C0C0A4",
-31001 => x"C0C0BFB0F9C0C0F9",
-31000 => x"C0C0BFB0F9C0C0C0",
-30999 => x"C0C0BFB0C0909090",
-30998 => x"C0C0BFB0C0909080",
-30997 => x"C0C0BFB0C09090F8",
-30996 => x"C0C0BFB0C0909082",
-30995 => x"C0C0BFB0C0909092",
-30994 => x"C0C0BFB0C0909099",
-30993 => x"C0C0BFB0C09090B0",
-30992 => x"C0C0BFB0C09090A4",
-30991 => x"C0C0BFB0C09090F9",
-30990 => x"C0C0BFB0C09090C0",
-30989 => x"C0C0BFB0C0908090",
-30988 => x"C0C0BFB0C0908080",
-30987 => x"C0C0BFB0C09080F8",
-30986 => x"C0C0BFB0C0908082",
-30985 => x"C0C0BFB0C0908092",
-30984 => x"C0C0BFB0C0908099",
-30983 => x"C0C0BFB0C09080B0",
-30982 => x"C0C0BFB0C09080A4",
-30981 => x"C0C0BFB0C09080F9",
-30980 => x"C0C0BFB0C09080C0",
-30979 => x"C0C0BFB0C090F890",
-30978 => x"C0C0BFB0C090F880",
-30977 => x"C0C0BFB0C090F8F8",
-30976 => x"C0C0BFB0C090F882",
-30975 => x"C0C0BFB0C090F892",
-30974 => x"C0C0BFB0C090F899",
-30973 => x"C0C0BFB0C090F8B0",
-30972 => x"C0C0BFB0C090F8A4",
-30971 => x"C0C0BFB0C090F8F9",
-30970 => x"C0C0BFB0C090F8C0",
-30969 => x"C0C0BFB0C0908290",
-30968 => x"C0C0BFB0C0908280",
-30967 => x"C0C0BFB0C09082F8",
-30966 => x"C0C0BFB0C0908282",
-30965 => x"C0C0BFB0C0908292",
-30964 => x"C0C0BFB0C0908299",
-30963 => x"C0C0BFB0C09082B0",
-30962 => x"C0C0BFB0C09082A4",
-30961 => x"C0C0BFB0C09082F9",
-30960 => x"C0C0BFB0C09082C0",
-30959 => x"C0C0BFB0C0909290",
-30958 => x"C0C0BFB0C0909280",
-30957 => x"C0C0BFB0C09092F8",
-30956 => x"C0C0BFB0C0909282",
-30955 => x"C0C0BFB0C0909292",
-30954 => x"C0C0BFB0C0909299",
-30953 => x"C0C0BFB0C09092B0",
-30952 => x"C0C0BFB0C09092A4",
-30951 => x"C0C0BFB0C09092F9",
-30950 => x"C0C0BFB0C09092C0",
-30949 => x"C0C0BFB0C0909990",
-30948 => x"C0C0BFB0C0909980",
-30947 => x"C0C0BFB0C09099F8",
-30946 => x"C0C0BFB0C0909982",
-30945 => x"C0C0BFB0C0909992",
-30944 => x"C0C0BFB0C0909999",
-30943 => x"C0C0BFB0C09099B0",
-30942 => x"C0C0BFB0C09099A4",
-30941 => x"C0C0BFB0C09099F9",
-30940 => x"C0C0BFB0C09099C0",
-30939 => x"C0C0BFB0C090B090",
-30938 => x"C0C0BFB0C090B080",
-30937 => x"C0C0BFB0C090B0F8",
-30936 => x"C0C0BFB0C090B082",
-30935 => x"C0C0BFB0C090B092",
-30934 => x"C0C0BFB0C090B099",
-30933 => x"C0C0BFB0C090B0B0",
-30932 => x"C0C0BFB0C090B0A4",
-30931 => x"C0C0BFB0C090B0F9",
-30930 => x"C0C0BFB0C090B0C0",
-30929 => x"C0C0BFB0C090A490",
-30928 => x"C0C0BFB0C090A480",
-30927 => x"C0C0BFB0C090A4F8",
-30926 => x"C0C0BFB0C090A482",
-30925 => x"C0C0BFB0C090A492",
-30924 => x"C0C0BFB0C090A499",
-30923 => x"C0C0BFB0C090A4B0",
-30922 => x"C0C0BFB0C090A4A4",
-30921 => x"C0C0BFB0C090A4F9",
-30920 => x"C0C0BFB0C090A4C0",
-30919 => x"C0C0BFB0C090F990",
-30918 => x"C0C0BFB0C090F980",
-30917 => x"C0C0BFB0C090F9F8",
-30916 => x"C0C0BFB0C090F982",
-30915 => x"C0C0BFB0C090F992",
-30914 => x"C0C0BFB0C090F999",
-30913 => x"C0C0BFB0C090F9B0",
-30912 => x"C0C0BFB0C090F9A4",
-30911 => x"C0C0BFB0C090F9F9",
-30910 => x"C0C0BFB0C090F9C0",
-30909 => x"C0C0BFB0C090C090",
-30908 => x"C0C0BFB0C090C080",
-30907 => x"C0C0BFB0C090C0F8",
-30906 => x"C0C0BFB0C090C082",
-30905 => x"C0C0BFB0C090C092",
-30904 => x"C0C0BFB0C090C099",
-30903 => x"C0C0BFB0C090C0B0",
-30902 => x"C0C0BFB0C090C0A4",
-30901 => x"C0C0BFB0C090C0F9",
-30900 => x"C0C0BFB0C090C0C0",
-30899 => x"C0C0BFB0C0809090",
-30898 => x"C0C0BFB0C0809080",
-30897 => x"C0C0BFB0C08090F8",
-30896 => x"C0C0BFB0C0809082",
-30895 => x"C0C0BFB0C0809092",
-30894 => x"C0C0BFB0C0809099",
-30893 => x"C0C0BFB0C08090B0",
-30892 => x"C0C0BFB0C08090A4",
-30891 => x"C0C0BFB0C08090F9",
-30890 => x"C0C0BFB0C08090C0",
-30889 => x"C0C0BFB0C0808090",
-30888 => x"C0C0BFB0C0808080",
-30887 => x"C0C0BFB0C08080F8",
-30886 => x"C0C0BFB0C0808082",
-30885 => x"C0C0BFB0C0808092",
-30884 => x"C0C0BFB0C0808099",
-30883 => x"C0C0BFB0C08080B0",
-30882 => x"C0C0BFB0C08080A4",
-30881 => x"C0C0BFB0C08080F9",
-30880 => x"C0C0BFB0C08080C0",
-30879 => x"C0C0BFB0C080F890",
-30878 => x"C0C0BFB0C080F880",
-30877 => x"C0C0BFB0C080F8F8",
-30876 => x"C0C0BFB0C080F882",
-30875 => x"C0C0BFB0C080F892",
-30874 => x"C0C0BFB0C080F899",
-30873 => x"C0C0BFB0C080F8B0",
-30872 => x"C0C0BFB0C080F8A4",
-30871 => x"C0C0BFB0C080F8F9",
-30870 => x"C0C0BFB0C080F8C0",
-30869 => x"C0C0BFB0C0808290",
-30868 => x"C0C0BFB0C0808280",
-30867 => x"C0C0BFB0C08082F8",
-30866 => x"C0C0BFB0C0808282",
-30865 => x"C0C0BFB0C0808292",
-30864 => x"C0C0BFB0C0808299",
-30863 => x"C0C0BFB0C08082B0",
-30862 => x"C0C0BFB0C08082A4",
-30861 => x"C0C0BFB0C08082F9",
-30860 => x"C0C0BFB0C08082C0",
-30859 => x"C0C0BFB0C0809290",
-30858 => x"C0C0BFB0C0809280",
-30857 => x"C0C0BFB0C08092F8",
-30856 => x"C0C0BFB0C0809282",
-30855 => x"C0C0BFB0C0809292",
-30854 => x"C0C0BFB0C0809299",
-30853 => x"C0C0BFB0C08092B0",
-30852 => x"C0C0BFB0C08092A4",
-30851 => x"C0C0BFB0C08092F9",
-30850 => x"C0C0BFB0C08092C0",
-30849 => x"C0C0BFB0C0809990",
-30848 => x"C0C0BFB0C0809980",
-30847 => x"C0C0BFB0C08099F8",
-30846 => x"C0C0BFB0C0809982",
-30845 => x"C0C0BFB0C0809992",
-30844 => x"C0C0BFB0C0809999",
-30843 => x"C0C0BFB0C08099B0",
-30842 => x"C0C0BFB0C08099A4",
-30841 => x"C0C0BFB0C08099F9",
-30840 => x"C0C0BFB0C08099C0",
-30839 => x"C0C0BFB0C080B090",
-30838 => x"C0C0BFB0C080B080",
-30837 => x"C0C0BFB0C080B0F8",
-30836 => x"C0C0BFB0C080B082",
-30835 => x"C0C0BFB0C080B092",
-30834 => x"C0C0BFB0C080B099",
-30833 => x"C0C0BFB0C080B0B0",
-30832 => x"C0C0BFB0C080B0A4",
-30831 => x"C0C0BFB0C080B0F9",
-30830 => x"C0C0BFB0C080B0C0",
-30829 => x"C0C0BFB0C080A490",
-30828 => x"C0C0BFB0C080A480",
-30827 => x"C0C0BFB0C080A4F8",
-30826 => x"C0C0BFB0C080A482",
-30825 => x"C0C0BFB0C080A492",
-30824 => x"C0C0BFB0C080A499",
-30823 => x"C0C0BFB0C080A4B0",
-30822 => x"C0C0BFB0C080A4A4",
-30821 => x"C0C0BFB0C080A4F9",
-30820 => x"C0C0BFB0C080A4C0",
-30819 => x"C0C0BFB0C080F990",
-30818 => x"C0C0BFB0C080F980",
-30817 => x"C0C0BFB0C080F9F8",
-30816 => x"C0C0BFB0C080F982",
-30815 => x"C0C0BFB0C080F992",
-30814 => x"C0C0BFB0C080F999",
-30813 => x"C0C0BFB0C080F9B0",
-30812 => x"C0C0BFB0C080F9A4",
-30811 => x"C0C0BFB0C080F9F9",
-30810 => x"C0C0BFB0C080F9C0",
-30809 => x"C0C0BFB0C080C090",
-30808 => x"C0C0BFB0C080C080",
-30807 => x"C0C0BFB0C080C0F8",
-30806 => x"C0C0BFB0C080C082",
-30805 => x"C0C0BFB0C080C092",
-30804 => x"C0C0BFB0C080C099",
-30803 => x"C0C0BFB0C080C0B0",
-30802 => x"C0C0BFB0C080C0A4",
-30801 => x"C0C0BFB0C080C0F9",
-30800 => x"C0C0BFB0C080C0C0",
-30799 => x"C0C0BFB0C0F89090",
-30798 => x"C0C0BFB0C0F89080",
-30797 => x"C0C0BFB0C0F890F8",
-30796 => x"C0C0BFB0C0F89082",
-30795 => x"C0C0BFB0C0F89092",
-30794 => x"C0C0BFB0C0F89099",
-30793 => x"C0C0BFB0C0F890B0",
-30792 => x"C0C0BFB0C0F890A4",
-30791 => x"C0C0BFB0C0F890F9",
-30790 => x"C0C0BFB0C0F890C0",
-30789 => x"C0C0BFB0C0F88090",
-30788 => x"C0C0BFB0C0F88080",
-30787 => x"C0C0BFB0C0F880F8",
-30786 => x"C0C0BFB0C0F88082",
-30785 => x"C0C0BFB0C0F88092",
-30784 => x"C0C0BFB0C0F88099",
-30783 => x"C0C0BFB0C0F880B0",
-30782 => x"C0C0BFB0C0F880A4",
-30781 => x"C0C0BFB0C0F880F9",
-30780 => x"C0C0BFB0C0F880C0",
-30779 => x"C0C0BFB0C0F8F890",
-30778 => x"C0C0BFB0C0F8F880",
-30777 => x"C0C0BFB0C0F8F8F8",
-30776 => x"C0C0BFB0C0F8F882",
-30775 => x"C0C0BFB0C0F8F892",
-30774 => x"C0C0BFB0C0F8F899",
-30773 => x"C0C0BFB0C0F8F8B0",
-30772 => x"C0C0BFB0C0F8F8A4",
-30771 => x"C0C0BFB0C0F8F8F9",
-30770 => x"C0C0BFB0C0F8F8C0",
-30769 => x"C0C0BFB0C0F88290",
-30768 => x"C0C0BFB0C0F88280",
-30767 => x"C0C0BFB0C0F882F8",
-30766 => x"C0C0BFB0C0F88282",
-30765 => x"C0C0BFB0C0F88292",
-30764 => x"C0C0BFB0C0F88299",
-30763 => x"C0C0BFB0C0F882B0",
-30762 => x"C0C0BFB0C0F882A4",
-30761 => x"C0C0BFB0C0F882F9",
-30760 => x"C0C0BFB0C0F882C0",
-30759 => x"C0C0BFB0C0F89290",
-30758 => x"C0C0BFB0C0F89280",
-30757 => x"C0C0BFB0C0F892F8",
-30756 => x"C0C0BFB0C0F89282",
-30755 => x"C0C0BFB0C0F89292",
-30754 => x"C0C0BFB0C0F89299",
-30753 => x"C0C0BFB0C0F892B0",
-30752 => x"C0C0BFB0C0F892A4",
-30751 => x"C0C0BFB0C0F892F9",
-30750 => x"C0C0BFB0C0F892C0",
-30749 => x"C0C0BFB0C0F89990",
-30748 => x"C0C0BFB0C0F89980",
-30747 => x"C0C0BFB0C0F899F8",
-30746 => x"C0C0BFB0C0F89982",
-30745 => x"C0C0BFB0C0F89992",
-30744 => x"C0C0BFB0C0F89999",
-30743 => x"C0C0BFB0C0F899B0",
-30742 => x"C0C0BFB0C0F899A4",
-30741 => x"C0C0BFB0C0F899F9",
-30740 => x"C0C0BFB0C0F899C0",
-30739 => x"C0C0BFB0C0F8B090",
-30738 => x"C0C0BFB0C0F8B080",
-30737 => x"C0C0BFB0C0F8B0F8",
-30736 => x"C0C0BFB0C0F8B082",
-30735 => x"C0C0BFB0C0F8B092",
-30734 => x"C0C0BFB0C0F8B099",
-30733 => x"C0C0BFB0C0F8B0B0",
-30732 => x"C0C0BFB0C0F8B0A4",
-30731 => x"C0C0BFB0C0F8B0F9",
-30730 => x"C0C0BFB0C0F8B0C0",
-30729 => x"C0C0BFB0C0F8A490",
-30728 => x"C0C0BFB0C0F8A480",
-30727 => x"C0C0BFB0C0F8A4F8",
-30726 => x"C0C0BFB0C0F8A482",
-30725 => x"C0C0BFB0C0F8A492",
-30724 => x"C0C0BFB0C0F8A499",
-30723 => x"C0C0BFB0C0F8A4B0",
-30722 => x"C0C0BFB0C0F8A4A4",
-30721 => x"C0C0BFB0C0F8A4F9",
-30720 => x"C0C0BFB0C0F8A4C0",
-30719 => x"C0C0BFB0C0F8F990",
-30718 => x"C0C0BFB0C0F8F980",
-30717 => x"C0C0BFB0C0F8F9F8",
-30716 => x"C0C0BFB0C0F8F982",
-30715 => x"C0C0BFB0C0F8F992",
-30714 => x"C0C0BFB0C0F8F999",
-30713 => x"C0C0BFB0C0F8F9B0",
-30712 => x"C0C0BFB0C0F8F9A4",
-30711 => x"C0C0BFB0C0F8F9F9",
-30710 => x"C0C0BFB0C0F8F9C0",
-30709 => x"C0C0BFB0C0F8C090",
-30708 => x"C0C0BFB0C0F8C080",
-30707 => x"C0C0BFB0C0F8C0F8",
-30706 => x"C0C0BFB0C0F8C082",
-30705 => x"C0C0BFB0C0F8C092",
-30704 => x"C0C0BFB0C0F8C099",
-30703 => x"C0C0BFB0C0F8C0B0",
-30702 => x"C0C0BFB0C0F8C0A4",
-30701 => x"C0C0BFB0C0F8C0F9",
-30700 => x"C0C0BFB0C0F8C0C0",
-30699 => x"C0C0BFB0C0829090",
-30698 => x"C0C0BFB0C0829080",
-30697 => x"C0C0BFB0C08290F8",
-30696 => x"C0C0BFB0C0829082",
-30695 => x"C0C0BFB0C0829092",
-30694 => x"C0C0BFB0C0829099",
-30693 => x"C0C0BFB0C08290B0",
-30692 => x"C0C0BFB0C08290A4",
-30691 => x"C0C0BFB0C08290F9",
-30690 => x"C0C0BFB0C08290C0",
-30689 => x"C0C0BFB0C0828090",
-30688 => x"C0C0BFB0C0828080",
-30687 => x"C0C0BFB0C08280F8",
-30686 => x"C0C0BFB0C0828082",
-30685 => x"C0C0BFB0C0828092",
-30684 => x"C0C0BFB0C0828099",
-30683 => x"C0C0BFB0C08280B0",
-30682 => x"C0C0BFB0C08280A4",
-30681 => x"C0C0BFB0C08280F9",
-30680 => x"C0C0BFB0C08280C0",
-30679 => x"C0C0BFB0C082F890",
-30678 => x"C0C0BFB0C082F880",
-30677 => x"C0C0BFB0C082F8F8",
-30676 => x"C0C0BFB0C082F882",
-30675 => x"C0C0BFB0C082F892",
-30674 => x"C0C0BFB0C082F899",
-30673 => x"C0C0BFB0C082F8B0",
-30672 => x"C0C0BFB0C082F8A4",
-30671 => x"C0C0BFB0C082F8F9",
-30670 => x"C0C0BFB0C082F8C0",
-30669 => x"C0C0BFB0C0828290",
-30668 => x"C0C0BFB0C0828280",
-30667 => x"C0C0BFB0C08282F8",
-30666 => x"C0C0BFB0C0828282",
-30665 => x"C0C0BFB0C0828292",
-30664 => x"C0C0BFB0C0828299",
-30663 => x"C0C0BFB0C08282B0",
-30662 => x"C0C0BFB0C08282A4",
-30661 => x"C0C0BFB0C08282F9",
-30660 => x"C0C0BFB0C08282C0",
-30659 => x"C0C0BFB0C0829290",
-30658 => x"C0C0BFB0C0829280",
-30657 => x"C0C0BFB0C08292F8",
-30656 => x"C0C0BFB0C0829282",
-30655 => x"C0C0BFB0C0829292",
-30654 => x"C0C0BFB0C0829299",
-30653 => x"C0C0BFB0C08292B0",
-30652 => x"C0C0BFB0C08292A4",
-30651 => x"C0C0BFB0C08292F9",
-30650 => x"C0C0BFB0C08292C0",
-30649 => x"C0C0BFB0C0829990",
-30648 => x"C0C0BFB0C0829980",
-30647 => x"C0C0BFB0C08299F8",
-30646 => x"C0C0BFB0C0829982",
-30645 => x"C0C0BFB0C0829992",
-30644 => x"C0C0BFB0C0829999",
-30643 => x"C0C0BFB0C08299B0",
-30642 => x"C0C0BFB0C08299A4",
-30641 => x"C0C0BFB0C08299F9",
-30640 => x"C0C0BFB0C08299C0",
-30639 => x"C0C0BFB0C082B090",
-30638 => x"C0C0BFB0C082B080",
-30637 => x"C0C0BFB0C082B0F8",
-30636 => x"C0C0BFB0C082B082",
-30635 => x"C0C0BFB0C082B092",
-30634 => x"C0C0BFB0C082B099",
-30633 => x"C0C0BFB0C082B0B0",
-30632 => x"C0C0BFB0C082B0A4",
-30631 => x"C0C0BFB0C082B0F9",
-30630 => x"C0C0BFB0C082B0C0",
-30629 => x"C0C0BFB0C082A490",
-30628 => x"C0C0BFB0C082A480",
-30627 => x"C0C0BFB0C082A4F8",
-30626 => x"C0C0BFB0C082A482",
-30625 => x"C0C0BFB0C082A492",
-30624 => x"C0C0BFB0C082A499",
-30623 => x"C0C0BFB0C082A4B0",
-30622 => x"C0C0BFB0C082A4A4",
-30621 => x"C0C0BFB0C082A4F9",
-30620 => x"C0C0BFB0C082A4C0",
-30619 => x"C0C0BFB0C082F990",
-30618 => x"C0C0BFB0C082F980",
-30617 => x"C0C0BFB0C082F9F8",
-30616 => x"C0C0BFB0C082F982",
-30615 => x"C0C0BFB0C082F992",
-30614 => x"C0C0BFB0C082F999",
-30613 => x"C0C0BFB0C082F9B0",
-30612 => x"C0C0BFB0C082F9A4",
-30611 => x"C0C0BFB0C082F9F9",
-30610 => x"C0C0BFB0C082F9C0",
-30609 => x"C0C0BFB0C082C090",
-30608 => x"C0C0BFB0C082C080",
-30607 => x"C0C0BFB0C082C0F8",
-30606 => x"C0C0BFB0C082C082",
-30605 => x"C0C0BFB0C082C092",
-30604 => x"C0C0BFB0C082C099",
-30603 => x"C0C0BFB0C082C0B0",
-30602 => x"C0C0BFB0C082C0A4",
-30601 => x"C0C0BFB0C082C0F9",
-30600 => x"C0C0BFB0C082C0C0",
-30599 => x"C0C0BFB0C0929090",
-30598 => x"C0C0BFB0C0929080",
-30597 => x"C0C0BFB0C09290F8",
-30596 => x"C0C0BFB0C0929082",
-30595 => x"C0C0BFB0C0929092",
-30594 => x"C0C0BFB0C0929099",
-30593 => x"C0C0BFB0C09290B0",
-30592 => x"C0C0BFB0C09290A4",
-30591 => x"C0C0BFB0C09290F9",
-30590 => x"C0C0BFB0C09290C0",
-30589 => x"C0C0BFB0C0928090",
-30588 => x"C0C0BFB0C0928080",
-30587 => x"C0C0BFB0C09280F8",
-30586 => x"C0C0BFB0C0928082",
-30585 => x"C0C0BFB0C0928092",
-30584 => x"C0C0BFB0C0928099",
-30583 => x"C0C0BFB0C09280B0",
-30582 => x"C0C0BFB0C09280A4",
-30581 => x"C0C0BFB0C09280F9",
-30580 => x"C0C0BFB0C09280C0",
-30579 => x"C0C0BFB0C092F890",
-30578 => x"C0C0BFB0C092F880",
-30577 => x"C0C0BFB0C092F8F8",
-30576 => x"C0C0BFB0C092F882",
-30575 => x"C0C0BFB0C092F892",
-30574 => x"C0C0BFB0C092F899",
-30573 => x"C0C0BFB0C092F8B0",
-30572 => x"C0C0BFB0C092F8A4",
-30571 => x"C0C0BFB0C092F8F9",
-30570 => x"C0C0BFB0C092F8C0",
-30569 => x"C0C0BFB0C0928290",
-30568 => x"C0C0BFB0C0928280",
-30567 => x"C0C0BFB0C09282F8",
-30566 => x"C0C0BFB0C0928282",
-30565 => x"C0C0BFB0C0928292",
-30564 => x"C0C0BFB0C0928299",
-30563 => x"C0C0BFB0C09282B0",
-30562 => x"C0C0BFB0C09282A4",
-30561 => x"C0C0BFB0C09282F9",
-30560 => x"C0C0BFB0C09282C0",
-30559 => x"C0C0BFB0C0929290",
-30558 => x"C0C0BFB0C0929280",
-30557 => x"C0C0BFB0C09292F8",
-30556 => x"C0C0BFB0C0929282",
-30555 => x"C0C0BFB0C0929292",
-30554 => x"C0C0BFB0C0929299",
-30553 => x"C0C0BFB0C09292B0",
-30552 => x"C0C0BFB0C09292A4",
-30551 => x"C0C0BFB0C09292F9",
-30550 => x"C0C0BFB0C09292C0",
-30549 => x"C0C0BFB0C0929990",
-30548 => x"C0C0BFB0C0929980",
-30547 => x"C0C0BFB0C09299F8",
-30546 => x"C0C0BFB0C0929982",
-30545 => x"C0C0BFB0C0929992",
-30544 => x"C0C0BFB0C0929999",
-30543 => x"C0C0BFB0C09299B0",
-30542 => x"C0C0BFB0C09299A4",
-30541 => x"C0C0BFB0C09299F9",
-30540 => x"C0C0BFB0C09299C0",
-30539 => x"C0C0BFB0C092B090",
-30538 => x"C0C0BFB0C092B080",
-30537 => x"C0C0BFB0C092B0F8",
-30536 => x"C0C0BFB0C092B082",
-30535 => x"C0C0BFB0C092B092",
-30534 => x"C0C0BFB0C092B099",
-30533 => x"C0C0BFB0C092B0B0",
-30532 => x"C0C0BFB0C092B0A4",
-30531 => x"C0C0BFB0C092B0F9",
-30530 => x"C0C0BFB0C092B0C0",
-30529 => x"C0C0BFB0C092A490",
-30528 => x"C0C0BFB0C092A480",
-30527 => x"C0C0BFB0C092A4F8",
-30526 => x"C0C0BFB0C092A482",
-30525 => x"C0C0BFB0C092A492",
-30524 => x"C0C0BFB0C092A499",
-30523 => x"C0C0BFB0C092A4B0",
-30522 => x"C0C0BFB0C092A4A4",
-30521 => x"C0C0BFB0C092A4F9",
-30520 => x"C0C0BFB0C092A4C0",
-30519 => x"C0C0BFB0C092F990",
-30518 => x"C0C0BFB0C092F980",
-30517 => x"C0C0BFB0C092F9F8",
-30516 => x"C0C0BFB0C092F982",
-30515 => x"C0C0BFB0C092F992",
-30514 => x"C0C0BFB0C092F999",
-30513 => x"C0C0BFB0C092F9B0",
-30512 => x"C0C0BFB0C092F9A4",
-30511 => x"C0C0BFB0C092F9F9",
-30510 => x"C0C0BFB0C092F9C0",
-30509 => x"C0C0BFB0C092C090",
-30508 => x"C0C0BFB0C092C080",
-30507 => x"C0C0BFB0C092C0F8",
-30506 => x"C0C0BFB0C092C082",
-30505 => x"C0C0BFB0C092C092",
-30504 => x"C0C0BFB0C092C099",
-30503 => x"C0C0BFB0C092C0B0",
-30502 => x"C0C0BFB0C092C0A4",
-30501 => x"C0C0BFB0C092C0F9",
-30500 => x"C0C0BFB0C092C0C0",
-30499 => x"C0C0BFB0C0999090",
-30498 => x"C0C0BFB0C0999080",
-30497 => x"C0C0BFB0C09990F8",
-30496 => x"C0C0BFB0C0999082",
-30495 => x"C0C0BFB0C0999092",
-30494 => x"C0C0BFB0C0999099",
-30493 => x"C0C0BFB0C09990B0",
-30492 => x"C0C0BFB0C09990A4",
-30491 => x"C0C0BFB0C09990F9",
-30490 => x"C0C0BFB0C09990C0",
-30489 => x"C0C0BFB0C0998090",
-30488 => x"C0C0BFB0C0998080",
-30487 => x"C0C0BFB0C09980F8",
-30486 => x"C0C0BFB0C0998082",
-30485 => x"C0C0BFB0C0998092",
-30484 => x"C0C0BFB0C0998099",
-30483 => x"C0C0BFB0C09980B0",
-30482 => x"C0C0BFB0C09980A4",
-30481 => x"C0C0BFB0C09980F9",
-30480 => x"C0C0BFB0C09980C0",
-30479 => x"C0C0BFB0C099F890",
-30478 => x"C0C0BFB0C099F880",
-30477 => x"C0C0BFB0C099F8F8",
-30476 => x"C0C0BFB0C099F882",
-30475 => x"C0C0BFB0C099F892",
-30474 => x"C0C0BFB0C099F899",
-30473 => x"C0C0BFB0C099F8B0",
-30472 => x"C0C0BFB0C099F8A4",
-30471 => x"C0C0BFB0C099F8F9",
-30470 => x"C0C0BFB0C099F8C0",
-30469 => x"C0C0BFB0C0998290",
-30468 => x"C0C0BFB0C0998280",
-30467 => x"C0C0BFB0C09982F8",
-30466 => x"C0C0BFB0C0998282",
-30465 => x"C0C0BFB0C0998292",
-30464 => x"C0C0BFB0C0998299",
-30463 => x"C0C0BFB0C09982B0",
-30462 => x"C0C0BFB0C09982A4",
-30461 => x"C0C0BFB0C09982F9",
-30460 => x"C0C0BFB0C09982C0",
-30459 => x"C0C0BFB0C0999290",
-30458 => x"C0C0BFB0C0999280",
-30457 => x"C0C0BFB0C09992F8",
-30456 => x"C0C0BFB0C0999282",
-30455 => x"C0C0BFB0C0999292",
-30454 => x"C0C0BFB0C0999299",
-30453 => x"C0C0BFB0C09992B0",
-30452 => x"C0C0BFB0C09992A4",
-30451 => x"C0C0BFB0C09992F9",
-30450 => x"C0C0BFB0C09992C0",
-30449 => x"C0C0BFB0C0999990",
-30448 => x"C0C0BFB0C0999980",
-30447 => x"C0C0BFB0C09999F8",
-30446 => x"C0C0BFB0C0999982",
-30445 => x"C0C0BFB0C0999992",
-30444 => x"C0C0BFB0C0999999",
-30443 => x"C0C0BFB0C09999B0",
-30442 => x"C0C0BFB0C09999A4",
-30441 => x"C0C0BFB0C09999F9",
-30440 => x"C0C0BFB0C09999C0",
-30439 => x"C0C0BFB0C099B090",
-30438 => x"C0C0BFB0C099B080",
-30437 => x"C0C0BFB0C099B0F8",
-30436 => x"C0C0BFB0C099B082",
-30435 => x"C0C0BFB0C099B092",
-30434 => x"C0C0BFB0C099B099",
-30433 => x"C0C0BFB0C099B0B0",
-30432 => x"C0C0BFB0C099B0A4",
-30431 => x"C0C0BFB0C099B0F9",
-30430 => x"C0C0BFB0C099B0C0",
-30429 => x"C0C0BFB0C099A490",
-30428 => x"C0C0BFB0C099A480",
-30427 => x"C0C0BFB0C099A4F8",
-30426 => x"C0C0BFB0C099A482",
-30425 => x"C0C0BFB0C099A492",
-30424 => x"C0C0BFB0C099A499",
-30423 => x"C0C0BFB0C099A4B0",
-30422 => x"C0C0BFB0C099A4A4",
-30421 => x"C0C0BFB0C099A4F9",
-30420 => x"C0C0BFB0C099A4C0",
-30419 => x"C0C0BFB0C099F990",
-30418 => x"C0C0BFB0C099F980",
-30417 => x"C0C0BFB0C099F9F8",
-30416 => x"C0C0BFB0C099F982",
-30415 => x"C0C0BFB0C099F992",
-30414 => x"C0C0BFB0C099F999",
-30413 => x"C0C0BFB0C099F9B0",
-30412 => x"C0C0BFB0C099F9A4",
-30411 => x"C0C0BFB0C099F9F9",
-30410 => x"C0C0BFB0C099F9C0",
-30409 => x"C0C0BFB0C099C090",
-30408 => x"C0C0BFB0C099C080",
-30407 => x"C0C0BFB0C099C0F8",
-30406 => x"C0C0BFB0C099C082",
-30405 => x"C0C0BFB0C099C092",
-30404 => x"C0C0BFB0C099C099",
-30403 => x"C0C0BFB0C099C0B0",
-30402 => x"C0C0BFB0C099C0A4",
-30401 => x"C0C0BFB0C099C0F9",
-30400 => x"C0C0BFB0C099C0C0",
-30399 => x"C0C0BFB0C0B09090",
-30398 => x"C0C0BFB0C0B09080",
-30397 => x"C0C0BFB0C0B090F8",
-30396 => x"C0C0BFB0C0B09082",
-30395 => x"C0C0BFB0C0B09092",
-30394 => x"C0C0BFB0C0B09099",
-30393 => x"C0C0BFB0C0B090B0",
-30392 => x"C0C0BFB0C0B090A4",
-30391 => x"C0C0BFB0C0B090F9",
-30390 => x"C0C0BFB0C0B090C0",
-30389 => x"C0C0BFB0C0B08090",
-30388 => x"C0C0BFB0C0B08080",
-30387 => x"C0C0BFB0C0B080F8",
-30386 => x"C0C0BFB0C0B08082",
-30385 => x"C0C0BFB0C0B08092",
-30384 => x"C0C0BFB0C0B08099",
-30383 => x"C0C0BFB0C0B080B0",
-30382 => x"C0C0BFB0C0B080A4",
-30381 => x"C0C0BFB0C0B080F9",
-30380 => x"C0C0BFB0C0B080C0",
-30379 => x"C0C0BFB0C0B0F890",
-30378 => x"C0C0BFB0C0B0F880",
-30377 => x"C0C0BFB0C0B0F8F8",
-30376 => x"C0C0BFB0C0B0F882",
-30375 => x"C0C0BFB0C0B0F892",
-30374 => x"C0C0BFB0C0B0F899",
-30373 => x"C0C0BFB0C0B0F8B0",
-30372 => x"C0C0BFB0C0B0F8A4",
-30371 => x"C0C0BFB0C0B0F8F9",
-30370 => x"C0C0BFB0C0B0F8C0",
-30369 => x"C0C0BFB0C0B08290",
-30368 => x"C0C0BFB0C0B08280",
-30367 => x"C0C0BFB0C0B082F8",
-30366 => x"C0C0BFB0C0B08282",
-30365 => x"C0C0BFB0C0B08292",
-30364 => x"C0C0BFB0C0B08299",
-30363 => x"C0C0BFB0C0B082B0",
-30362 => x"C0C0BFB0C0B082A4",
-30361 => x"C0C0BFB0C0B082F9",
-30360 => x"C0C0BFB0C0B082C0",
-30359 => x"C0C0BFB0C0B09290",
-30358 => x"C0C0BFB0C0B09280",
-30357 => x"C0C0BFB0C0B092F8",
-30356 => x"C0C0BFB0C0B09282",
-30355 => x"C0C0BFB0C0B09292",
-30354 => x"C0C0BFB0C0B09299",
-30353 => x"C0C0BFB0C0B092B0",
-30352 => x"C0C0BFB0C0B092A4",
-30351 => x"C0C0BFB0C0B092F9",
-30350 => x"C0C0BFB0C0B092C0",
-30349 => x"C0C0BFB0C0B09990",
-30348 => x"C0C0BFB0C0B09980",
-30347 => x"C0C0BFB0C0B099F8",
-30346 => x"C0C0BFB0C0B09982",
-30345 => x"C0C0BFB0C0B09992",
-30344 => x"C0C0BFB0C0B09999",
-30343 => x"C0C0BFB0C0B099B0",
-30342 => x"C0C0BFB0C0B099A4",
-30341 => x"C0C0BFB0C0B099F9",
-30340 => x"C0C0BFB0C0B099C0",
-30339 => x"C0C0BFB0C0B0B090",
-30338 => x"C0C0BFB0C0B0B080",
-30337 => x"C0C0BFB0C0B0B0F8",
-30336 => x"C0C0BFB0C0B0B082",
-30335 => x"C0C0BFB0C0B0B092",
-30334 => x"C0C0BFB0C0B0B099",
-30333 => x"C0C0BFB0C0B0B0B0",
-30332 => x"C0C0BFB0C0B0B0A4",
-30331 => x"C0C0BFB0C0B0B0F9",
-30330 => x"C0C0BFB0C0B0B0C0",
-30329 => x"C0C0BFB0C0B0A490",
-30328 => x"C0C0BFB0C0B0A480",
-30327 => x"C0C0BFB0C0B0A4F8",
-30326 => x"C0C0BFB0C0B0A482",
-30325 => x"C0C0BFB0C0B0A492",
-30324 => x"C0C0BFB0C0B0A499",
-30323 => x"C0C0BFB0C0B0A4B0",
-30322 => x"C0C0BFB0C0B0A4A4",
-30321 => x"C0C0BFB0C0B0A4F9",
-30320 => x"C0C0BFB0C0B0A4C0",
-30319 => x"C0C0BFB0C0B0F990",
-30318 => x"C0C0BFB0C0B0F980",
-30317 => x"C0C0BFB0C0B0F9F8",
-30316 => x"C0C0BFB0C0B0F982",
-30315 => x"C0C0BFB0C0B0F992",
-30314 => x"C0C0BFB0C0B0F999",
-30313 => x"C0C0BFB0C0B0F9B0",
-30312 => x"C0C0BFB0C0B0F9A4",
-30311 => x"C0C0BFB0C0B0F9F9",
-30310 => x"C0C0BFB0C0B0F9C0",
-30309 => x"C0C0BFB0C0B0C090",
-30308 => x"C0C0BFB0C0B0C080",
-30307 => x"C0C0BFB0C0B0C0F8",
-30306 => x"C0C0BFB0C0B0C082",
-30305 => x"C0C0BFB0C0B0C092",
-30304 => x"C0C0BFB0C0B0C099",
-30303 => x"C0C0BFB0C0B0C0B0",
-30302 => x"C0C0BFB0C0B0C0A4",
-30301 => x"C0C0BFB0C0B0C0F9",
-30300 => x"C0C0BFB0C0B0C0C0",
-30299 => x"C0C0BFB0C0A49090",
-30298 => x"C0C0BFB0C0A49080",
-30297 => x"C0C0BFB0C0A490F8",
-30296 => x"C0C0BFB0C0A49082",
-30295 => x"C0C0BFB0C0A49092",
-30294 => x"C0C0BFB0C0A49099",
-30293 => x"C0C0BFB0C0A490B0",
-30292 => x"C0C0BFB0C0A490A4",
-30291 => x"C0C0BFB0C0A490F9",
-30290 => x"C0C0BFB0C0A490C0",
-30289 => x"C0C0BFB0C0A48090",
-30288 => x"C0C0BFB0C0A48080",
-30287 => x"C0C0BFB0C0A480F8",
-30286 => x"C0C0BFB0C0A48082",
-30285 => x"C0C0BFB0C0A48092",
-30284 => x"C0C0BFB0C0A48099",
-30283 => x"C0C0BFB0C0A480B0",
-30282 => x"C0C0BFB0C0A480A4",
-30281 => x"C0C0BFB0C0A480F9",
-30280 => x"C0C0BFB0C0A480C0",
-30279 => x"C0C0BFB0C0A4F890",
-30278 => x"C0C0BFB0C0A4F880",
-30277 => x"C0C0BFB0C0A4F8F8",
-30276 => x"C0C0BFB0C0A4F882",
-30275 => x"C0C0BFB0C0A4F892",
-30274 => x"C0C0BFB0C0A4F899",
-30273 => x"C0C0BFB0C0A4F8B0",
-30272 => x"C0C0BFB0C0A4F8A4",
-30271 => x"C0C0BFB0C0A4F8F9",
-30270 => x"C0C0BFB0C0A4F8C0",
-30269 => x"C0C0BFB0C0A48290",
-30268 => x"C0C0BFB0C0A48280",
-30267 => x"C0C0BFB0C0A482F8",
-30266 => x"C0C0BFB0C0A48282",
-30265 => x"C0C0BFB0C0A48292",
-30264 => x"C0C0BFB0C0A48299",
-30263 => x"C0C0BFB0C0A482B0",
-30262 => x"C0C0BFB0C0A482A4",
-30261 => x"C0C0BFB0C0A482F9",
-30260 => x"C0C0BFB0C0A482C0",
-30259 => x"C0C0BFB0C0A49290",
-30258 => x"C0C0BFB0C0A49280",
-30257 => x"C0C0BFB0C0A492F8",
-30256 => x"C0C0BFB0C0A49282",
-30255 => x"C0C0BFB0C0A49292",
-30254 => x"C0C0BFB0C0A49299",
-30253 => x"C0C0BFB0C0A492B0",
-30252 => x"C0C0BFB0C0A492A4",
-30251 => x"C0C0BFB0C0A492F9",
-30250 => x"C0C0BFB0C0A492C0",
-30249 => x"C0C0BFB0C0A49990",
-30248 => x"C0C0BFB0C0A49980",
-30247 => x"C0C0BFB0C0A499F8",
-30246 => x"C0C0BFB0C0A49982",
-30245 => x"C0C0BFB0C0A49992",
-30244 => x"C0C0BFB0C0A49999",
-30243 => x"C0C0BFB0C0A499B0",
-30242 => x"C0C0BFB0C0A499A4",
-30241 => x"C0C0BFB0C0A499F9",
-30240 => x"C0C0BFB0C0A499C0",
-30239 => x"C0C0BFB0C0A4B090",
-30238 => x"C0C0BFB0C0A4B080",
-30237 => x"C0C0BFB0C0A4B0F8",
-30236 => x"C0C0BFB0C0A4B082",
-30235 => x"C0C0BFB0C0A4B092",
-30234 => x"C0C0BFB0C0A4B099",
-30233 => x"C0C0BFB0C0A4B0B0",
-30232 => x"C0C0BFB0C0A4B0A4",
-30231 => x"C0C0BFB0C0A4B0F9",
-30230 => x"C0C0BFB0C0A4B0C0",
-30229 => x"C0C0BFB0C0A4A490",
-30228 => x"C0C0BFB0C0A4A480",
-30227 => x"C0C0BFB0C0A4A4F8",
-30226 => x"C0C0BFB0C0A4A482",
-30225 => x"C0C0BFB0C0A4A492",
-30224 => x"C0C0BFB0C0A4A499",
-30223 => x"C0C0BFB0C0A4A4B0",
-30222 => x"C0C0BFB0C0A4A4A4",
-30221 => x"C0C0BFB0C0A4A4F9",
-30220 => x"C0C0BFB0C0A4A4C0",
-30219 => x"C0C0BFB0C0A4F990",
-30218 => x"C0C0BFB0C0A4F980",
-30217 => x"C0C0BFB0C0A4F9F8",
-30216 => x"C0C0BFB0C0A4F982",
-30215 => x"C0C0BFB0C0A4F992",
-30214 => x"C0C0BFB0C0A4F999",
-30213 => x"C0C0BFB0C0A4F9B0",
-30212 => x"C0C0BFB0C0A4F9A4",
-30211 => x"C0C0BFB0C0A4F9F9",
-30210 => x"C0C0BFB0C0A4F9C0",
-30209 => x"C0C0BFB0C0A4C090",
-30208 => x"C0C0BFB0C0A4C080",
-30207 => x"C0C0BFB0C0A4C0F8",
-30206 => x"C0C0BFB0C0A4C082",
-30205 => x"C0C0BFB0C0A4C092",
-30204 => x"C0C0BFB0C0A4C099",
-30203 => x"C0C0BFB0C0A4C0B0",
-30202 => x"C0C0BFB0C0A4C0A4",
-30201 => x"C0C0BFB0C0A4C0F9",
-30200 => x"C0C0BFB0C0A4C0C0",
-30199 => x"C0C0BFB0C0F99090",
-30198 => x"C0C0BFB0C0F99080",
-30197 => x"C0C0BFB0C0F990F8",
-30196 => x"C0C0BFB0C0F99082",
-30195 => x"C0C0BFB0C0F99092",
-30194 => x"C0C0BFB0C0F99099",
-30193 => x"C0C0BFB0C0F990B0",
-30192 => x"C0C0BFB0C0F990A4",
-30191 => x"C0C0BFB0C0F990F9",
-30190 => x"C0C0BFB0C0F990C0",
-30189 => x"C0C0BFB0C0F98090",
-30188 => x"C0C0BFB0C0F98080",
-30187 => x"C0C0BFB0C0F980F8",
-30186 => x"C0C0BFB0C0F98082",
-30185 => x"C0C0BFB0C0F98092",
-30184 => x"C0C0BFB0C0F98099",
-30183 => x"C0C0BFB0C0F980B0",
-30182 => x"C0C0BFB0C0F980A4",
-30181 => x"C0C0BFB0C0F980F9",
-30180 => x"C0C0BFB0C0F980C0",
-30179 => x"C0C0BFB0C0F9F890",
-30178 => x"C0C0BFB0C0F9F880",
-30177 => x"C0C0BFB0C0F9F8F8",
-30176 => x"C0C0BFB0C0F9F882",
-30175 => x"C0C0BFB0C0F9F892",
-30174 => x"C0C0BFB0C0F9F899",
-30173 => x"C0C0BFB0C0F9F8B0",
-30172 => x"C0C0BFB0C0F9F8A4",
-30171 => x"C0C0BFB0C0F9F8F9",
-30170 => x"C0C0BFB0C0F9F8C0",
-30169 => x"C0C0BFB0C0F98290",
-30168 => x"C0C0BFB0C0F98280",
-30167 => x"C0C0BFB0C0F982F8",
-30166 => x"C0C0BFB0C0F98282",
-30165 => x"C0C0BFB0C0F98292",
-30164 => x"C0C0BFB0C0F98299",
-30163 => x"C0C0BFB0C0F982B0",
-30162 => x"C0C0BFB0C0F982A4",
-30161 => x"C0C0BFB0C0F982F9",
-30160 => x"C0C0BFB0C0F982C0",
-30159 => x"C0C0BFB0C0F99290",
-30158 => x"C0C0BFB0C0F99280",
-30157 => x"C0C0BFB0C0F992F8",
-30156 => x"C0C0BFB0C0F99282",
-30155 => x"C0C0BFB0C0F99292",
-30154 => x"C0C0BFB0C0F99299",
-30153 => x"C0C0BFB0C0F992B0",
-30152 => x"C0C0BFB0C0F992A4",
-30151 => x"C0C0BFB0C0F992F9",
-30150 => x"C0C0BFB0C0F992C0",
-30149 => x"C0C0BFB0C0F99990",
-30148 => x"C0C0BFB0C0F99980",
-30147 => x"C0C0BFB0C0F999F8",
-30146 => x"C0C0BFB0C0F99982",
-30145 => x"C0C0BFB0C0F99992",
-30144 => x"C0C0BFB0C0F99999",
-30143 => x"C0C0BFB0C0F999B0",
-30142 => x"C0C0BFB0C0F999A4",
-30141 => x"C0C0BFB0C0F999F9",
-30140 => x"C0C0BFB0C0F999C0",
-30139 => x"C0C0BFB0C0F9B090",
-30138 => x"C0C0BFB0C0F9B080",
-30137 => x"C0C0BFB0C0F9B0F8",
-30136 => x"C0C0BFB0C0F9B082",
-30135 => x"C0C0BFB0C0F9B092",
-30134 => x"C0C0BFB0C0F9B099",
-30133 => x"C0C0BFB0C0F9B0B0",
-30132 => x"C0C0BFB0C0F9B0A4",
-30131 => x"C0C0BFB0C0F9B0F9",
-30130 => x"C0C0BFB0C0F9B0C0",
-30129 => x"C0C0BFB0C0F9A490",
-30128 => x"C0C0BFB0C0F9A480",
-30127 => x"C0C0BFB0C0F9A4F8",
-30126 => x"C0C0BFB0C0F9A482",
-30125 => x"C0C0BFB0C0F9A492",
-30124 => x"C0C0BFB0C0F9A499",
-30123 => x"C0C0BFB0C0F9A4B0",
-30122 => x"C0C0BFB0C0F9A4A4",
-30121 => x"C0C0BFB0C0F9A4F9",
-30120 => x"C0C0BFB0C0F9A4C0",
-30119 => x"C0C0BFB0C0F9F990",
-30118 => x"C0C0BFB0C0F9F980",
-30117 => x"C0C0BFB0C0F9F9F8",
-30116 => x"C0C0BFB0C0F9F982",
-30115 => x"C0C0BFB0C0F9F992",
-30114 => x"C0C0BFB0C0F9F999",
-30113 => x"C0C0BFB0C0F9F9B0",
-30112 => x"C0C0BFB0C0F9F9A4",
-30111 => x"C0C0BFB0C0F9F9F9",
-30110 => x"C0C0BFB0C0F9F9C0",
-30109 => x"C0C0BFB0C0F9C090",
-30108 => x"C0C0BFB0C0F9C080",
-30107 => x"C0C0BFB0C0F9C0F8",
-30106 => x"C0C0BFB0C0F9C082",
-30105 => x"C0C0BFB0C0F9C092",
-30104 => x"C0C0BFB0C0F9C099",
-30103 => x"C0C0BFB0C0F9C0B0",
-30102 => x"C0C0BFB0C0F9C0A4",
-30101 => x"C0C0BFB0C0F9C0F9",
-30100 => x"C0C0BFB0C0F9C0C0",
-30099 => x"C0C0BFB0C0C09090",
-30098 => x"C0C0BFB0C0C09080",
-30097 => x"C0C0BFB0C0C090F8",
-30096 => x"C0C0BFB0C0C09082",
-30095 => x"C0C0BFB0C0C09092",
-30094 => x"C0C0BFB0C0C09099",
-30093 => x"C0C0BFB0C0C090B0",
-30092 => x"C0C0BFB0C0C090A4",
-30091 => x"C0C0BFB0C0C090F9",
-30090 => x"C0C0BFB0C0C090C0",
-30089 => x"C0C0BFB0C0C08090",
-30088 => x"C0C0BFB0C0C08080",
-30087 => x"C0C0BFB0C0C080F8",
-30086 => x"C0C0BFB0C0C08082",
-30085 => x"C0C0BFB0C0C08092",
-30084 => x"C0C0BFB0C0C08099",
-30083 => x"C0C0BFB0C0C080B0",
-30082 => x"C0C0BFB0C0C080A4",
-30081 => x"C0C0BFB0C0C080F9",
-30080 => x"C0C0BFB0C0C080C0",
-30079 => x"C0C0BFB0C0C0F890",
-30078 => x"C0C0BFB0C0C0F880",
-30077 => x"C0C0BFB0C0C0F8F8",
-30076 => x"C0C0BFB0C0C0F882",
-30075 => x"C0C0BFB0C0C0F892",
-30074 => x"C0C0BFB0C0C0F899",
-30073 => x"C0C0BFB0C0C0F8B0",
-30072 => x"C0C0BFB0C0C0F8A4",
-30071 => x"C0C0BFB0C0C0F8F9",
-30070 => x"C0C0BFB0C0C0F8C0",
-30069 => x"C0C0BFB0C0C08290",
-30068 => x"C0C0BFB0C0C08280",
-30067 => x"C0C0BFB0C0C082F8",
-30066 => x"C0C0BFB0C0C08282",
-30065 => x"C0C0BFB0C0C08292",
-30064 => x"C0C0BFB0C0C08299",
-30063 => x"C0C0BFB0C0C082B0",
-30062 => x"C0C0BFB0C0C082A4",
-30061 => x"C0C0BFB0C0C082F9",
-30060 => x"C0C0BFB0C0C082C0",
-30059 => x"C0C0BFB0C0C09290",
-30058 => x"C0C0BFB0C0C09280",
-30057 => x"C0C0BFB0C0C092F8",
-30056 => x"C0C0BFB0C0C09282",
-30055 => x"C0C0BFB0C0C09292",
-30054 => x"C0C0BFB0C0C09299",
-30053 => x"C0C0BFB0C0C092B0",
-30052 => x"C0C0BFB0C0C092A4",
-30051 => x"C0C0BFB0C0C092F9",
-30050 => x"C0C0BFB0C0C092C0",
-30049 => x"C0C0BFB0C0C09990",
-30048 => x"C0C0BFB0C0C09980",
-30047 => x"C0C0BFB0C0C099F8",
-30046 => x"C0C0BFB0C0C09982",
-30045 => x"C0C0BFB0C0C09992",
-30044 => x"C0C0BFB0C0C09999",
-30043 => x"C0C0BFB0C0C099B0",
-30042 => x"C0C0BFB0C0C099A4",
-30041 => x"C0C0BFB0C0C099F9",
-30040 => x"C0C0BFB0C0C099C0",
-30039 => x"C0C0BFB0C0C0B090",
-30038 => x"C0C0BFB0C0C0B080",
-30037 => x"C0C0BFB0C0C0B0F8",
-30036 => x"C0C0BFB0C0C0B082",
-30035 => x"C0C0BFB0C0C0B092",
-30034 => x"C0C0BFB0C0C0B099",
-30033 => x"C0C0BFB0C0C0B0B0",
-30032 => x"C0C0BFB0C0C0B0A4",
-30031 => x"C0C0BFB0C0C0B0F9",
-30030 => x"C0C0BFB0C0C0B0C0",
-30029 => x"C0C0BFB0C0C0A490",
-30028 => x"C0C0BFB0C0C0A480",
-30027 => x"C0C0BFB0C0C0A4F8",
-30026 => x"C0C0BFB0C0C0A482",
-30025 => x"C0C0BFB0C0C0A492",
-30024 => x"C0C0BFB0C0C0A499",
-30023 => x"C0C0BFB0C0C0A4B0",
-30022 => x"C0C0BFB0C0C0A4A4",
-30021 => x"C0C0BFB0C0C0A4F9",
-30020 => x"C0C0BFB0C0C0A4C0",
-30019 => x"C0C0BFB0C0C0F990",
-30018 => x"C0C0BFB0C0C0F980",
-30017 => x"C0C0BFB0C0C0F9F8",
-30016 => x"C0C0BFB0C0C0F982",
-30015 => x"C0C0BFB0C0C0F992",
-30014 => x"C0C0BFB0C0C0F999",
-30013 => x"C0C0BFB0C0C0F9B0",
-30012 => x"C0C0BFB0C0C0F9A4",
-30011 => x"C0C0BFB0C0C0F9F9",
-30010 => x"C0C0BFB0C0C0F9C0",
-30009 => x"C0C0BFB0C0C0C090",
-30008 => x"C0C0BFB0C0C0C080",
-30007 => x"C0C0BFB0C0C0C0F8",
-30006 => x"C0C0BFB0C0C0C082",
-30005 => x"C0C0BFB0C0C0C092",
-30004 => x"C0C0BFB0C0C0C099",
-30003 => x"C0C0BFB0C0C0C0B0",
-30002 => x"C0C0BFB0C0C0C0A4",
-30001 => x"C0C0BFB0C0C0C0F9",
-30000 => x"C0C0BFB0C0C0C0C0",
-29999 => x"C0C0BFA490909090",
-29998 => x"C0C0BFA490909080",
-29997 => x"C0C0BFA4909090F8",
-29996 => x"C0C0BFA490909082",
-29995 => x"C0C0BFA490909092",
-29994 => x"C0C0BFA490909099",
-29993 => x"C0C0BFA4909090B0",
-29992 => x"C0C0BFA4909090A4",
-29991 => x"C0C0BFA4909090F9",
-29990 => x"C0C0BFA4909090C0",
-29989 => x"C0C0BFA490908090",
-29988 => x"C0C0BFA490908080",
-29987 => x"C0C0BFA4909080F8",
-29986 => x"C0C0BFA490908082",
-29985 => x"C0C0BFA490908092",
-29984 => x"C0C0BFA490908099",
-29983 => x"C0C0BFA4909080B0",
-29982 => x"C0C0BFA4909080A4",
-29981 => x"C0C0BFA4909080F9",
-29980 => x"C0C0BFA4909080C0",
-29979 => x"C0C0BFA49090F890",
-29978 => x"C0C0BFA49090F880",
-29977 => x"C0C0BFA49090F8F8",
-29976 => x"C0C0BFA49090F882",
-29975 => x"C0C0BFA49090F892",
-29974 => x"C0C0BFA49090F899",
-29973 => x"C0C0BFA49090F8B0",
-29972 => x"C0C0BFA49090F8A4",
-29971 => x"C0C0BFA49090F8F9",
-29970 => x"C0C0BFA49090F8C0",
-29969 => x"C0C0BFA490908290",
-29968 => x"C0C0BFA490908280",
-29967 => x"C0C0BFA4909082F8",
-29966 => x"C0C0BFA490908282",
-29965 => x"C0C0BFA490908292",
-29964 => x"C0C0BFA490908299",
-29963 => x"C0C0BFA4909082B0",
-29962 => x"C0C0BFA4909082A4",
-29961 => x"C0C0BFA4909082F9",
-29960 => x"C0C0BFA4909082C0",
-29959 => x"C0C0BFA490909290",
-29958 => x"C0C0BFA490909280",
-29957 => x"C0C0BFA4909092F8",
-29956 => x"C0C0BFA490909282",
-29955 => x"C0C0BFA490909292",
-29954 => x"C0C0BFA490909299",
-29953 => x"C0C0BFA4909092B0",
-29952 => x"C0C0BFA4909092A4",
-29951 => x"C0C0BFA4909092F9",
-29950 => x"C0C0BFA4909092C0",
-29949 => x"C0C0BFA490909990",
-29948 => x"C0C0BFA490909980",
-29947 => x"C0C0BFA4909099F8",
-29946 => x"C0C0BFA490909982",
-29945 => x"C0C0BFA490909992",
-29944 => x"C0C0BFA490909999",
-29943 => x"C0C0BFA4909099B0",
-29942 => x"C0C0BFA4909099A4",
-29941 => x"C0C0BFA4909099F9",
-29940 => x"C0C0BFA4909099C0",
-29939 => x"C0C0BFA49090B090",
-29938 => x"C0C0BFA49090B080",
-29937 => x"C0C0BFA49090B0F8",
-29936 => x"C0C0BFA49090B082",
-29935 => x"C0C0BFA49090B092",
-29934 => x"C0C0BFA49090B099",
-29933 => x"C0C0BFA49090B0B0",
-29932 => x"C0C0BFA49090B0A4",
-29931 => x"C0C0BFA49090B0F9",
-29930 => x"C0C0BFA49090B0C0",
-29929 => x"C0C0BFA49090A490",
-29928 => x"C0C0BFA49090A480",
-29927 => x"C0C0BFA49090A4F8",
-29926 => x"C0C0BFA49090A482",
-29925 => x"C0C0BFA49090A492",
-29924 => x"C0C0BFA49090A499",
-29923 => x"C0C0BFA49090A4B0",
-29922 => x"C0C0BFA49090A4A4",
-29921 => x"C0C0BFA49090A4F9",
-29920 => x"C0C0BFA49090A4C0",
-29919 => x"C0C0BFA49090F990",
-29918 => x"C0C0BFA49090F980",
-29917 => x"C0C0BFA49090F9F8",
-29916 => x"C0C0BFA49090F982",
-29915 => x"C0C0BFA49090F992",
-29914 => x"C0C0BFA49090F999",
-29913 => x"C0C0BFA49090F9B0",
-29912 => x"C0C0BFA49090F9A4",
-29911 => x"C0C0BFA49090F9F9",
-29910 => x"C0C0BFA49090F9C0",
-29909 => x"C0C0BFA49090C090",
-29908 => x"C0C0BFA49090C080",
-29907 => x"C0C0BFA49090C0F8",
-29906 => x"C0C0BFA49090C082",
-29905 => x"C0C0BFA49090C092",
-29904 => x"C0C0BFA49090C099",
-29903 => x"C0C0BFA49090C0B0",
-29902 => x"C0C0BFA49090C0A4",
-29901 => x"C0C0BFA49090C0F9",
-29900 => x"C0C0BFA49090C0C0",
-29899 => x"C0C0BFA490809090",
-29898 => x"C0C0BFA490809080",
-29897 => x"C0C0BFA4908090F8",
-29896 => x"C0C0BFA490809082",
-29895 => x"C0C0BFA490809092",
-29894 => x"C0C0BFA490809099",
-29893 => x"C0C0BFA4908090B0",
-29892 => x"C0C0BFA4908090A4",
-29891 => x"C0C0BFA4908090F9",
-29890 => x"C0C0BFA4908090C0",
-29889 => x"C0C0BFA490808090",
-29888 => x"C0C0BFA490808080",
-29887 => x"C0C0BFA4908080F8",
-29886 => x"C0C0BFA490808082",
-29885 => x"C0C0BFA490808092",
-29884 => x"C0C0BFA490808099",
-29883 => x"C0C0BFA4908080B0",
-29882 => x"C0C0BFA4908080A4",
-29881 => x"C0C0BFA4908080F9",
-29880 => x"C0C0BFA4908080C0",
-29879 => x"C0C0BFA49080F890",
-29878 => x"C0C0BFA49080F880",
-29877 => x"C0C0BFA49080F8F8",
-29876 => x"C0C0BFA49080F882",
-29875 => x"C0C0BFA49080F892",
-29874 => x"C0C0BFA49080F899",
-29873 => x"C0C0BFA49080F8B0",
-29872 => x"C0C0BFA49080F8A4",
-29871 => x"C0C0BFA49080F8F9",
-29870 => x"C0C0BFA49080F8C0",
-29869 => x"C0C0BFA490808290",
-29868 => x"C0C0BFA490808280",
-29867 => x"C0C0BFA4908082F8",
-29866 => x"C0C0BFA490808282",
-29865 => x"C0C0BFA490808292",
-29864 => x"C0C0BFA490808299",
-29863 => x"C0C0BFA4908082B0",
-29862 => x"C0C0BFA4908082A4",
-29861 => x"C0C0BFA4908082F9",
-29860 => x"C0C0BFA4908082C0",
-29859 => x"C0C0BFA490809290",
-29858 => x"C0C0BFA490809280",
-29857 => x"C0C0BFA4908092F8",
-29856 => x"C0C0BFA490809282",
-29855 => x"C0C0BFA490809292",
-29854 => x"C0C0BFA490809299",
-29853 => x"C0C0BFA4908092B0",
-29852 => x"C0C0BFA4908092A4",
-29851 => x"C0C0BFA4908092F9",
-29850 => x"C0C0BFA4908092C0",
-29849 => x"C0C0BFA490809990",
-29848 => x"C0C0BFA490809980",
-29847 => x"C0C0BFA4908099F8",
-29846 => x"C0C0BFA490809982",
-29845 => x"C0C0BFA490809992",
-29844 => x"C0C0BFA490809999",
-29843 => x"C0C0BFA4908099B0",
-29842 => x"C0C0BFA4908099A4",
-29841 => x"C0C0BFA4908099F9",
-29840 => x"C0C0BFA4908099C0",
-29839 => x"C0C0BFA49080B090",
-29838 => x"C0C0BFA49080B080",
-29837 => x"C0C0BFA49080B0F8",
-29836 => x"C0C0BFA49080B082",
-29835 => x"C0C0BFA49080B092",
-29834 => x"C0C0BFA49080B099",
-29833 => x"C0C0BFA49080B0B0",
-29832 => x"C0C0BFA49080B0A4",
-29831 => x"C0C0BFA49080B0F9",
-29830 => x"C0C0BFA49080B0C0",
-29829 => x"C0C0BFA49080A490",
-29828 => x"C0C0BFA49080A480",
-29827 => x"C0C0BFA49080A4F8",
-29826 => x"C0C0BFA49080A482",
-29825 => x"C0C0BFA49080A492",
-29824 => x"C0C0BFA49080A499",
-29823 => x"C0C0BFA49080A4B0",
-29822 => x"C0C0BFA49080A4A4",
-29821 => x"C0C0BFA49080A4F9",
-29820 => x"C0C0BFA49080A4C0",
-29819 => x"C0C0BFA49080F990",
-29818 => x"C0C0BFA49080F980",
-29817 => x"C0C0BFA49080F9F8",
-29816 => x"C0C0BFA49080F982",
-29815 => x"C0C0BFA49080F992",
-29814 => x"C0C0BFA49080F999",
-29813 => x"C0C0BFA49080F9B0",
-29812 => x"C0C0BFA49080F9A4",
-29811 => x"C0C0BFA49080F9F9",
-29810 => x"C0C0BFA49080F9C0",
-29809 => x"C0C0BFA49080C090",
-29808 => x"C0C0BFA49080C080",
-29807 => x"C0C0BFA49080C0F8",
-29806 => x"C0C0BFA49080C082",
-29805 => x"C0C0BFA49080C092",
-29804 => x"C0C0BFA49080C099",
-29803 => x"C0C0BFA49080C0B0",
-29802 => x"C0C0BFA49080C0A4",
-29801 => x"C0C0BFA49080C0F9",
-29800 => x"C0C0BFA49080C0C0",
-29799 => x"C0C0BFA490F89090",
-29798 => x"C0C0BFA490F89080",
-29797 => x"C0C0BFA490F890F8",
-29796 => x"C0C0BFA490F89082",
-29795 => x"C0C0BFA490F89092",
-29794 => x"C0C0BFA490F89099",
-29793 => x"C0C0BFA490F890B0",
-29792 => x"C0C0BFA490F890A4",
-29791 => x"C0C0BFA490F890F9",
-29790 => x"C0C0BFA490F890C0",
-29789 => x"C0C0BFA490F88090",
-29788 => x"C0C0BFA490F88080",
-29787 => x"C0C0BFA490F880F8",
-29786 => x"C0C0BFA490F88082",
-29785 => x"C0C0BFA490F88092",
-29784 => x"C0C0BFA490F88099",
-29783 => x"C0C0BFA490F880B0",
-29782 => x"C0C0BFA490F880A4",
-29781 => x"C0C0BFA490F880F9",
-29780 => x"C0C0BFA490F880C0",
-29779 => x"C0C0BFA490F8F890",
-29778 => x"C0C0BFA490F8F880",
-29777 => x"C0C0BFA490F8F8F8",
-29776 => x"C0C0BFA490F8F882",
-29775 => x"C0C0BFA490F8F892",
-29774 => x"C0C0BFA490F8F899",
-29773 => x"C0C0BFA490F8F8B0",
-29772 => x"C0C0BFA490F8F8A4",
-29771 => x"C0C0BFA490F8F8F9",
-29770 => x"C0C0BFA490F8F8C0",
-29769 => x"C0C0BFA490F88290",
-29768 => x"C0C0BFA490F88280",
-29767 => x"C0C0BFA490F882F8",
-29766 => x"C0C0BFA490F88282",
-29765 => x"C0C0BFA490F88292",
-29764 => x"C0C0BFA490F88299",
-29763 => x"C0C0BFA490F882B0",
-29762 => x"C0C0BFA490F882A4",
-29761 => x"C0C0BFA490F882F9",
-29760 => x"C0C0BFA490F882C0",
-29759 => x"C0C0BFA490F89290",
-29758 => x"C0C0BFA490F89280",
-29757 => x"C0C0BFA490F892F8",
-29756 => x"C0C0BFA490F89282",
-29755 => x"C0C0BFA490F89292",
-29754 => x"C0C0BFA490F89299",
-29753 => x"C0C0BFA490F892B0",
-29752 => x"C0C0BFA490F892A4",
-29751 => x"C0C0BFA490F892F9",
-29750 => x"C0C0BFA490F892C0",
-29749 => x"C0C0BFA490F89990",
-29748 => x"C0C0BFA490F89980",
-29747 => x"C0C0BFA490F899F8",
-29746 => x"C0C0BFA490F89982",
-29745 => x"C0C0BFA490F89992",
-29744 => x"C0C0BFA490F89999",
-29743 => x"C0C0BFA490F899B0",
-29742 => x"C0C0BFA490F899A4",
-29741 => x"C0C0BFA490F899F9",
-29740 => x"C0C0BFA490F899C0",
-29739 => x"C0C0BFA490F8B090",
-29738 => x"C0C0BFA490F8B080",
-29737 => x"C0C0BFA490F8B0F8",
-29736 => x"C0C0BFA490F8B082",
-29735 => x"C0C0BFA490F8B092",
-29734 => x"C0C0BFA490F8B099",
-29733 => x"C0C0BFA490F8B0B0",
-29732 => x"C0C0BFA490F8B0A4",
-29731 => x"C0C0BFA490F8B0F9",
-29730 => x"C0C0BFA490F8B0C0",
-29729 => x"C0C0BFA490F8A490",
-29728 => x"C0C0BFA490F8A480",
-29727 => x"C0C0BFA490F8A4F8",
-29726 => x"C0C0BFA490F8A482",
-29725 => x"C0C0BFA490F8A492",
-29724 => x"C0C0BFA490F8A499",
-29723 => x"C0C0BFA490F8A4B0",
-29722 => x"C0C0BFA490F8A4A4",
-29721 => x"C0C0BFA490F8A4F9",
-29720 => x"C0C0BFA490F8A4C0",
-29719 => x"C0C0BFA490F8F990",
-29718 => x"C0C0BFA490F8F980",
-29717 => x"C0C0BFA490F8F9F8",
-29716 => x"C0C0BFA490F8F982",
-29715 => x"C0C0BFA490F8F992",
-29714 => x"C0C0BFA490F8F999",
-29713 => x"C0C0BFA490F8F9B0",
-29712 => x"C0C0BFA490F8F9A4",
-29711 => x"C0C0BFA490F8F9F9",
-29710 => x"C0C0BFA490F8F9C0",
-29709 => x"C0C0BFA490F8C090",
-29708 => x"C0C0BFA490F8C080",
-29707 => x"C0C0BFA490F8C0F8",
-29706 => x"C0C0BFA490F8C082",
-29705 => x"C0C0BFA490F8C092",
-29704 => x"C0C0BFA490F8C099",
-29703 => x"C0C0BFA490F8C0B0",
-29702 => x"C0C0BFA490F8C0A4",
-29701 => x"C0C0BFA490F8C0F9",
-29700 => x"C0C0BFA490F8C0C0",
-29699 => x"C0C0BFA490829090",
-29698 => x"C0C0BFA490829080",
-29697 => x"C0C0BFA4908290F8",
-29696 => x"C0C0BFA490829082",
-29695 => x"C0C0BFA490829092",
-29694 => x"C0C0BFA490829099",
-29693 => x"C0C0BFA4908290B0",
-29692 => x"C0C0BFA4908290A4",
-29691 => x"C0C0BFA4908290F9",
-29690 => x"C0C0BFA4908290C0",
-29689 => x"C0C0BFA490828090",
-29688 => x"C0C0BFA490828080",
-29687 => x"C0C0BFA4908280F8",
-29686 => x"C0C0BFA490828082",
-29685 => x"C0C0BFA490828092",
-29684 => x"C0C0BFA490828099",
-29683 => x"C0C0BFA4908280B0",
-29682 => x"C0C0BFA4908280A4",
-29681 => x"C0C0BFA4908280F9",
-29680 => x"C0C0BFA4908280C0",
-29679 => x"C0C0BFA49082F890",
-29678 => x"C0C0BFA49082F880",
-29677 => x"C0C0BFA49082F8F8",
-29676 => x"C0C0BFA49082F882",
-29675 => x"C0C0BFA49082F892",
-29674 => x"C0C0BFA49082F899",
-29673 => x"C0C0BFA49082F8B0",
-29672 => x"C0C0BFA49082F8A4",
-29671 => x"C0C0BFA49082F8F9",
-29670 => x"C0C0BFA49082F8C0",
-29669 => x"C0C0BFA490828290",
-29668 => x"C0C0BFA490828280",
-29667 => x"C0C0BFA4908282F8",
-29666 => x"C0C0BFA490828282",
-29665 => x"C0C0BFA490828292",
-29664 => x"C0C0BFA490828299",
-29663 => x"C0C0BFA4908282B0",
-29662 => x"C0C0BFA4908282A4",
-29661 => x"C0C0BFA4908282F9",
-29660 => x"C0C0BFA4908282C0",
-29659 => x"C0C0BFA490829290",
-29658 => x"C0C0BFA490829280",
-29657 => x"C0C0BFA4908292F8",
-29656 => x"C0C0BFA490829282",
-29655 => x"C0C0BFA490829292",
-29654 => x"C0C0BFA490829299",
-29653 => x"C0C0BFA4908292B0",
-29652 => x"C0C0BFA4908292A4",
-29651 => x"C0C0BFA4908292F9",
-29650 => x"C0C0BFA4908292C0",
-29649 => x"C0C0BFA490829990",
-29648 => x"C0C0BFA490829980",
-29647 => x"C0C0BFA4908299F8",
-29646 => x"C0C0BFA490829982",
-29645 => x"C0C0BFA490829992",
-29644 => x"C0C0BFA490829999",
-29643 => x"C0C0BFA4908299B0",
-29642 => x"C0C0BFA4908299A4",
-29641 => x"C0C0BFA4908299F9",
-29640 => x"C0C0BFA4908299C0",
-29639 => x"C0C0BFA49082B090",
-29638 => x"C0C0BFA49082B080",
-29637 => x"C0C0BFA49082B0F8",
-29636 => x"C0C0BFA49082B082",
-29635 => x"C0C0BFA49082B092",
-29634 => x"C0C0BFA49082B099",
-29633 => x"C0C0BFA49082B0B0",
-29632 => x"C0C0BFA49082B0A4",
-29631 => x"C0C0BFA49082B0F9",
-29630 => x"C0C0BFA49082B0C0",
-29629 => x"C0C0BFA49082A490",
-29628 => x"C0C0BFA49082A480",
-29627 => x"C0C0BFA49082A4F8",
-29626 => x"C0C0BFA49082A482",
-29625 => x"C0C0BFA49082A492",
-29624 => x"C0C0BFA49082A499",
-29623 => x"C0C0BFA49082A4B0",
-29622 => x"C0C0BFA49082A4A4",
-29621 => x"C0C0BFA49082A4F9",
-29620 => x"C0C0BFA49082A4C0",
-29619 => x"C0C0BFA49082F990",
-29618 => x"C0C0BFA49082F980",
-29617 => x"C0C0BFA49082F9F8",
-29616 => x"C0C0BFA49082F982",
-29615 => x"C0C0BFA49082F992",
-29614 => x"C0C0BFA49082F999",
-29613 => x"C0C0BFA49082F9B0",
-29612 => x"C0C0BFA49082F9A4",
-29611 => x"C0C0BFA49082F9F9",
-29610 => x"C0C0BFA49082F9C0",
-29609 => x"C0C0BFA49082C090",
-29608 => x"C0C0BFA49082C080",
-29607 => x"C0C0BFA49082C0F8",
-29606 => x"C0C0BFA49082C082",
-29605 => x"C0C0BFA49082C092",
-29604 => x"C0C0BFA49082C099",
-29603 => x"C0C0BFA49082C0B0",
-29602 => x"C0C0BFA49082C0A4",
-29601 => x"C0C0BFA49082C0F9",
-29600 => x"C0C0BFA49082C0C0",
-29599 => x"C0C0BFA490929090",
-29598 => x"C0C0BFA490929080",
-29597 => x"C0C0BFA4909290F8",
-29596 => x"C0C0BFA490929082",
-29595 => x"C0C0BFA490929092",
-29594 => x"C0C0BFA490929099",
-29593 => x"C0C0BFA4909290B0",
-29592 => x"C0C0BFA4909290A4",
-29591 => x"C0C0BFA4909290F9",
-29590 => x"C0C0BFA4909290C0",
-29589 => x"C0C0BFA490928090",
-29588 => x"C0C0BFA490928080",
-29587 => x"C0C0BFA4909280F8",
-29586 => x"C0C0BFA490928082",
-29585 => x"C0C0BFA490928092",
-29584 => x"C0C0BFA490928099",
-29583 => x"C0C0BFA4909280B0",
-29582 => x"C0C0BFA4909280A4",
-29581 => x"C0C0BFA4909280F9",
-29580 => x"C0C0BFA4909280C0",
-29579 => x"C0C0BFA49092F890",
-29578 => x"C0C0BFA49092F880",
-29577 => x"C0C0BFA49092F8F8",
-29576 => x"C0C0BFA49092F882",
-29575 => x"C0C0BFA49092F892",
-29574 => x"C0C0BFA49092F899",
-29573 => x"C0C0BFA49092F8B0",
-29572 => x"C0C0BFA49092F8A4",
-29571 => x"C0C0BFA49092F8F9",
-29570 => x"C0C0BFA49092F8C0",
-29569 => x"C0C0BFA490928290",
-29568 => x"C0C0BFA490928280",
-29567 => x"C0C0BFA4909282F8",
-29566 => x"C0C0BFA490928282",
-29565 => x"C0C0BFA490928292",
-29564 => x"C0C0BFA490928299",
-29563 => x"C0C0BFA4909282B0",
-29562 => x"C0C0BFA4909282A4",
-29561 => x"C0C0BFA4909282F9",
-29560 => x"C0C0BFA4909282C0",
-29559 => x"C0C0BFA490929290",
-29558 => x"C0C0BFA490929280",
-29557 => x"C0C0BFA4909292F8",
-29556 => x"C0C0BFA490929282",
-29555 => x"C0C0BFA490929292",
-29554 => x"C0C0BFA490929299",
-29553 => x"C0C0BFA4909292B0",
-29552 => x"C0C0BFA4909292A4",
-29551 => x"C0C0BFA4909292F9",
-29550 => x"C0C0BFA4909292C0",
-29549 => x"C0C0BFA490929990",
-29548 => x"C0C0BFA490929980",
-29547 => x"C0C0BFA4909299F8",
-29546 => x"C0C0BFA490929982",
-29545 => x"C0C0BFA490929992",
-29544 => x"C0C0BFA490929999",
-29543 => x"C0C0BFA4909299B0",
-29542 => x"C0C0BFA4909299A4",
-29541 => x"C0C0BFA4909299F9",
-29540 => x"C0C0BFA4909299C0",
-29539 => x"C0C0BFA49092B090",
-29538 => x"C0C0BFA49092B080",
-29537 => x"C0C0BFA49092B0F8",
-29536 => x"C0C0BFA49092B082",
-29535 => x"C0C0BFA49092B092",
-29534 => x"C0C0BFA49092B099",
-29533 => x"C0C0BFA49092B0B0",
-29532 => x"C0C0BFA49092B0A4",
-29531 => x"C0C0BFA49092B0F9",
-29530 => x"C0C0BFA49092B0C0",
-29529 => x"C0C0BFA49092A490",
-29528 => x"C0C0BFA49092A480",
-29527 => x"C0C0BFA49092A4F8",
-29526 => x"C0C0BFA49092A482",
-29525 => x"C0C0BFA49092A492",
-29524 => x"C0C0BFA49092A499",
-29523 => x"C0C0BFA49092A4B0",
-29522 => x"C0C0BFA49092A4A4",
-29521 => x"C0C0BFA49092A4F9",
-29520 => x"C0C0BFA49092A4C0",
-29519 => x"C0C0BFA49092F990",
-29518 => x"C0C0BFA49092F980",
-29517 => x"C0C0BFA49092F9F8",
-29516 => x"C0C0BFA49092F982",
-29515 => x"C0C0BFA49092F992",
-29514 => x"C0C0BFA49092F999",
-29513 => x"C0C0BFA49092F9B0",
-29512 => x"C0C0BFA49092F9A4",
-29511 => x"C0C0BFA49092F9F9",
-29510 => x"C0C0BFA49092F9C0",
-29509 => x"C0C0BFA49092C090",
-29508 => x"C0C0BFA49092C080",
-29507 => x"C0C0BFA49092C0F8",
-29506 => x"C0C0BFA49092C082",
-29505 => x"C0C0BFA49092C092",
-29504 => x"C0C0BFA49092C099",
-29503 => x"C0C0BFA49092C0B0",
-29502 => x"C0C0BFA49092C0A4",
-29501 => x"C0C0BFA49092C0F9",
-29500 => x"C0C0BFA49092C0C0",
-29499 => x"C0C0BFA490999090",
-29498 => x"C0C0BFA490999080",
-29497 => x"C0C0BFA4909990F8",
-29496 => x"C0C0BFA490999082",
-29495 => x"C0C0BFA490999092",
-29494 => x"C0C0BFA490999099",
-29493 => x"C0C0BFA4909990B0",
-29492 => x"C0C0BFA4909990A4",
-29491 => x"C0C0BFA4909990F9",
-29490 => x"C0C0BFA4909990C0",
-29489 => x"C0C0BFA490998090",
-29488 => x"C0C0BFA490998080",
-29487 => x"C0C0BFA4909980F8",
-29486 => x"C0C0BFA490998082",
-29485 => x"C0C0BFA490998092",
-29484 => x"C0C0BFA490998099",
-29483 => x"C0C0BFA4909980B0",
-29482 => x"C0C0BFA4909980A4",
-29481 => x"C0C0BFA4909980F9",
-29480 => x"C0C0BFA4909980C0",
-29479 => x"C0C0BFA49099F890",
-29478 => x"C0C0BFA49099F880",
-29477 => x"C0C0BFA49099F8F8",
-29476 => x"C0C0BFA49099F882",
-29475 => x"C0C0BFA49099F892",
-29474 => x"C0C0BFA49099F899",
-29473 => x"C0C0BFA49099F8B0",
-29472 => x"C0C0BFA49099F8A4",
-29471 => x"C0C0BFA49099F8F9",
-29470 => x"C0C0BFA49099F8C0",
-29469 => x"C0C0BFA490998290",
-29468 => x"C0C0BFA490998280",
-29467 => x"C0C0BFA4909982F8",
-29466 => x"C0C0BFA490998282",
-29465 => x"C0C0BFA490998292",
-29464 => x"C0C0BFA490998299",
-29463 => x"C0C0BFA4909982B0",
-29462 => x"C0C0BFA4909982A4",
-29461 => x"C0C0BFA4909982F9",
-29460 => x"C0C0BFA4909982C0",
-29459 => x"C0C0BFA490999290",
-29458 => x"C0C0BFA490999280",
-29457 => x"C0C0BFA4909992F8",
-29456 => x"C0C0BFA490999282",
-29455 => x"C0C0BFA490999292",
-29454 => x"C0C0BFA490999299",
-29453 => x"C0C0BFA4909992B0",
-29452 => x"C0C0BFA4909992A4",
-29451 => x"C0C0BFA4909992F9",
-29450 => x"C0C0BFA4909992C0",
-29449 => x"C0C0BFA490999990",
-29448 => x"C0C0BFA490999980",
-29447 => x"C0C0BFA4909999F8",
-29446 => x"C0C0BFA490999982",
-29445 => x"C0C0BFA490999992",
-29444 => x"C0C0BFA490999999",
-29443 => x"C0C0BFA4909999B0",
-29442 => x"C0C0BFA4909999A4",
-29441 => x"C0C0BFA4909999F9",
-29440 => x"C0C0BFA4909999C0",
-29439 => x"C0C0BFA49099B090",
-29438 => x"C0C0BFA49099B080",
-29437 => x"C0C0BFA49099B0F8",
-29436 => x"C0C0BFA49099B082",
-29435 => x"C0C0BFA49099B092",
-29434 => x"C0C0BFA49099B099",
-29433 => x"C0C0BFA49099B0B0",
-29432 => x"C0C0BFA49099B0A4",
-29431 => x"C0C0BFA49099B0F9",
-29430 => x"C0C0BFA49099B0C0",
-29429 => x"C0C0BFA49099A490",
-29428 => x"C0C0BFA49099A480",
-29427 => x"C0C0BFA49099A4F8",
-29426 => x"C0C0BFA49099A482",
-29425 => x"C0C0BFA49099A492",
-29424 => x"C0C0BFA49099A499",
-29423 => x"C0C0BFA49099A4B0",
-29422 => x"C0C0BFA49099A4A4",
-29421 => x"C0C0BFA49099A4F9",
-29420 => x"C0C0BFA49099A4C0",
-29419 => x"C0C0BFA49099F990",
-29418 => x"C0C0BFA49099F980",
-29417 => x"C0C0BFA49099F9F8",
-29416 => x"C0C0BFA49099F982",
-29415 => x"C0C0BFA49099F992",
-29414 => x"C0C0BFA49099F999",
-29413 => x"C0C0BFA49099F9B0",
-29412 => x"C0C0BFA49099F9A4",
-29411 => x"C0C0BFA49099F9F9",
-29410 => x"C0C0BFA49099F9C0",
-29409 => x"C0C0BFA49099C090",
-29408 => x"C0C0BFA49099C080",
-29407 => x"C0C0BFA49099C0F8",
-29406 => x"C0C0BFA49099C082",
-29405 => x"C0C0BFA49099C092",
-29404 => x"C0C0BFA49099C099",
-29403 => x"C0C0BFA49099C0B0",
-29402 => x"C0C0BFA49099C0A4",
-29401 => x"C0C0BFA49099C0F9",
-29400 => x"C0C0BFA49099C0C0",
-29399 => x"C0C0BFA490B09090",
-29398 => x"C0C0BFA490B09080",
-29397 => x"C0C0BFA490B090F8",
-29396 => x"C0C0BFA490B09082",
-29395 => x"C0C0BFA490B09092",
-29394 => x"C0C0BFA490B09099",
-29393 => x"C0C0BFA490B090B0",
-29392 => x"C0C0BFA490B090A4",
-29391 => x"C0C0BFA490B090F9",
-29390 => x"C0C0BFA490B090C0",
-29389 => x"C0C0BFA490B08090",
-29388 => x"C0C0BFA490B08080",
-29387 => x"C0C0BFA490B080F8",
-29386 => x"C0C0BFA490B08082",
-29385 => x"C0C0BFA490B08092",
-29384 => x"C0C0BFA490B08099",
-29383 => x"C0C0BFA490B080B0",
-29382 => x"C0C0BFA490B080A4",
-29381 => x"C0C0BFA490B080F9",
-29380 => x"C0C0BFA490B080C0",
-29379 => x"C0C0BFA490B0F890",
-29378 => x"C0C0BFA490B0F880",
-29377 => x"C0C0BFA490B0F8F8",
-29376 => x"C0C0BFA490B0F882",
-29375 => x"C0C0BFA490B0F892",
-29374 => x"C0C0BFA490B0F899",
-29373 => x"C0C0BFA490B0F8B0",
-29372 => x"C0C0BFA490B0F8A4",
-29371 => x"C0C0BFA490B0F8F9",
-29370 => x"C0C0BFA490B0F8C0",
-29369 => x"C0C0BFA490B08290",
-29368 => x"C0C0BFA490B08280",
-29367 => x"C0C0BFA490B082F8",
-29366 => x"C0C0BFA490B08282",
-29365 => x"C0C0BFA490B08292",
-29364 => x"C0C0BFA490B08299",
-29363 => x"C0C0BFA490B082B0",
-29362 => x"C0C0BFA490B082A4",
-29361 => x"C0C0BFA490B082F9",
-29360 => x"C0C0BFA490B082C0",
-29359 => x"C0C0BFA490B09290",
-29358 => x"C0C0BFA490B09280",
-29357 => x"C0C0BFA490B092F8",
-29356 => x"C0C0BFA490B09282",
-29355 => x"C0C0BFA490B09292",
-29354 => x"C0C0BFA490B09299",
-29353 => x"C0C0BFA490B092B0",
-29352 => x"C0C0BFA490B092A4",
-29351 => x"C0C0BFA490B092F9",
-29350 => x"C0C0BFA490B092C0",
-29349 => x"C0C0BFA490B09990",
-29348 => x"C0C0BFA490B09980",
-29347 => x"C0C0BFA490B099F8",
-29346 => x"C0C0BFA490B09982",
-29345 => x"C0C0BFA490B09992",
-29344 => x"C0C0BFA490B09999",
-29343 => x"C0C0BFA490B099B0",
-29342 => x"C0C0BFA490B099A4",
-29341 => x"C0C0BFA490B099F9",
-29340 => x"C0C0BFA490B099C0",
-29339 => x"C0C0BFA490B0B090",
-29338 => x"C0C0BFA490B0B080",
-29337 => x"C0C0BFA490B0B0F8",
-29336 => x"C0C0BFA490B0B082",
-29335 => x"C0C0BFA490B0B092",
-29334 => x"C0C0BFA490B0B099",
-29333 => x"C0C0BFA490B0B0B0",
-29332 => x"C0C0BFA490B0B0A4",
-29331 => x"C0C0BFA490B0B0F9",
-29330 => x"C0C0BFA490B0B0C0",
-29329 => x"C0C0BFA490B0A490",
-29328 => x"C0C0BFA490B0A480",
-29327 => x"C0C0BFA490B0A4F8",
-29326 => x"C0C0BFA490B0A482",
-29325 => x"C0C0BFA490B0A492",
-29324 => x"C0C0BFA490B0A499",
-29323 => x"C0C0BFA490B0A4B0",
-29322 => x"C0C0BFA490B0A4A4",
-29321 => x"C0C0BFA490B0A4F9",
-29320 => x"C0C0BFA490B0A4C0",
-29319 => x"C0C0BFA490B0F990",
-29318 => x"C0C0BFA490B0F980",
-29317 => x"C0C0BFA490B0F9F8",
-29316 => x"C0C0BFA490B0F982",
-29315 => x"C0C0BFA490B0F992",
-29314 => x"C0C0BFA490B0F999",
-29313 => x"C0C0BFA490B0F9B0",
-29312 => x"C0C0BFA490B0F9A4",
-29311 => x"C0C0BFA490B0F9F9",
-29310 => x"C0C0BFA490B0F9C0",
-29309 => x"C0C0BFA490B0C090",
-29308 => x"C0C0BFA490B0C080",
-29307 => x"C0C0BFA490B0C0F8",
-29306 => x"C0C0BFA490B0C082",
-29305 => x"C0C0BFA490B0C092",
-29304 => x"C0C0BFA490B0C099",
-29303 => x"C0C0BFA490B0C0B0",
-29302 => x"C0C0BFA490B0C0A4",
-29301 => x"C0C0BFA490B0C0F9",
-29300 => x"C0C0BFA490B0C0C0",
-29299 => x"C0C0BFA490A49090",
-29298 => x"C0C0BFA490A49080",
-29297 => x"C0C0BFA490A490F8",
-29296 => x"C0C0BFA490A49082",
-29295 => x"C0C0BFA490A49092",
-29294 => x"C0C0BFA490A49099",
-29293 => x"C0C0BFA490A490B0",
-29292 => x"C0C0BFA490A490A4",
-29291 => x"C0C0BFA490A490F9",
-29290 => x"C0C0BFA490A490C0",
-29289 => x"C0C0BFA490A48090",
-29288 => x"C0C0BFA490A48080",
-29287 => x"C0C0BFA490A480F8",
-29286 => x"C0C0BFA490A48082",
-29285 => x"C0C0BFA490A48092",
-29284 => x"C0C0BFA490A48099",
-29283 => x"C0C0BFA490A480B0",
-29282 => x"C0C0BFA490A480A4",
-29281 => x"C0C0BFA490A480F9",
-29280 => x"C0C0BFA490A480C0",
-29279 => x"C0C0BFA490A4F890",
-29278 => x"C0C0BFA490A4F880",
-29277 => x"C0C0BFA490A4F8F8",
-29276 => x"C0C0BFA490A4F882",
-29275 => x"C0C0BFA490A4F892",
-29274 => x"C0C0BFA490A4F899",
-29273 => x"C0C0BFA490A4F8B0",
-29272 => x"C0C0BFA490A4F8A4",
-29271 => x"C0C0BFA490A4F8F9",
-29270 => x"C0C0BFA490A4F8C0",
-29269 => x"C0C0BFA490A48290",
-29268 => x"C0C0BFA490A48280",
-29267 => x"C0C0BFA490A482F8",
-29266 => x"C0C0BFA490A48282",
-29265 => x"C0C0BFA490A48292",
-29264 => x"C0C0BFA490A48299",
-29263 => x"C0C0BFA490A482B0",
-29262 => x"C0C0BFA490A482A4",
-29261 => x"C0C0BFA490A482F9",
-29260 => x"C0C0BFA490A482C0",
-29259 => x"C0C0BFA490A49290",
-29258 => x"C0C0BFA490A49280",
-29257 => x"C0C0BFA490A492F8",
-29256 => x"C0C0BFA490A49282",
-29255 => x"C0C0BFA490A49292",
-29254 => x"C0C0BFA490A49299",
-29253 => x"C0C0BFA490A492B0",
-29252 => x"C0C0BFA490A492A4",
-29251 => x"C0C0BFA490A492F9",
-29250 => x"C0C0BFA490A492C0",
-29249 => x"C0C0BFA490A49990",
-29248 => x"C0C0BFA490A49980",
-29247 => x"C0C0BFA490A499F8",
-29246 => x"C0C0BFA490A49982",
-29245 => x"C0C0BFA490A49992",
-29244 => x"C0C0BFA490A49999",
-29243 => x"C0C0BFA490A499B0",
-29242 => x"C0C0BFA490A499A4",
-29241 => x"C0C0BFA490A499F9",
-29240 => x"C0C0BFA490A499C0",
-29239 => x"C0C0BFA490A4B090",
-29238 => x"C0C0BFA490A4B080",
-29237 => x"C0C0BFA490A4B0F8",
-29236 => x"C0C0BFA490A4B082",
-29235 => x"C0C0BFA490A4B092",
-29234 => x"C0C0BFA490A4B099",
-29233 => x"C0C0BFA490A4B0B0",
-29232 => x"C0C0BFA490A4B0A4",
-29231 => x"C0C0BFA490A4B0F9",
-29230 => x"C0C0BFA490A4B0C0",
-29229 => x"C0C0BFA490A4A490",
-29228 => x"C0C0BFA490A4A480",
-29227 => x"C0C0BFA490A4A4F8",
-29226 => x"C0C0BFA490A4A482",
-29225 => x"C0C0BFA490A4A492",
-29224 => x"C0C0BFA490A4A499",
-29223 => x"C0C0BFA490A4A4B0",
-29222 => x"C0C0BFA490A4A4A4",
-29221 => x"C0C0BFA490A4A4F9",
-29220 => x"C0C0BFA490A4A4C0",
-29219 => x"C0C0BFA490A4F990",
-29218 => x"C0C0BFA490A4F980",
-29217 => x"C0C0BFA490A4F9F8",
-29216 => x"C0C0BFA490A4F982",
-29215 => x"C0C0BFA490A4F992",
-29214 => x"C0C0BFA490A4F999",
-29213 => x"C0C0BFA490A4F9B0",
-29212 => x"C0C0BFA490A4F9A4",
-29211 => x"C0C0BFA490A4F9F9",
-29210 => x"C0C0BFA490A4F9C0",
-29209 => x"C0C0BFA490A4C090",
-29208 => x"C0C0BFA490A4C080",
-29207 => x"C0C0BFA490A4C0F8",
-29206 => x"C0C0BFA490A4C082",
-29205 => x"C0C0BFA490A4C092",
-29204 => x"C0C0BFA490A4C099",
-29203 => x"C0C0BFA490A4C0B0",
-29202 => x"C0C0BFA490A4C0A4",
-29201 => x"C0C0BFA490A4C0F9",
-29200 => x"C0C0BFA490A4C0C0",
-29199 => x"C0C0BFA490F99090",
-29198 => x"C0C0BFA490F99080",
-29197 => x"C0C0BFA490F990F8",
-29196 => x"C0C0BFA490F99082",
-29195 => x"C0C0BFA490F99092",
-29194 => x"C0C0BFA490F99099",
-29193 => x"C0C0BFA490F990B0",
-29192 => x"C0C0BFA490F990A4",
-29191 => x"C0C0BFA490F990F9",
-29190 => x"C0C0BFA490F990C0",
-29189 => x"C0C0BFA490F98090",
-29188 => x"C0C0BFA490F98080",
-29187 => x"C0C0BFA490F980F8",
-29186 => x"C0C0BFA490F98082",
-29185 => x"C0C0BFA490F98092",
-29184 => x"C0C0BFA490F98099",
-29183 => x"C0C0BFA490F980B0",
-29182 => x"C0C0BFA490F980A4",
-29181 => x"C0C0BFA490F980F9",
-29180 => x"C0C0BFA490F980C0",
-29179 => x"C0C0BFA490F9F890",
-29178 => x"C0C0BFA490F9F880",
-29177 => x"C0C0BFA490F9F8F8",
-29176 => x"C0C0BFA490F9F882",
-29175 => x"C0C0BFA490F9F892",
-29174 => x"C0C0BFA490F9F899",
-29173 => x"C0C0BFA490F9F8B0",
-29172 => x"C0C0BFA490F9F8A4",
-29171 => x"C0C0BFA490F9F8F9",
-29170 => x"C0C0BFA490F9F8C0",
-29169 => x"C0C0BFA490F98290",
-29168 => x"C0C0BFA490F98280",
-29167 => x"C0C0BFA490F982F8",
-29166 => x"C0C0BFA490F98282",
-29165 => x"C0C0BFA490F98292",
-29164 => x"C0C0BFA490F98299",
-29163 => x"C0C0BFA490F982B0",
-29162 => x"C0C0BFA490F982A4",
-29161 => x"C0C0BFA490F982F9",
-29160 => x"C0C0BFA490F982C0",
-29159 => x"C0C0BFA490F99290",
-29158 => x"C0C0BFA490F99280",
-29157 => x"C0C0BFA490F992F8",
-29156 => x"C0C0BFA490F99282",
-29155 => x"C0C0BFA490F99292",
-29154 => x"C0C0BFA490F99299",
-29153 => x"C0C0BFA490F992B0",
-29152 => x"C0C0BFA490F992A4",
-29151 => x"C0C0BFA490F992F9",
-29150 => x"C0C0BFA490F992C0",
-29149 => x"C0C0BFA490F99990",
-29148 => x"C0C0BFA490F99980",
-29147 => x"C0C0BFA490F999F8",
-29146 => x"C0C0BFA490F99982",
-29145 => x"C0C0BFA490F99992",
-29144 => x"C0C0BFA490F99999",
-29143 => x"C0C0BFA490F999B0",
-29142 => x"C0C0BFA490F999A4",
-29141 => x"C0C0BFA490F999F9",
-29140 => x"C0C0BFA490F999C0",
-29139 => x"C0C0BFA490F9B090",
-29138 => x"C0C0BFA490F9B080",
-29137 => x"C0C0BFA490F9B0F8",
-29136 => x"C0C0BFA490F9B082",
-29135 => x"C0C0BFA490F9B092",
-29134 => x"C0C0BFA490F9B099",
-29133 => x"C0C0BFA490F9B0B0",
-29132 => x"C0C0BFA490F9B0A4",
-29131 => x"C0C0BFA490F9B0F9",
-29130 => x"C0C0BFA490F9B0C0",
-29129 => x"C0C0BFA490F9A490",
-29128 => x"C0C0BFA490F9A480",
-29127 => x"C0C0BFA490F9A4F8",
-29126 => x"C0C0BFA490F9A482",
-29125 => x"C0C0BFA490F9A492",
-29124 => x"C0C0BFA490F9A499",
-29123 => x"C0C0BFA490F9A4B0",
-29122 => x"C0C0BFA490F9A4A4",
-29121 => x"C0C0BFA490F9A4F9",
-29120 => x"C0C0BFA490F9A4C0",
-29119 => x"C0C0BFA490F9F990",
-29118 => x"C0C0BFA490F9F980",
-29117 => x"C0C0BFA490F9F9F8",
-29116 => x"C0C0BFA490F9F982",
-29115 => x"C0C0BFA490F9F992",
-29114 => x"C0C0BFA490F9F999",
-29113 => x"C0C0BFA490F9F9B0",
-29112 => x"C0C0BFA490F9F9A4",
-29111 => x"C0C0BFA490F9F9F9",
-29110 => x"C0C0BFA490F9F9C0",
-29109 => x"C0C0BFA490F9C090",
-29108 => x"C0C0BFA490F9C080",
-29107 => x"C0C0BFA490F9C0F8",
-29106 => x"C0C0BFA490F9C082",
-29105 => x"C0C0BFA490F9C092",
-29104 => x"C0C0BFA490F9C099",
-29103 => x"C0C0BFA490F9C0B0",
-29102 => x"C0C0BFA490F9C0A4",
-29101 => x"C0C0BFA490F9C0F9",
-29100 => x"C0C0BFA490F9C0C0",
-29099 => x"C0C0BFA490C09090",
-29098 => x"C0C0BFA490C09080",
-29097 => x"C0C0BFA490C090F8",
-29096 => x"C0C0BFA490C09082",
-29095 => x"C0C0BFA490C09092",
-29094 => x"C0C0BFA490C09099",
-29093 => x"C0C0BFA490C090B0",
-29092 => x"C0C0BFA490C090A4",
-29091 => x"C0C0BFA490C090F9",
-29090 => x"C0C0BFA490C090C0",
-29089 => x"C0C0BFA490C08090",
-29088 => x"C0C0BFA490C08080",
-29087 => x"C0C0BFA490C080F8",
-29086 => x"C0C0BFA490C08082",
-29085 => x"C0C0BFA490C08092",
-29084 => x"C0C0BFA490C08099",
-29083 => x"C0C0BFA490C080B0",
-29082 => x"C0C0BFA490C080A4",
-29081 => x"C0C0BFA490C080F9",
-29080 => x"C0C0BFA490C080C0",
-29079 => x"C0C0BFA490C0F890",
-29078 => x"C0C0BFA490C0F880",
-29077 => x"C0C0BFA490C0F8F8",
-29076 => x"C0C0BFA490C0F882",
-29075 => x"C0C0BFA490C0F892",
-29074 => x"C0C0BFA490C0F899",
-29073 => x"C0C0BFA490C0F8B0",
-29072 => x"C0C0BFA490C0F8A4",
-29071 => x"C0C0BFA490C0F8F9",
-29070 => x"C0C0BFA490C0F8C0",
-29069 => x"C0C0BFA490C08290",
-29068 => x"C0C0BFA490C08280",
-29067 => x"C0C0BFA490C082F8",
-29066 => x"C0C0BFA490C08282",
-29065 => x"C0C0BFA490C08292",
-29064 => x"C0C0BFA490C08299",
-29063 => x"C0C0BFA490C082B0",
-29062 => x"C0C0BFA490C082A4",
-29061 => x"C0C0BFA490C082F9",
-29060 => x"C0C0BFA490C082C0",
-29059 => x"C0C0BFA490C09290",
-29058 => x"C0C0BFA490C09280",
-29057 => x"C0C0BFA490C092F8",
-29056 => x"C0C0BFA490C09282",
-29055 => x"C0C0BFA490C09292",
-29054 => x"C0C0BFA490C09299",
-29053 => x"C0C0BFA490C092B0",
-29052 => x"C0C0BFA490C092A4",
-29051 => x"C0C0BFA490C092F9",
-29050 => x"C0C0BFA490C092C0",
-29049 => x"C0C0BFA490C09990",
-29048 => x"C0C0BFA490C09980",
-29047 => x"C0C0BFA490C099F8",
-29046 => x"C0C0BFA490C09982",
-29045 => x"C0C0BFA490C09992",
-29044 => x"C0C0BFA490C09999",
-29043 => x"C0C0BFA490C099B0",
-29042 => x"C0C0BFA490C099A4",
-29041 => x"C0C0BFA490C099F9",
-29040 => x"C0C0BFA490C099C0",
-29039 => x"C0C0BFA490C0B090",
-29038 => x"C0C0BFA490C0B080",
-29037 => x"C0C0BFA490C0B0F8",
-29036 => x"C0C0BFA490C0B082",
-29035 => x"C0C0BFA490C0B092",
-29034 => x"C0C0BFA490C0B099",
-29033 => x"C0C0BFA490C0B0B0",
-29032 => x"C0C0BFA490C0B0A4",
-29031 => x"C0C0BFA490C0B0F9",
-29030 => x"C0C0BFA490C0B0C0",
-29029 => x"C0C0BFA490C0A490",
-29028 => x"C0C0BFA490C0A480",
-29027 => x"C0C0BFA490C0A4F8",
-29026 => x"C0C0BFA490C0A482",
-29025 => x"C0C0BFA490C0A492",
-29024 => x"C0C0BFA490C0A499",
-29023 => x"C0C0BFA490C0A4B0",
-29022 => x"C0C0BFA490C0A4A4",
-29021 => x"C0C0BFA490C0A4F9",
-29020 => x"C0C0BFA490C0A4C0",
-29019 => x"C0C0BFA490C0F990",
-29018 => x"C0C0BFA490C0F980",
-29017 => x"C0C0BFA490C0F9F8",
-29016 => x"C0C0BFA490C0F982",
-29015 => x"C0C0BFA490C0F992",
-29014 => x"C0C0BFA490C0F999",
-29013 => x"C0C0BFA490C0F9B0",
-29012 => x"C0C0BFA490C0F9A4",
-29011 => x"C0C0BFA490C0F9F9",
-29010 => x"C0C0BFA490C0F9C0",
-29009 => x"C0C0BFA490C0C090",
-29008 => x"C0C0BFA490C0C080",
-29007 => x"C0C0BFA490C0C0F8",
-29006 => x"C0C0BFA490C0C082",
-29005 => x"C0C0BFA490C0C092",
-29004 => x"C0C0BFA490C0C099",
-29003 => x"C0C0BFA490C0C0B0",
-29002 => x"C0C0BFA490C0C0A4",
-29001 => x"C0C0BFA490C0C0F9",
-29000 => x"C0C0BFA490C0C0C0",
-28999 => x"C0C0BFA480909090",
-28998 => x"C0C0BFA480909080",
-28997 => x"C0C0BFA4809090F8",
-28996 => x"C0C0BFA480909082",
-28995 => x"C0C0BFA480909092",
-28994 => x"C0C0BFA480909099",
-28993 => x"C0C0BFA4809090B0",
-28992 => x"C0C0BFA4809090A4",
-28991 => x"C0C0BFA4809090F9",
-28990 => x"C0C0BFA4809090C0",
-28989 => x"C0C0BFA480908090",
-28988 => x"C0C0BFA480908080",
-28987 => x"C0C0BFA4809080F8",
-28986 => x"C0C0BFA480908082",
-28985 => x"C0C0BFA480908092",
-28984 => x"C0C0BFA480908099",
-28983 => x"C0C0BFA4809080B0",
-28982 => x"C0C0BFA4809080A4",
-28981 => x"C0C0BFA4809080F9",
-28980 => x"C0C0BFA4809080C0",
-28979 => x"C0C0BFA48090F890",
-28978 => x"C0C0BFA48090F880",
-28977 => x"C0C0BFA48090F8F8",
-28976 => x"C0C0BFA48090F882",
-28975 => x"C0C0BFA48090F892",
-28974 => x"C0C0BFA48090F899",
-28973 => x"C0C0BFA48090F8B0",
-28972 => x"C0C0BFA48090F8A4",
-28971 => x"C0C0BFA48090F8F9",
-28970 => x"C0C0BFA48090F8C0",
-28969 => x"C0C0BFA480908290",
-28968 => x"C0C0BFA480908280",
-28967 => x"C0C0BFA4809082F8",
-28966 => x"C0C0BFA480908282",
-28965 => x"C0C0BFA480908292",
-28964 => x"C0C0BFA480908299",
-28963 => x"C0C0BFA4809082B0",
-28962 => x"C0C0BFA4809082A4",
-28961 => x"C0C0BFA4809082F9",
-28960 => x"C0C0BFA4809082C0",
-28959 => x"C0C0BFA480909290",
-28958 => x"C0C0BFA480909280",
-28957 => x"C0C0BFA4809092F8",
-28956 => x"C0C0BFA480909282",
-28955 => x"C0C0BFA480909292",
-28954 => x"C0C0BFA480909299",
-28953 => x"C0C0BFA4809092B0",
-28952 => x"C0C0BFA4809092A4",
-28951 => x"C0C0BFA4809092F9",
-28950 => x"C0C0BFA4809092C0",
-28949 => x"C0C0BFA480909990",
-28948 => x"C0C0BFA480909980",
-28947 => x"C0C0BFA4809099F8",
-28946 => x"C0C0BFA480909982",
-28945 => x"C0C0BFA480909992",
-28944 => x"C0C0BFA480909999",
-28943 => x"C0C0BFA4809099B0",
-28942 => x"C0C0BFA4809099A4",
-28941 => x"C0C0BFA4809099F9",
-28940 => x"C0C0BFA4809099C0",
-28939 => x"C0C0BFA48090B090",
-28938 => x"C0C0BFA48090B080",
-28937 => x"C0C0BFA48090B0F8",
-28936 => x"C0C0BFA48090B082",
-28935 => x"C0C0BFA48090B092",
-28934 => x"C0C0BFA48090B099",
-28933 => x"C0C0BFA48090B0B0",
-28932 => x"C0C0BFA48090B0A4",
-28931 => x"C0C0BFA48090B0F9",
-28930 => x"C0C0BFA48090B0C0",
-28929 => x"C0C0BFA48090A490",
-28928 => x"C0C0BFA48090A480",
-28927 => x"C0C0BFA48090A4F8",
-28926 => x"C0C0BFA48090A482",
-28925 => x"C0C0BFA48090A492",
-28924 => x"C0C0BFA48090A499",
-28923 => x"C0C0BFA48090A4B0",
-28922 => x"C0C0BFA48090A4A4",
-28921 => x"C0C0BFA48090A4F9",
-28920 => x"C0C0BFA48090A4C0",
-28919 => x"C0C0BFA48090F990",
-28918 => x"C0C0BFA48090F980",
-28917 => x"C0C0BFA48090F9F8",
-28916 => x"C0C0BFA48090F982",
-28915 => x"C0C0BFA48090F992",
-28914 => x"C0C0BFA48090F999",
-28913 => x"C0C0BFA48090F9B0",
-28912 => x"C0C0BFA48090F9A4",
-28911 => x"C0C0BFA48090F9F9",
-28910 => x"C0C0BFA48090F9C0",
-28909 => x"C0C0BFA48090C090",
-28908 => x"C0C0BFA48090C080",
-28907 => x"C0C0BFA48090C0F8",
-28906 => x"C0C0BFA48090C082",
-28905 => x"C0C0BFA48090C092",
-28904 => x"C0C0BFA48090C099",
-28903 => x"C0C0BFA48090C0B0",
-28902 => x"C0C0BFA48090C0A4",
-28901 => x"C0C0BFA48090C0F9",
-28900 => x"C0C0BFA48090C0C0",
-28899 => x"C0C0BFA480809090",
-28898 => x"C0C0BFA480809080",
-28897 => x"C0C0BFA4808090F8",
-28896 => x"C0C0BFA480809082",
-28895 => x"C0C0BFA480809092",
-28894 => x"C0C0BFA480809099",
-28893 => x"C0C0BFA4808090B0",
-28892 => x"C0C0BFA4808090A4",
-28891 => x"C0C0BFA4808090F9",
-28890 => x"C0C0BFA4808090C0",
-28889 => x"C0C0BFA480808090",
-28888 => x"C0C0BFA480808080",
-28887 => x"C0C0BFA4808080F8",
-28886 => x"C0C0BFA480808082",
-28885 => x"C0C0BFA480808092",
-28884 => x"C0C0BFA480808099",
-28883 => x"C0C0BFA4808080B0",
-28882 => x"C0C0BFA4808080A4",
-28881 => x"C0C0BFA4808080F9",
-28880 => x"C0C0BFA4808080C0",
-28879 => x"C0C0BFA48080F890",
-28878 => x"C0C0BFA48080F880",
-28877 => x"C0C0BFA48080F8F8",
-28876 => x"C0C0BFA48080F882",
-28875 => x"C0C0BFA48080F892",
-28874 => x"C0C0BFA48080F899",
-28873 => x"C0C0BFA48080F8B0",
-28872 => x"C0C0BFA48080F8A4",
-28871 => x"C0C0BFA48080F8F9",
-28870 => x"C0C0BFA48080F8C0",
-28869 => x"C0C0BFA480808290",
-28868 => x"C0C0BFA480808280",
-28867 => x"C0C0BFA4808082F8",
-28866 => x"C0C0BFA480808282",
-28865 => x"C0C0BFA480808292",
-28864 => x"C0C0BFA480808299",
-28863 => x"C0C0BFA4808082B0",
-28862 => x"C0C0BFA4808082A4",
-28861 => x"C0C0BFA4808082F9",
-28860 => x"C0C0BFA4808082C0",
-28859 => x"C0C0BFA480809290",
-28858 => x"C0C0BFA480809280",
-28857 => x"C0C0BFA4808092F8",
-28856 => x"C0C0BFA480809282",
-28855 => x"C0C0BFA480809292",
-28854 => x"C0C0BFA480809299",
-28853 => x"C0C0BFA4808092B0",
-28852 => x"C0C0BFA4808092A4",
-28851 => x"C0C0BFA4808092F9",
-28850 => x"C0C0BFA4808092C0",
-28849 => x"C0C0BFA480809990",
-28848 => x"C0C0BFA480809980",
-28847 => x"C0C0BFA4808099F8",
-28846 => x"C0C0BFA480809982",
-28845 => x"C0C0BFA480809992",
-28844 => x"C0C0BFA480809999",
-28843 => x"C0C0BFA4808099B0",
-28842 => x"C0C0BFA4808099A4",
-28841 => x"C0C0BFA4808099F9",
-28840 => x"C0C0BFA4808099C0",
-28839 => x"C0C0BFA48080B090",
-28838 => x"C0C0BFA48080B080",
-28837 => x"C0C0BFA48080B0F8",
-28836 => x"C0C0BFA48080B082",
-28835 => x"C0C0BFA48080B092",
-28834 => x"C0C0BFA48080B099",
-28833 => x"C0C0BFA48080B0B0",
-28832 => x"C0C0BFA48080B0A4",
-28831 => x"C0C0BFA48080B0F9",
-28830 => x"C0C0BFA48080B0C0",
-28829 => x"C0C0BFA48080A490",
-28828 => x"C0C0BFA48080A480",
-28827 => x"C0C0BFA48080A4F8",
-28826 => x"C0C0BFA48080A482",
-28825 => x"C0C0BFA48080A492",
-28824 => x"C0C0BFA48080A499",
-28823 => x"C0C0BFA48080A4B0",
-28822 => x"C0C0BFA48080A4A4",
-28821 => x"C0C0BFA48080A4F9",
-28820 => x"C0C0BFA48080A4C0",
-28819 => x"C0C0BFA48080F990",
-28818 => x"C0C0BFA48080F980",
-28817 => x"C0C0BFA48080F9F8",
-28816 => x"C0C0BFA48080F982",
-28815 => x"C0C0BFA48080F992",
-28814 => x"C0C0BFA48080F999",
-28813 => x"C0C0BFA48080F9B0",
-28812 => x"C0C0BFA48080F9A4",
-28811 => x"C0C0BFA48080F9F9",
-28810 => x"C0C0BFA48080F9C0",
-28809 => x"C0C0BFA48080C090",
-28808 => x"C0C0BFA48080C080",
-28807 => x"C0C0BFA48080C0F8",
-28806 => x"C0C0BFA48080C082",
-28805 => x"C0C0BFA48080C092",
-28804 => x"C0C0BFA48080C099",
-28803 => x"C0C0BFA48080C0B0",
-28802 => x"C0C0BFA48080C0A4",
-28801 => x"C0C0BFA48080C0F9",
-28800 => x"C0C0BFA48080C0C0",
-28799 => x"C0C0BFA480F89090",
-28798 => x"C0C0BFA480F89080",
-28797 => x"C0C0BFA480F890F8",
-28796 => x"C0C0BFA480F89082",
-28795 => x"C0C0BFA480F89092",
-28794 => x"C0C0BFA480F89099",
-28793 => x"C0C0BFA480F890B0",
-28792 => x"C0C0BFA480F890A4",
-28791 => x"C0C0BFA480F890F9",
-28790 => x"C0C0BFA480F890C0",
-28789 => x"C0C0BFA480F88090",
-28788 => x"C0C0BFA480F88080",
-28787 => x"C0C0BFA480F880F8",
-28786 => x"C0C0BFA480F88082",
-28785 => x"C0C0BFA480F88092",
-28784 => x"C0C0BFA480F88099",
-28783 => x"C0C0BFA480F880B0",
-28782 => x"C0C0BFA480F880A4",
-28781 => x"C0C0BFA480F880F9",
-28780 => x"C0C0BFA480F880C0",
-28779 => x"C0C0BFA480F8F890",
-28778 => x"C0C0BFA480F8F880",
-28777 => x"C0C0BFA480F8F8F8",
-28776 => x"C0C0BFA480F8F882",
-28775 => x"C0C0BFA480F8F892",
-28774 => x"C0C0BFA480F8F899",
-28773 => x"C0C0BFA480F8F8B0",
-28772 => x"C0C0BFA480F8F8A4",
-28771 => x"C0C0BFA480F8F8F9",
-28770 => x"C0C0BFA480F8F8C0",
-28769 => x"C0C0BFA480F88290",
-28768 => x"C0C0BFA480F88280",
-28767 => x"C0C0BFA480F882F8",
-28766 => x"C0C0BFA480F88282",
-28765 => x"C0C0BFA480F88292",
-28764 => x"C0C0BFA480F88299",
-28763 => x"C0C0BFA480F882B0",
-28762 => x"C0C0BFA480F882A4",
-28761 => x"C0C0BFA480F882F9",
-28760 => x"C0C0BFA480F882C0",
-28759 => x"C0C0BFA480F89290",
-28758 => x"C0C0BFA480F89280",
-28757 => x"C0C0BFA480F892F8",
-28756 => x"C0C0BFA480F89282",
-28755 => x"C0C0BFA480F89292",
-28754 => x"C0C0BFA480F89299",
-28753 => x"C0C0BFA480F892B0",
-28752 => x"C0C0BFA480F892A4",
-28751 => x"C0C0BFA480F892F9",
-28750 => x"C0C0BFA480F892C0",
-28749 => x"C0C0BFA480F89990",
-28748 => x"C0C0BFA480F89980",
-28747 => x"C0C0BFA480F899F8",
-28746 => x"C0C0BFA480F89982",
-28745 => x"C0C0BFA480F89992",
-28744 => x"C0C0BFA480F89999",
-28743 => x"C0C0BFA480F899B0",
-28742 => x"C0C0BFA480F899A4",
-28741 => x"C0C0BFA480F899F9",
-28740 => x"C0C0BFA480F899C0",
-28739 => x"C0C0BFA480F8B090",
-28738 => x"C0C0BFA480F8B080",
-28737 => x"C0C0BFA480F8B0F8",
-28736 => x"C0C0BFA480F8B082",
-28735 => x"C0C0BFA480F8B092",
-28734 => x"C0C0BFA480F8B099",
-28733 => x"C0C0BFA480F8B0B0",
-28732 => x"C0C0BFA480F8B0A4",
-28731 => x"C0C0BFA480F8B0F9",
-28730 => x"C0C0BFA480F8B0C0",
-28729 => x"C0C0BFA480F8A490",
-28728 => x"C0C0BFA480F8A480",
-28727 => x"C0C0BFA480F8A4F8",
-28726 => x"C0C0BFA480F8A482",
-28725 => x"C0C0BFA480F8A492",
-28724 => x"C0C0BFA480F8A499",
-28723 => x"C0C0BFA480F8A4B0",
-28722 => x"C0C0BFA480F8A4A4",
-28721 => x"C0C0BFA480F8A4F9",
-28720 => x"C0C0BFA480F8A4C0",
-28719 => x"C0C0BFA480F8F990",
-28718 => x"C0C0BFA480F8F980",
-28717 => x"C0C0BFA480F8F9F8",
-28716 => x"C0C0BFA480F8F982",
-28715 => x"C0C0BFA480F8F992",
-28714 => x"C0C0BFA480F8F999",
-28713 => x"C0C0BFA480F8F9B0",
-28712 => x"C0C0BFA480F8F9A4",
-28711 => x"C0C0BFA480F8F9F9",
-28710 => x"C0C0BFA480F8F9C0",
-28709 => x"C0C0BFA480F8C090",
-28708 => x"C0C0BFA480F8C080",
-28707 => x"C0C0BFA480F8C0F8",
-28706 => x"C0C0BFA480F8C082",
-28705 => x"C0C0BFA480F8C092",
-28704 => x"C0C0BFA480F8C099",
-28703 => x"C0C0BFA480F8C0B0",
-28702 => x"C0C0BFA480F8C0A4",
-28701 => x"C0C0BFA480F8C0F9",
-28700 => x"C0C0BFA480F8C0C0",
-28699 => x"C0C0BFA480829090",
-28698 => x"C0C0BFA480829080",
-28697 => x"C0C0BFA4808290F8",
-28696 => x"C0C0BFA480829082",
-28695 => x"C0C0BFA480829092",
-28694 => x"C0C0BFA480829099",
-28693 => x"C0C0BFA4808290B0",
-28692 => x"C0C0BFA4808290A4",
-28691 => x"C0C0BFA4808290F9",
-28690 => x"C0C0BFA4808290C0",
-28689 => x"C0C0BFA480828090",
-28688 => x"C0C0BFA480828080",
-28687 => x"C0C0BFA4808280F8",
-28686 => x"C0C0BFA480828082",
-28685 => x"C0C0BFA480828092",
-28684 => x"C0C0BFA480828099",
-28683 => x"C0C0BFA4808280B0",
-28682 => x"C0C0BFA4808280A4",
-28681 => x"C0C0BFA4808280F9",
-28680 => x"C0C0BFA4808280C0",
-28679 => x"C0C0BFA48082F890",
-28678 => x"C0C0BFA48082F880",
-28677 => x"C0C0BFA48082F8F8",
-28676 => x"C0C0BFA48082F882",
-28675 => x"C0C0BFA48082F892",
-28674 => x"C0C0BFA48082F899",
-28673 => x"C0C0BFA48082F8B0",
-28672 => x"C0C0BFA48082F8A4",
-28671 => x"C0C0BFA48082F8F9",
-28670 => x"C0C0BFA48082F8C0",
-28669 => x"C0C0BFA480828290",
-28668 => x"C0C0BFA480828280",
-28667 => x"C0C0BFA4808282F8",
-28666 => x"C0C0BFA480828282",
-28665 => x"C0C0BFA480828292",
-28664 => x"C0C0BFA480828299",
-28663 => x"C0C0BFA4808282B0",
-28662 => x"C0C0BFA4808282A4",
-28661 => x"C0C0BFA4808282F9",
-28660 => x"C0C0BFA4808282C0",
-28659 => x"C0C0BFA480829290",
-28658 => x"C0C0BFA480829280",
-28657 => x"C0C0BFA4808292F8",
-28656 => x"C0C0BFA480829282",
-28655 => x"C0C0BFA480829292",
-28654 => x"C0C0BFA480829299",
-28653 => x"C0C0BFA4808292B0",
-28652 => x"C0C0BFA4808292A4",
-28651 => x"C0C0BFA4808292F9",
-28650 => x"C0C0BFA4808292C0",
-28649 => x"C0C0BFA480829990",
-28648 => x"C0C0BFA480829980",
-28647 => x"C0C0BFA4808299F8",
-28646 => x"C0C0BFA480829982",
-28645 => x"C0C0BFA480829992",
-28644 => x"C0C0BFA480829999",
-28643 => x"C0C0BFA4808299B0",
-28642 => x"C0C0BFA4808299A4",
-28641 => x"C0C0BFA4808299F9",
-28640 => x"C0C0BFA4808299C0",
-28639 => x"C0C0BFA48082B090",
-28638 => x"C0C0BFA48082B080",
-28637 => x"C0C0BFA48082B0F8",
-28636 => x"C0C0BFA48082B082",
-28635 => x"C0C0BFA48082B092",
-28634 => x"C0C0BFA48082B099",
-28633 => x"C0C0BFA48082B0B0",
-28632 => x"C0C0BFA48082B0A4",
-28631 => x"C0C0BFA48082B0F9",
-28630 => x"C0C0BFA48082B0C0",
-28629 => x"C0C0BFA48082A490",
-28628 => x"C0C0BFA48082A480",
-28627 => x"C0C0BFA48082A4F8",
-28626 => x"C0C0BFA48082A482",
-28625 => x"C0C0BFA48082A492",
-28624 => x"C0C0BFA48082A499",
-28623 => x"C0C0BFA48082A4B0",
-28622 => x"C0C0BFA48082A4A4",
-28621 => x"C0C0BFA48082A4F9",
-28620 => x"C0C0BFA48082A4C0",
-28619 => x"C0C0BFA48082F990",
-28618 => x"C0C0BFA48082F980",
-28617 => x"C0C0BFA48082F9F8",
-28616 => x"C0C0BFA48082F982",
-28615 => x"C0C0BFA48082F992",
-28614 => x"C0C0BFA48082F999",
-28613 => x"C0C0BFA48082F9B0",
-28612 => x"C0C0BFA48082F9A4",
-28611 => x"C0C0BFA48082F9F9",
-28610 => x"C0C0BFA48082F9C0",
-28609 => x"C0C0BFA48082C090",
-28608 => x"C0C0BFA48082C080",
-28607 => x"C0C0BFA48082C0F8",
-28606 => x"C0C0BFA48082C082",
-28605 => x"C0C0BFA48082C092",
-28604 => x"C0C0BFA48082C099",
-28603 => x"C0C0BFA48082C0B0",
-28602 => x"C0C0BFA48082C0A4",
-28601 => x"C0C0BFA48082C0F9",
-28600 => x"C0C0BFA48082C0C0",
-28599 => x"C0C0BFA480929090",
-28598 => x"C0C0BFA480929080",
-28597 => x"C0C0BFA4809290F8",
-28596 => x"C0C0BFA480929082",
-28595 => x"C0C0BFA480929092",
-28594 => x"C0C0BFA480929099",
-28593 => x"C0C0BFA4809290B0",
-28592 => x"C0C0BFA4809290A4",
-28591 => x"C0C0BFA4809290F9",
-28590 => x"C0C0BFA4809290C0",
-28589 => x"C0C0BFA480928090",
-28588 => x"C0C0BFA480928080",
-28587 => x"C0C0BFA4809280F8",
-28586 => x"C0C0BFA480928082",
-28585 => x"C0C0BFA480928092",
-28584 => x"C0C0BFA480928099",
-28583 => x"C0C0BFA4809280B0",
-28582 => x"C0C0BFA4809280A4",
-28581 => x"C0C0BFA4809280F9",
-28580 => x"C0C0BFA4809280C0",
-28579 => x"C0C0BFA48092F890",
-28578 => x"C0C0BFA48092F880",
-28577 => x"C0C0BFA48092F8F8",
-28576 => x"C0C0BFA48092F882",
-28575 => x"C0C0BFA48092F892",
-28574 => x"C0C0BFA48092F899",
-28573 => x"C0C0BFA48092F8B0",
-28572 => x"C0C0BFA48092F8A4",
-28571 => x"C0C0BFA48092F8F9",
-28570 => x"C0C0BFA48092F8C0",
-28569 => x"C0C0BFA480928290",
-28568 => x"C0C0BFA480928280",
-28567 => x"C0C0BFA4809282F8",
-28566 => x"C0C0BFA480928282",
-28565 => x"C0C0BFA480928292",
-28564 => x"C0C0BFA480928299",
-28563 => x"C0C0BFA4809282B0",
-28562 => x"C0C0BFA4809282A4",
-28561 => x"C0C0BFA4809282F9",
-28560 => x"C0C0BFA4809282C0",
-28559 => x"C0C0BFA480929290",
-28558 => x"C0C0BFA480929280",
-28557 => x"C0C0BFA4809292F8",
-28556 => x"C0C0BFA480929282",
-28555 => x"C0C0BFA480929292",
-28554 => x"C0C0BFA480929299",
-28553 => x"C0C0BFA4809292B0",
-28552 => x"C0C0BFA4809292A4",
-28551 => x"C0C0BFA4809292F9",
-28550 => x"C0C0BFA4809292C0",
-28549 => x"C0C0BFA480929990",
-28548 => x"C0C0BFA480929980",
-28547 => x"C0C0BFA4809299F8",
-28546 => x"C0C0BFA480929982",
-28545 => x"C0C0BFA480929992",
-28544 => x"C0C0BFA480929999",
-28543 => x"C0C0BFA4809299B0",
-28542 => x"C0C0BFA4809299A4",
-28541 => x"C0C0BFA4809299F9",
-28540 => x"C0C0BFA4809299C0",
-28539 => x"C0C0BFA48092B090",
-28538 => x"C0C0BFA48092B080",
-28537 => x"C0C0BFA48092B0F8",
-28536 => x"C0C0BFA48092B082",
-28535 => x"C0C0BFA48092B092",
-28534 => x"C0C0BFA48092B099",
-28533 => x"C0C0BFA48092B0B0",
-28532 => x"C0C0BFA48092B0A4",
-28531 => x"C0C0BFA48092B0F9",
-28530 => x"C0C0BFA48092B0C0",
-28529 => x"C0C0BFA48092A490",
-28528 => x"C0C0BFA48092A480",
-28527 => x"C0C0BFA48092A4F8",
-28526 => x"C0C0BFA48092A482",
-28525 => x"C0C0BFA48092A492",
-28524 => x"C0C0BFA48092A499",
-28523 => x"C0C0BFA48092A4B0",
-28522 => x"C0C0BFA48092A4A4",
-28521 => x"C0C0BFA48092A4F9",
-28520 => x"C0C0BFA48092A4C0",
-28519 => x"C0C0BFA48092F990",
-28518 => x"C0C0BFA48092F980",
-28517 => x"C0C0BFA48092F9F8",
-28516 => x"C0C0BFA48092F982",
-28515 => x"C0C0BFA48092F992",
-28514 => x"C0C0BFA48092F999",
-28513 => x"C0C0BFA48092F9B0",
-28512 => x"C0C0BFA48092F9A4",
-28511 => x"C0C0BFA48092F9F9",
-28510 => x"C0C0BFA48092F9C0",
-28509 => x"C0C0BFA48092C090",
-28508 => x"C0C0BFA48092C080",
-28507 => x"C0C0BFA48092C0F8",
-28506 => x"C0C0BFA48092C082",
-28505 => x"C0C0BFA48092C092",
-28504 => x"C0C0BFA48092C099",
-28503 => x"C0C0BFA48092C0B0",
-28502 => x"C0C0BFA48092C0A4",
-28501 => x"C0C0BFA48092C0F9",
-28500 => x"C0C0BFA48092C0C0",
-28499 => x"C0C0BFA480999090",
-28498 => x"C0C0BFA480999080",
-28497 => x"C0C0BFA4809990F8",
-28496 => x"C0C0BFA480999082",
-28495 => x"C0C0BFA480999092",
-28494 => x"C0C0BFA480999099",
-28493 => x"C0C0BFA4809990B0",
-28492 => x"C0C0BFA4809990A4",
-28491 => x"C0C0BFA4809990F9",
-28490 => x"C0C0BFA4809990C0",
-28489 => x"C0C0BFA480998090",
-28488 => x"C0C0BFA480998080",
-28487 => x"C0C0BFA4809980F8",
-28486 => x"C0C0BFA480998082",
-28485 => x"C0C0BFA480998092",
-28484 => x"C0C0BFA480998099",
-28483 => x"C0C0BFA4809980B0",
-28482 => x"C0C0BFA4809980A4",
-28481 => x"C0C0BFA4809980F9",
-28480 => x"C0C0BFA4809980C0",
-28479 => x"C0C0BFA48099F890",
-28478 => x"C0C0BFA48099F880",
-28477 => x"C0C0BFA48099F8F8",
-28476 => x"C0C0BFA48099F882",
-28475 => x"C0C0BFA48099F892",
-28474 => x"C0C0BFA48099F899",
-28473 => x"C0C0BFA48099F8B0",
-28472 => x"C0C0BFA48099F8A4",
-28471 => x"C0C0BFA48099F8F9",
-28470 => x"C0C0BFA48099F8C0",
-28469 => x"C0C0BFA480998290",
-28468 => x"C0C0BFA480998280",
-28467 => x"C0C0BFA4809982F8",
-28466 => x"C0C0BFA480998282",
-28465 => x"C0C0BFA480998292",
-28464 => x"C0C0BFA480998299",
-28463 => x"C0C0BFA4809982B0",
-28462 => x"C0C0BFA4809982A4",
-28461 => x"C0C0BFA4809982F9",
-28460 => x"C0C0BFA4809982C0",
-28459 => x"C0C0BFA480999290",
-28458 => x"C0C0BFA480999280",
-28457 => x"C0C0BFA4809992F8",
-28456 => x"C0C0BFA480999282",
-28455 => x"C0C0BFA480999292",
-28454 => x"C0C0BFA480999299",
-28453 => x"C0C0BFA4809992B0",
-28452 => x"C0C0BFA4809992A4",
-28451 => x"C0C0BFA4809992F9",
-28450 => x"C0C0BFA4809992C0",
-28449 => x"C0C0BFA480999990",
-28448 => x"C0C0BFA480999980",
-28447 => x"C0C0BFA4809999F8",
-28446 => x"C0C0BFA480999982",
-28445 => x"C0C0BFA480999992",
-28444 => x"C0C0BFA480999999",
-28443 => x"C0C0BFA4809999B0",
-28442 => x"C0C0BFA4809999A4",
-28441 => x"C0C0BFA4809999F9",
-28440 => x"C0C0BFA4809999C0",
-28439 => x"C0C0BFA48099B090",
-28438 => x"C0C0BFA48099B080",
-28437 => x"C0C0BFA48099B0F8",
-28436 => x"C0C0BFA48099B082",
-28435 => x"C0C0BFA48099B092",
-28434 => x"C0C0BFA48099B099",
-28433 => x"C0C0BFA48099B0B0",
-28432 => x"C0C0BFA48099B0A4",
-28431 => x"C0C0BFA48099B0F9",
-28430 => x"C0C0BFA48099B0C0",
-28429 => x"C0C0BFA48099A490",
-28428 => x"C0C0BFA48099A480",
-28427 => x"C0C0BFA48099A4F8",
-28426 => x"C0C0BFA48099A482",
-28425 => x"C0C0BFA48099A492",
-28424 => x"C0C0BFA48099A499",
-28423 => x"C0C0BFA48099A4B0",
-28422 => x"C0C0BFA48099A4A4",
-28421 => x"C0C0BFA48099A4F9",
-28420 => x"C0C0BFA48099A4C0",
-28419 => x"C0C0BFA48099F990",
-28418 => x"C0C0BFA48099F980",
-28417 => x"C0C0BFA48099F9F8",
-28416 => x"C0C0BFA48099F982",
-28415 => x"C0C0BFA48099F992",
-28414 => x"C0C0BFA48099F999",
-28413 => x"C0C0BFA48099F9B0",
-28412 => x"C0C0BFA48099F9A4",
-28411 => x"C0C0BFA48099F9F9",
-28410 => x"C0C0BFA48099F9C0",
-28409 => x"C0C0BFA48099C090",
-28408 => x"C0C0BFA48099C080",
-28407 => x"C0C0BFA48099C0F8",
-28406 => x"C0C0BFA48099C082",
-28405 => x"C0C0BFA48099C092",
-28404 => x"C0C0BFA48099C099",
-28403 => x"C0C0BFA48099C0B0",
-28402 => x"C0C0BFA48099C0A4",
-28401 => x"C0C0BFA48099C0F9",
-28400 => x"C0C0BFA48099C0C0",
-28399 => x"C0C0BFA480B09090",
-28398 => x"C0C0BFA480B09080",
-28397 => x"C0C0BFA480B090F8",
-28396 => x"C0C0BFA480B09082",
-28395 => x"C0C0BFA480B09092",
-28394 => x"C0C0BFA480B09099",
-28393 => x"C0C0BFA480B090B0",
-28392 => x"C0C0BFA480B090A4",
-28391 => x"C0C0BFA480B090F9",
-28390 => x"C0C0BFA480B090C0",
-28389 => x"C0C0BFA480B08090",
-28388 => x"C0C0BFA480B08080",
-28387 => x"C0C0BFA480B080F8",
-28386 => x"C0C0BFA480B08082",
-28385 => x"C0C0BFA480B08092",
-28384 => x"C0C0BFA480B08099",
-28383 => x"C0C0BFA480B080B0",
-28382 => x"C0C0BFA480B080A4",
-28381 => x"C0C0BFA480B080F9",
-28380 => x"C0C0BFA480B080C0",
-28379 => x"C0C0BFA480B0F890",
-28378 => x"C0C0BFA480B0F880",
-28377 => x"C0C0BFA480B0F8F8",
-28376 => x"C0C0BFA480B0F882",
-28375 => x"C0C0BFA480B0F892",
-28374 => x"C0C0BFA480B0F899",
-28373 => x"C0C0BFA480B0F8B0",
-28372 => x"C0C0BFA480B0F8A4",
-28371 => x"C0C0BFA480B0F8F9",
-28370 => x"C0C0BFA480B0F8C0",
-28369 => x"C0C0BFA480B08290",
-28368 => x"C0C0BFA480B08280",
-28367 => x"C0C0BFA480B082F8",
-28366 => x"C0C0BFA480B08282",
-28365 => x"C0C0BFA480B08292",
-28364 => x"C0C0BFA480B08299",
-28363 => x"C0C0BFA480B082B0",
-28362 => x"C0C0BFA480B082A4",
-28361 => x"C0C0BFA480B082F9",
-28360 => x"C0C0BFA480B082C0",
-28359 => x"C0C0BFA480B09290",
-28358 => x"C0C0BFA480B09280",
-28357 => x"C0C0BFA480B092F8",
-28356 => x"C0C0BFA480B09282",
-28355 => x"C0C0BFA480B09292",
-28354 => x"C0C0BFA480B09299",
-28353 => x"C0C0BFA480B092B0",
-28352 => x"C0C0BFA480B092A4",
-28351 => x"C0C0BFA480B092F9",
-28350 => x"C0C0BFA480B092C0",
-28349 => x"C0C0BFA480B09990",
-28348 => x"C0C0BFA480B09980",
-28347 => x"C0C0BFA480B099F8",
-28346 => x"C0C0BFA480B09982",
-28345 => x"C0C0BFA480B09992",
-28344 => x"C0C0BFA480B09999",
-28343 => x"C0C0BFA480B099B0",
-28342 => x"C0C0BFA480B099A4",
-28341 => x"C0C0BFA480B099F9",
-28340 => x"C0C0BFA480B099C0",
-28339 => x"C0C0BFA480B0B090",
-28338 => x"C0C0BFA480B0B080",
-28337 => x"C0C0BFA480B0B0F8",
-28336 => x"C0C0BFA480B0B082",
-28335 => x"C0C0BFA480B0B092",
-28334 => x"C0C0BFA480B0B099",
-28333 => x"C0C0BFA480B0B0B0",
-28332 => x"C0C0BFA480B0B0A4",
-28331 => x"C0C0BFA480B0B0F9",
-28330 => x"C0C0BFA480B0B0C0",
-28329 => x"C0C0BFA480B0A490",
-28328 => x"C0C0BFA480B0A480",
-28327 => x"C0C0BFA480B0A4F8",
-28326 => x"C0C0BFA480B0A482",
-28325 => x"C0C0BFA480B0A492",
-28324 => x"C0C0BFA480B0A499",
-28323 => x"C0C0BFA480B0A4B0",
-28322 => x"C0C0BFA480B0A4A4",
-28321 => x"C0C0BFA480B0A4F9",
-28320 => x"C0C0BFA480B0A4C0",
-28319 => x"C0C0BFA480B0F990",
-28318 => x"C0C0BFA480B0F980",
-28317 => x"C0C0BFA480B0F9F8",
-28316 => x"C0C0BFA480B0F982",
-28315 => x"C0C0BFA480B0F992",
-28314 => x"C0C0BFA480B0F999",
-28313 => x"C0C0BFA480B0F9B0",
-28312 => x"C0C0BFA480B0F9A4",
-28311 => x"C0C0BFA480B0F9F9",
-28310 => x"C0C0BFA480B0F9C0",
-28309 => x"C0C0BFA480B0C090",
-28308 => x"C0C0BFA480B0C080",
-28307 => x"C0C0BFA480B0C0F8",
-28306 => x"C0C0BFA480B0C082",
-28305 => x"C0C0BFA480B0C092",
-28304 => x"C0C0BFA480B0C099",
-28303 => x"C0C0BFA480B0C0B0",
-28302 => x"C0C0BFA480B0C0A4",
-28301 => x"C0C0BFA480B0C0F9",
-28300 => x"C0C0BFA480B0C0C0",
-28299 => x"C0C0BFA480A49090",
-28298 => x"C0C0BFA480A49080",
-28297 => x"C0C0BFA480A490F8",
-28296 => x"C0C0BFA480A49082",
-28295 => x"C0C0BFA480A49092",
-28294 => x"C0C0BFA480A49099",
-28293 => x"C0C0BFA480A490B0",
-28292 => x"C0C0BFA480A490A4",
-28291 => x"C0C0BFA480A490F9",
-28290 => x"C0C0BFA480A490C0",
-28289 => x"C0C0BFA480A48090",
-28288 => x"C0C0BFA480A48080",
-28287 => x"C0C0BFA480A480F8",
-28286 => x"C0C0BFA480A48082",
-28285 => x"C0C0BFA480A48092",
-28284 => x"C0C0BFA480A48099",
-28283 => x"C0C0BFA480A480B0",
-28282 => x"C0C0BFA480A480A4",
-28281 => x"C0C0BFA480A480F9",
-28280 => x"C0C0BFA480A480C0",
-28279 => x"C0C0BFA480A4F890",
-28278 => x"C0C0BFA480A4F880",
-28277 => x"C0C0BFA480A4F8F8",
-28276 => x"C0C0BFA480A4F882",
-28275 => x"C0C0BFA480A4F892",
-28274 => x"C0C0BFA480A4F899",
-28273 => x"C0C0BFA480A4F8B0",
-28272 => x"C0C0BFA480A4F8A4",
-28271 => x"C0C0BFA480A4F8F9",
-28270 => x"C0C0BFA480A4F8C0",
-28269 => x"C0C0BFA480A48290",
-28268 => x"C0C0BFA480A48280",
-28267 => x"C0C0BFA480A482F8",
-28266 => x"C0C0BFA480A48282",
-28265 => x"C0C0BFA480A48292",
-28264 => x"C0C0BFA480A48299",
-28263 => x"C0C0BFA480A482B0",
-28262 => x"C0C0BFA480A482A4",
-28261 => x"C0C0BFA480A482F9",
-28260 => x"C0C0BFA480A482C0",
-28259 => x"C0C0BFA480A49290",
-28258 => x"C0C0BFA480A49280",
-28257 => x"C0C0BFA480A492F8",
-28256 => x"C0C0BFA480A49282",
-28255 => x"C0C0BFA480A49292",
-28254 => x"C0C0BFA480A49299",
-28253 => x"C0C0BFA480A492B0",
-28252 => x"C0C0BFA480A492A4",
-28251 => x"C0C0BFA480A492F9",
-28250 => x"C0C0BFA480A492C0",
-28249 => x"C0C0BFA480A49990",
-28248 => x"C0C0BFA480A49980",
-28247 => x"C0C0BFA480A499F8",
-28246 => x"C0C0BFA480A49982",
-28245 => x"C0C0BFA480A49992",
-28244 => x"C0C0BFA480A49999",
-28243 => x"C0C0BFA480A499B0",
-28242 => x"C0C0BFA480A499A4",
-28241 => x"C0C0BFA480A499F9",
-28240 => x"C0C0BFA480A499C0",
-28239 => x"C0C0BFA480A4B090",
-28238 => x"C0C0BFA480A4B080",
-28237 => x"C0C0BFA480A4B0F8",
-28236 => x"C0C0BFA480A4B082",
-28235 => x"C0C0BFA480A4B092",
-28234 => x"C0C0BFA480A4B099",
-28233 => x"C0C0BFA480A4B0B0",
-28232 => x"C0C0BFA480A4B0A4",
-28231 => x"C0C0BFA480A4B0F9",
-28230 => x"C0C0BFA480A4B0C0",
-28229 => x"C0C0BFA480A4A490",
-28228 => x"C0C0BFA480A4A480",
-28227 => x"C0C0BFA480A4A4F8",
-28226 => x"C0C0BFA480A4A482",
-28225 => x"C0C0BFA480A4A492",
-28224 => x"C0C0BFA480A4A499",
-28223 => x"C0C0BFA480A4A4B0",
-28222 => x"C0C0BFA480A4A4A4",
-28221 => x"C0C0BFA480A4A4F9",
-28220 => x"C0C0BFA480A4A4C0",
-28219 => x"C0C0BFA480A4F990",
-28218 => x"C0C0BFA480A4F980",
-28217 => x"C0C0BFA480A4F9F8",
-28216 => x"C0C0BFA480A4F982",
-28215 => x"C0C0BFA480A4F992",
-28214 => x"C0C0BFA480A4F999",
-28213 => x"C0C0BFA480A4F9B0",
-28212 => x"C0C0BFA480A4F9A4",
-28211 => x"C0C0BFA480A4F9F9",
-28210 => x"C0C0BFA480A4F9C0",
-28209 => x"C0C0BFA480A4C090",
-28208 => x"C0C0BFA480A4C080",
-28207 => x"C0C0BFA480A4C0F8",
-28206 => x"C0C0BFA480A4C082",
-28205 => x"C0C0BFA480A4C092",
-28204 => x"C0C0BFA480A4C099",
-28203 => x"C0C0BFA480A4C0B0",
-28202 => x"C0C0BFA480A4C0A4",
-28201 => x"C0C0BFA480A4C0F9",
-28200 => x"C0C0BFA480A4C0C0",
-28199 => x"C0C0BFA480F99090",
-28198 => x"C0C0BFA480F99080",
-28197 => x"C0C0BFA480F990F8",
-28196 => x"C0C0BFA480F99082",
-28195 => x"C0C0BFA480F99092",
-28194 => x"C0C0BFA480F99099",
-28193 => x"C0C0BFA480F990B0",
-28192 => x"C0C0BFA480F990A4",
-28191 => x"C0C0BFA480F990F9",
-28190 => x"C0C0BFA480F990C0",
-28189 => x"C0C0BFA480F98090",
-28188 => x"C0C0BFA480F98080",
-28187 => x"C0C0BFA480F980F8",
-28186 => x"C0C0BFA480F98082",
-28185 => x"C0C0BFA480F98092",
-28184 => x"C0C0BFA480F98099",
-28183 => x"C0C0BFA480F980B0",
-28182 => x"C0C0BFA480F980A4",
-28181 => x"C0C0BFA480F980F9",
-28180 => x"C0C0BFA480F980C0",
-28179 => x"C0C0BFA480F9F890",
-28178 => x"C0C0BFA480F9F880",
-28177 => x"C0C0BFA480F9F8F8",
-28176 => x"C0C0BFA480F9F882",
-28175 => x"C0C0BFA480F9F892",
-28174 => x"C0C0BFA480F9F899",
-28173 => x"C0C0BFA480F9F8B0",
-28172 => x"C0C0BFA480F9F8A4",
-28171 => x"C0C0BFA480F9F8F9",
-28170 => x"C0C0BFA480F9F8C0",
-28169 => x"C0C0BFA480F98290",
-28168 => x"C0C0BFA480F98280",
-28167 => x"C0C0BFA480F982F8",
-28166 => x"C0C0BFA480F98282",
-28165 => x"C0C0BFA480F98292",
-28164 => x"C0C0BFA480F98299",
-28163 => x"C0C0BFA480F982B0",
-28162 => x"C0C0BFA480F982A4",
-28161 => x"C0C0BFA480F982F9",
-28160 => x"C0C0BFA480F982C0",
-28159 => x"C0C0BFA480F99290",
-28158 => x"C0C0BFA480F99280",
-28157 => x"C0C0BFA480F992F8",
-28156 => x"C0C0BFA480F99282",
-28155 => x"C0C0BFA480F99292",
-28154 => x"C0C0BFA480F99299",
-28153 => x"C0C0BFA480F992B0",
-28152 => x"C0C0BFA480F992A4",
-28151 => x"C0C0BFA480F992F9",
-28150 => x"C0C0BFA480F992C0",
-28149 => x"C0C0BFA480F99990",
-28148 => x"C0C0BFA480F99980",
-28147 => x"C0C0BFA480F999F8",
-28146 => x"C0C0BFA480F99982",
-28145 => x"C0C0BFA480F99992",
-28144 => x"C0C0BFA480F99999",
-28143 => x"C0C0BFA480F999B0",
-28142 => x"C0C0BFA480F999A4",
-28141 => x"C0C0BFA480F999F9",
-28140 => x"C0C0BFA480F999C0",
-28139 => x"C0C0BFA480F9B090",
-28138 => x"C0C0BFA480F9B080",
-28137 => x"C0C0BFA480F9B0F8",
-28136 => x"C0C0BFA480F9B082",
-28135 => x"C0C0BFA480F9B092",
-28134 => x"C0C0BFA480F9B099",
-28133 => x"C0C0BFA480F9B0B0",
-28132 => x"C0C0BFA480F9B0A4",
-28131 => x"C0C0BFA480F9B0F9",
-28130 => x"C0C0BFA480F9B0C0",
-28129 => x"C0C0BFA480F9A490",
-28128 => x"C0C0BFA480F9A480",
-28127 => x"C0C0BFA480F9A4F8",
-28126 => x"C0C0BFA480F9A482",
-28125 => x"C0C0BFA480F9A492",
-28124 => x"C0C0BFA480F9A499",
-28123 => x"C0C0BFA480F9A4B0",
-28122 => x"C0C0BFA480F9A4A4",
-28121 => x"C0C0BFA480F9A4F9",
-28120 => x"C0C0BFA480F9A4C0",
-28119 => x"C0C0BFA480F9F990",
-28118 => x"C0C0BFA480F9F980",
-28117 => x"C0C0BFA480F9F9F8",
-28116 => x"C0C0BFA480F9F982",
-28115 => x"C0C0BFA480F9F992",
-28114 => x"C0C0BFA480F9F999",
-28113 => x"C0C0BFA480F9F9B0",
-28112 => x"C0C0BFA480F9F9A4",
-28111 => x"C0C0BFA480F9F9F9",
-28110 => x"C0C0BFA480F9F9C0",
-28109 => x"C0C0BFA480F9C090",
-28108 => x"C0C0BFA480F9C080",
-28107 => x"C0C0BFA480F9C0F8",
-28106 => x"C0C0BFA480F9C082",
-28105 => x"C0C0BFA480F9C092",
-28104 => x"C0C0BFA480F9C099",
-28103 => x"C0C0BFA480F9C0B0",
-28102 => x"C0C0BFA480F9C0A4",
-28101 => x"C0C0BFA480F9C0F9",
-28100 => x"C0C0BFA480F9C0C0",
-28099 => x"C0C0BFA480C09090",
-28098 => x"C0C0BFA480C09080",
-28097 => x"C0C0BFA480C090F8",
-28096 => x"C0C0BFA480C09082",
-28095 => x"C0C0BFA480C09092",
-28094 => x"C0C0BFA480C09099",
-28093 => x"C0C0BFA480C090B0",
-28092 => x"C0C0BFA480C090A4",
-28091 => x"C0C0BFA480C090F9",
-28090 => x"C0C0BFA480C090C0",
-28089 => x"C0C0BFA480C08090",
-28088 => x"C0C0BFA480C08080",
-28087 => x"C0C0BFA480C080F8",
-28086 => x"C0C0BFA480C08082",
-28085 => x"C0C0BFA480C08092",
-28084 => x"C0C0BFA480C08099",
-28083 => x"C0C0BFA480C080B0",
-28082 => x"C0C0BFA480C080A4",
-28081 => x"C0C0BFA480C080F9",
-28080 => x"C0C0BFA480C080C0",
-28079 => x"C0C0BFA480C0F890",
-28078 => x"C0C0BFA480C0F880",
-28077 => x"C0C0BFA480C0F8F8",
-28076 => x"C0C0BFA480C0F882",
-28075 => x"C0C0BFA480C0F892",
-28074 => x"C0C0BFA480C0F899",
-28073 => x"C0C0BFA480C0F8B0",
-28072 => x"C0C0BFA480C0F8A4",
-28071 => x"C0C0BFA480C0F8F9",
-28070 => x"C0C0BFA480C0F8C0",
-28069 => x"C0C0BFA480C08290",
-28068 => x"C0C0BFA480C08280",
-28067 => x"C0C0BFA480C082F8",
-28066 => x"C0C0BFA480C08282",
-28065 => x"C0C0BFA480C08292",
-28064 => x"C0C0BFA480C08299",
-28063 => x"C0C0BFA480C082B0",
-28062 => x"C0C0BFA480C082A4",
-28061 => x"C0C0BFA480C082F9",
-28060 => x"C0C0BFA480C082C0",
-28059 => x"C0C0BFA480C09290",
-28058 => x"C0C0BFA480C09280",
-28057 => x"C0C0BFA480C092F8",
-28056 => x"C0C0BFA480C09282",
-28055 => x"C0C0BFA480C09292",
-28054 => x"C0C0BFA480C09299",
-28053 => x"C0C0BFA480C092B0",
-28052 => x"C0C0BFA480C092A4",
-28051 => x"C0C0BFA480C092F9",
-28050 => x"C0C0BFA480C092C0",
-28049 => x"C0C0BFA480C09990",
-28048 => x"C0C0BFA480C09980",
-28047 => x"C0C0BFA480C099F8",
-28046 => x"C0C0BFA480C09982",
-28045 => x"C0C0BFA480C09992",
-28044 => x"C0C0BFA480C09999",
-28043 => x"C0C0BFA480C099B0",
-28042 => x"C0C0BFA480C099A4",
-28041 => x"C0C0BFA480C099F9",
-28040 => x"C0C0BFA480C099C0",
-28039 => x"C0C0BFA480C0B090",
-28038 => x"C0C0BFA480C0B080",
-28037 => x"C0C0BFA480C0B0F8",
-28036 => x"C0C0BFA480C0B082",
-28035 => x"C0C0BFA480C0B092",
-28034 => x"C0C0BFA480C0B099",
-28033 => x"C0C0BFA480C0B0B0",
-28032 => x"C0C0BFA480C0B0A4",
-28031 => x"C0C0BFA480C0B0F9",
-28030 => x"C0C0BFA480C0B0C0",
-28029 => x"C0C0BFA480C0A490",
-28028 => x"C0C0BFA480C0A480",
-28027 => x"C0C0BFA480C0A4F8",
-28026 => x"C0C0BFA480C0A482",
-28025 => x"C0C0BFA480C0A492",
-28024 => x"C0C0BFA480C0A499",
-28023 => x"C0C0BFA480C0A4B0",
-28022 => x"C0C0BFA480C0A4A4",
-28021 => x"C0C0BFA480C0A4F9",
-28020 => x"C0C0BFA480C0A4C0",
-28019 => x"C0C0BFA480C0F990",
-28018 => x"C0C0BFA480C0F980",
-28017 => x"C0C0BFA480C0F9F8",
-28016 => x"C0C0BFA480C0F982",
-28015 => x"C0C0BFA480C0F992",
-28014 => x"C0C0BFA480C0F999",
-28013 => x"C0C0BFA480C0F9B0",
-28012 => x"C0C0BFA480C0F9A4",
-28011 => x"C0C0BFA480C0F9F9",
-28010 => x"C0C0BFA480C0F9C0",
-28009 => x"C0C0BFA480C0C090",
-28008 => x"C0C0BFA480C0C080",
-28007 => x"C0C0BFA480C0C0F8",
-28006 => x"C0C0BFA480C0C082",
-28005 => x"C0C0BFA480C0C092",
-28004 => x"C0C0BFA480C0C099",
-28003 => x"C0C0BFA480C0C0B0",
-28002 => x"C0C0BFA480C0C0A4",
-28001 => x"C0C0BFA480C0C0F9",
-28000 => x"C0C0BFA480C0C0C0",
-27999 => x"C0C0BFA4F8909090",
-27998 => x"C0C0BFA4F8909080",
-27997 => x"C0C0BFA4F89090F8",
-27996 => x"C0C0BFA4F8909082",
-27995 => x"C0C0BFA4F8909092",
-27994 => x"C0C0BFA4F8909099",
-27993 => x"C0C0BFA4F89090B0",
-27992 => x"C0C0BFA4F89090A4",
-27991 => x"C0C0BFA4F89090F9",
-27990 => x"C0C0BFA4F89090C0",
-27989 => x"C0C0BFA4F8908090",
-27988 => x"C0C0BFA4F8908080",
-27987 => x"C0C0BFA4F89080F8",
-27986 => x"C0C0BFA4F8908082",
-27985 => x"C0C0BFA4F8908092",
-27984 => x"C0C0BFA4F8908099",
-27983 => x"C0C0BFA4F89080B0",
-27982 => x"C0C0BFA4F89080A4",
-27981 => x"C0C0BFA4F89080F9",
-27980 => x"C0C0BFA4F89080C0",
-27979 => x"C0C0BFA4F890F890",
-27978 => x"C0C0BFA4F890F880",
-27977 => x"C0C0BFA4F890F8F8",
-27976 => x"C0C0BFA4F890F882",
-27975 => x"C0C0BFA4F890F892",
-27974 => x"C0C0BFA4F890F899",
-27973 => x"C0C0BFA4F890F8B0",
-27972 => x"C0C0BFA4F890F8A4",
-27971 => x"C0C0BFA4F890F8F9",
-27970 => x"C0C0BFA4F890F8C0",
-27969 => x"C0C0BFA4F8908290",
-27968 => x"C0C0BFA4F8908280",
-27967 => x"C0C0BFA4F89082F8",
-27966 => x"C0C0BFA4F8908282",
-27965 => x"C0C0BFA4F8908292",
-27964 => x"C0C0BFA4F8908299",
-27963 => x"C0C0BFA4F89082B0",
-27962 => x"C0C0BFA4F89082A4",
-27961 => x"C0C0BFA4F89082F9",
-27960 => x"C0C0BFA4F89082C0",
-27959 => x"C0C0BFA4F8909290",
-27958 => x"C0C0BFA4F8909280",
-27957 => x"C0C0BFA4F89092F8",
-27956 => x"C0C0BFA4F8909282",
-27955 => x"C0C0BFA4F8909292",
-27954 => x"C0C0BFA4F8909299",
-27953 => x"C0C0BFA4F89092B0",
-27952 => x"C0C0BFA4F89092A4",
-27951 => x"C0C0BFA4F89092F9",
-27950 => x"C0C0BFA4F89092C0",
-27949 => x"C0C0BFA4F8909990",
-27948 => x"C0C0BFA4F8909980",
-27947 => x"C0C0BFA4F89099F8",
-27946 => x"C0C0BFA4F8909982",
-27945 => x"C0C0BFA4F8909992",
-27944 => x"C0C0BFA4F8909999",
-27943 => x"C0C0BFA4F89099B0",
-27942 => x"C0C0BFA4F89099A4",
-27941 => x"C0C0BFA4F89099F9",
-27940 => x"C0C0BFA4F89099C0",
-27939 => x"C0C0BFA4F890B090",
-27938 => x"C0C0BFA4F890B080",
-27937 => x"C0C0BFA4F890B0F8",
-27936 => x"C0C0BFA4F890B082",
-27935 => x"C0C0BFA4F890B092",
-27934 => x"C0C0BFA4F890B099",
-27933 => x"C0C0BFA4F890B0B0",
-27932 => x"C0C0BFA4F890B0A4",
-27931 => x"C0C0BFA4F890B0F9",
-27930 => x"C0C0BFA4F890B0C0",
-27929 => x"C0C0BFA4F890A490",
-27928 => x"C0C0BFA4F890A480",
-27927 => x"C0C0BFA4F890A4F8",
-27926 => x"C0C0BFA4F890A482",
-27925 => x"C0C0BFA4F890A492",
-27924 => x"C0C0BFA4F890A499",
-27923 => x"C0C0BFA4F890A4B0",
-27922 => x"C0C0BFA4F890A4A4",
-27921 => x"C0C0BFA4F890A4F9",
-27920 => x"C0C0BFA4F890A4C0",
-27919 => x"C0C0BFA4F890F990",
-27918 => x"C0C0BFA4F890F980",
-27917 => x"C0C0BFA4F890F9F8",
-27916 => x"C0C0BFA4F890F982",
-27915 => x"C0C0BFA4F890F992",
-27914 => x"C0C0BFA4F890F999",
-27913 => x"C0C0BFA4F890F9B0",
-27912 => x"C0C0BFA4F890F9A4",
-27911 => x"C0C0BFA4F890F9F9",
-27910 => x"C0C0BFA4F890F9C0",
-27909 => x"C0C0BFA4F890C090",
-27908 => x"C0C0BFA4F890C080",
-27907 => x"C0C0BFA4F890C0F8",
-27906 => x"C0C0BFA4F890C082",
-27905 => x"C0C0BFA4F890C092",
-27904 => x"C0C0BFA4F890C099",
-27903 => x"C0C0BFA4F890C0B0",
-27902 => x"C0C0BFA4F890C0A4",
-27901 => x"C0C0BFA4F890C0F9",
-27900 => x"C0C0BFA4F890C0C0",
-27899 => x"C0C0BFA4F8809090",
-27898 => x"C0C0BFA4F8809080",
-27897 => x"C0C0BFA4F88090F8",
-27896 => x"C0C0BFA4F8809082",
-27895 => x"C0C0BFA4F8809092",
-27894 => x"C0C0BFA4F8809099",
-27893 => x"C0C0BFA4F88090B0",
-27892 => x"C0C0BFA4F88090A4",
-27891 => x"C0C0BFA4F88090F9",
-27890 => x"C0C0BFA4F88090C0",
-27889 => x"C0C0BFA4F8808090",
-27888 => x"C0C0BFA4F8808080",
-27887 => x"C0C0BFA4F88080F8",
-27886 => x"C0C0BFA4F8808082",
-27885 => x"C0C0BFA4F8808092",
-27884 => x"C0C0BFA4F8808099",
-27883 => x"C0C0BFA4F88080B0",
-27882 => x"C0C0BFA4F88080A4",
-27881 => x"C0C0BFA4F88080F9",
-27880 => x"C0C0BFA4F88080C0",
-27879 => x"C0C0BFA4F880F890",
-27878 => x"C0C0BFA4F880F880",
-27877 => x"C0C0BFA4F880F8F8",
-27876 => x"C0C0BFA4F880F882",
-27875 => x"C0C0BFA4F880F892",
-27874 => x"C0C0BFA4F880F899",
-27873 => x"C0C0BFA4F880F8B0",
-27872 => x"C0C0BFA4F880F8A4",
-27871 => x"C0C0BFA4F880F8F9",
-27870 => x"C0C0BFA4F880F8C0",
-27869 => x"C0C0BFA4F8808290",
-27868 => x"C0C0BFA4F8808280",
-27867 => x"C0C0BFA4F88082F8",
-27866 => x"C0C0BFA4F8808282",
-27865 => x"C0C0BFA4F8808292",
-27864 => x"C0C0BFA4F8808299",
-27863 => x"C0C0BFA4F88082B0",
-27862 => x"C0C0BFA4F88082A4",
-27861 => x"C0C0BFA4F88082F9",
-27860 => x"C0C0BFA4F88082C0",
-27859 => x"C0C0BFA4F8809290",
-27858 => x"C0C0BFA4F8809280",
-27857 => x"C0C0BFA4F88092F8",
-27856 => x"C0C0BFA4F8809282",
-27855 => x"C0C0BFA4F8809292",
-27854 => x"C0C0BFA4F8809299",
-27853 => x"C0C0BFA4F88092B0",
-27852 => x"C0C0BFA4F88092A4",
-27851 => x"C0C0BFA4F88092F9",
-27850 => x"C0C0BFA4F88092C0",
-27849 => x"C0C0BFA4F8809990",
-27848 => x"C0C0BFA4F8809980",
-27847 => x"C0C0BFA4F88099F8",
-27846 => x"C0C0BFA4F8809982",
-27845 => x"C0C0BFA4F8809992",
-27844 => x"C0C0BFA4F8809999",
-27843 => x"C0C0BFA4F88099B0",
-27842 => x"C0C0BFA4F88099A4",
-27841 => x"C0C0BFA4F88099F9",
-27840 => x"C0C0BFA4F88099C0",
-27839 => x"C0C0BFA4F880B090",
-27838 => x"C0C0BFA4F880B080",
-27837 => x"C0C0BFA4F880B0F8",
-27836 => x"C0C0BFA4F880B082",
-27835 => x"C0C0BFA4F880B092",
-27834 => x"C0C0BFA4F880B099",
-27833 => x"C0C0BFA4F880B0B0",
-27832 => x"C0C0BFA4F880B0A4",
-27831 => x"C0C0BFA4F880B0F9",
-27830 => x"C0C0BFA4F880B0C0",
-27829 => x"C0C0BFA4F880A490",
-27828 => x"C0C0BFA4F880A480",
-27827 => x"C0C0BFA4F880A4F8",
-27826 => x"C0C0BFA4F880A482",
-27825 => x"C0C0BFA4F880A492",
-27824 => x"C0C0BFA4F880A499",
-27823 => x"C0C0BFA4F880A4B0",
-27822 => x"C0C0BFA4F880A4A4",
-27821 => x"C0C0BFA4F880A4F9",
-27820 => x"C0C0BFA4F880A4C0",
-27819 => x"C0C0BFA4F880F990",
-27818 => x"C0C0BFA4F880F980",
-27817 => x"C0C0BFA4F880F9F8",
-27816 => x"C0C0BFA4F880F982",
-27815 => x"C0C0BFA4F880F992",
-27814 => x"C0C0BFA4F880F999",
-27813 => x"C0C0BFA4F880F9B0",
-27812 => x"C0C0BFA4F880F9A4",
-27811 => x"C0C0BFA4F880F9F9",
-27810 => x"C0C0BFA4F880F9C0",
-27809 => x"C0C0BFA4F880C090",
-27808 => x"C0C0BFA4F880C080",
-27807 => x"C0C0BFA4F880C0F8",
-27806 => x"C0C0BFA4F880C082",
-27805 => x"C0C0BFA4F880C092",
-27804 => x"C0C0BFA4F880C099",
-27803 => x"C0C0BFA4F880C0B0",
-27802 => x"C0C0BFA4F880C0A4",
-27801 => x"C0C0BFA4F880C0F9",
-27800 => x"C0C0BFA4F880C0C0",
-27799 => x"C0C0BFA4F8F89090",
-27798 => x"C0C0BFA4F8F89080",
-27797 => x"C0C0BFA4F8F890F8",
-27796 => x"C0C0BFA4F8F89082",
-27795 => x"C0C0BFA4F8F89092",
-27794 => x"C0C0BFA4F8F89099",
-27793 => x"C0C0BFA4F8F890B0",
-27792 => x"C0C0BFA4F8F890A4",
-27791 => x"C0C0BFA4F8F890F9",
-27790 => x"C0C0BFA4F8F890C0",
-27789 => x"C0C0BFA4F8F88090",
-27788 => x"C0C0BFA4F8F88080",
-27787 => x"C0C0BFA4F8F880F8",
-27786 => x"C0C0BFA4F8F88082",
-27785 => x"C0C0BFA4F8F88092",
-27784 => x"C0C0BFA4F8F88099",
-27783 => x"C0C0BFA4F8F880B0",
-27782 => x"C0C0BFA4F8F880A4",
-27781 => x"C0C0BFA4F8F880F9",
-27780 => x"C0C0BFA4F8F880C0",
-27779 => x"C0C0BFA4F8F8F890",
-27778 => x"C0C0BFA4F8F8F880",
-27777 => x"C0C0BFA4F8F8F8F8",
-27776 => x"C0C0BFA4F8F8F882",
-27775 => x"C0C0BFA4F8F8F892",
-27774 => x"C0C0BFA4F8F8F899",
-27773 => x"C0C0BFA4F8F8F8B0",
-27772 => x"C0C0BFA4F8F8F8A4",
-27771 => x"C0C0BFA4F8F8F8F9",
-27770 => x"C0C0BFA4F8F8F8C0",
-27769 => x"C0C0BFA4F8F88290",
-27768 => x"C0C0BFA4F8F88280",
-27767 => x"C0C0BFA4F8F882F8",
-27766 => x"C0C0BFA4F8F88282",
-27765 => x"C0C0BFA4F8F88292",
-27764 => x"C0C0BFA4F8F88299",
-27763 => x"C0C0BFA4F8F882B0",
-27762 => x"C0C0BFA4F8F882A4",
-27761 => x"C0C0BFA4F8F882F9",
-27760 => x"C0C0BFA4F8F882C0",
-27759 => x"C0C0BFA4F8F89290",
-27758 => x"C0C0BFA4F8F89280",
-27757 => x"C0C0BFA4F8F892F8",
-27756 => x"C0C0BFA4F8F89282",
-27755 => x"C0C0BFA4F8F89292",
-27754 => x"C0C0BFA4F8F89299",
-27753 => x"C0C0BFA4F8F892B0",
-27752 => x"C0C0BFA4F8F892A4",
-27751 => x"C0C0BFA4F8F892F9",
-27750 => x"C0C0BFA4F8F892C0",
-27749 => x"C0C0BFA4F8F89990",
-27748 => x"C0C0BFA4F8F89980",
-27747 => x"C0C0BFA4F8F899F8",
-27746 => x"C0C0BFA4F8F89982",
-27745 => x"C0C0BFA4F8F89992",
-27744 => x"C0C0BFA4F8F89999",
-27743 => x"C0C0BFA4F8F899B0",
-27742 => x"C0C0BFA4F8F899A4",
-27741 => x"C0C0BFA4F8F899F9",
-27740 => x"C0C0BFA4F8F899C0",
-27739 => x"C0C0BFA4F8F8B090",
-27738 => x"C0C0BFA4F8F8B080",
-27737 => x"C0C0BFA4F8F8B0F8",
-27736 => x"C0C0BFA4F8F8B082",
-27735 => x"C0C0BFA4F8F8B092",
-27734 => x"C0C0BFA4F8F8B099",
-27733 => x"C0C0BFA4F8F8B0B0",
-27732 => x"C0C0BFA4F8F8B0A4",
-27731 => x"C0C0BFA4F8F8B0F9",
-27730 => x"C0C0BFA4F8F8B0C0",
-27729 => x"C0C0BFA4F8F8A490",
-27728 => x"C0C0BFA4F8F8A480",
-27727 => x"C0C0BFA4F8F8A4F8",
-27726 => x"C0C0BFA4F8F8A482",
-27725 => x"C0C0BFA4F8F8A492",
-27724 => x"C0C0BFA4F8F8A499",
-27723 => x"C0C0BFA4F8F8A4B0",
-27722 => x"C0C0BFA4F8F8A4A4",
-27721 => x"C0C0BFA4F8F8A4F9",
-27720 => x"C0C0BFA4F8F8A4C0",
-27719 => x"C0C0BFA4F8F8F990",
-27718 => x"C0C0BFA4F8F8F980",
-27717 => x"C0C0BFA4F8F8F9F8",
-27716 => x"C0C0BFA4F8F8F982",
-27715 => x"C0C0BFA4F8F8F992",
-27714 => x"C0C0BFA4F8F8F999",
-27713 => x"C0C0BFA4F8F8F9B0",
-27712 => x"C0C0BFA4F8F8F9A4",
-27711 => x"C0C0BFA4F8F8F9F9",
-27710 => x"C0C0BFA4F8F8F9C0",
-27709 => x"C0C0BFA4F8F8C090",
-27708 => x"C0C0BFA4F8F8C080",
-27707 => x"C0C0BFA4F8F8C0F8",
-27706 => x"C0C0BFA4F8F8C082",
-27705 => x"C0C0BFA4F8F8C092",
-27704 => x"C0C0BFA4F8F8C099",
-27703 => x"C0C0BFA4F8F8C0B0",
-27702 => x"C0C0BFA4F8F8C0A4",
-27701 => x"C0C0BFA4F8F8C0F9",
-27700 => x"C0C0BFA4F8F8C0C0",
-27699 => x"C0C0BFA4F8829090",
-27698 => x"C0C0BFA4F8829080",
-27697 => x"C0C0BFA4F88290F8",
-27696 => x"C0C0BFA4F8829082",
-27695 => x"C0C0BFA4F8829092",
-27694 => x"C0C0BFA4F8829099",
-27693 => x"C0C0BFA4F88290B0",
-27692 => x"C0C0BFA4F88290A4",
-27691 => x"C0C0BFA4F88290F9",
-27690 => x"C0C0BFA4F88290C0",
-27689 => x"C0C0BFA4F8828090",
-27688 => x"C0C0BFA4F8828080",
-27687 => x"C0C0BFA4F88280F8",
-27686 => x"C0C0BFA4F8828082",
-27685 => x"C0C0BFA4F8828092",
-27684 => x"C0C0BFA4F8828099",
-27683 => x"C0C0BFA4F88280B0",
-27682 => x"C0C0BFA4F88280A4",
-27681 => x"C0C0BFA4F88280F9",
-27680 => x"C0C0BFA4F88280C0",
-27679 => x"C0C0BFA4F882F890",
-27678 => x"C0C0BFA4F882F880",
-27677 => x"C0C0BFA4F882F8F8",
-27676 => x"C0C0BFA4F882F882",
-27675 => x"C0C0BFA4F882F892",
-27674 => x"C0C0BFA4F882F899",
-27673 => x"C0C0BFA4F882F8B0",
-27672 => x"C0C0BFA4F882F8A4",
-27671 => x"C0C0BFA4F882F8F9",
-27670 => x"C0C0BFA4F882F8C0",
-27669 => x"C0C0BFA4F8828290",
-27668 => x"C0C0BFA4F8828280",
-27667 => x"C0C0BFA4F88282F8",
-27666 => x"C0C0BFA4F8828282",
-27665 => x"C0C0BFA4F8828292",
-27664 => x"C0C0BFA4F8828299",
-27663 => x"C0C0BFA4F88282B0",
-27662 => x"C0C0BFA4F88282A4",
-27661 => x"C0C0BFA4F88282F9",
-27660 => x"C0C0BFA4F88282C0",
-27659 => x"C0C0BFA4F8829290",
-27658 => x"C0C0BFA4F8829280",
-27657 => x"C0C0BFA4F88292F8",
-27656 => x"C0C0BFA4F8829282",
-27655 => x"C0C0BFA4F8829292",
-27654 => x"C0C0BFA4F8829299",
-27653 => x"C0C0BFA4F88292B0",
-27652 => x"C0C0BFA4F88292A4",
-27651 => x"C0C0BFA4F88292F9",
-27650 => x"C0C0BFA4F88292C0",
-27649 => x"C0C0BFA4F8829990",
-27648 => x"C0C0BFA4F8829980",
-27647 => x"C0C0BFA4F88299F8",
-27646 => x"C0C0BFA4F8829982",
-27645 => x"C0C0BFA4F8829992",
-27644 => x"C0C0BFA4F8829999",
-27643 => x"C0C0BFA4F88299B0",
-27642 => x"C0C0BFA4F88299A4",
-27641 => x"C0C0BFA4F88299F9",
-27640 => x"C0C0BFA4F88299C0",
-27639 => x"C0C0BFA4F882B090",
-27638 => x"C0C0BFA4F882B080",
-27637 => x"C0C0BFA4F882B0F8",
-27636 => x"C0C0BFA4F882B082",
-27635 => x"C0C0BFA4F882B092",
-27634 => x"C0C0BFA4F882B099",
-27633 => x"C0C0BFA4F882B0B0",
-27632 => x"C0C0BFA4F882B0A4",
-27631 => x"C0C0BFA4F882B0F9",
-27630 => x"C0C0BFA4F882B0C0",
-27629 => x"C0C0BFA4F882A490",
-27628 => x"C0C0BFA4F882A480",
-27627 => x"C0C0BFA4F882A4F8",
-27626 => x"C0C0BFA4F882A482",
-27625 => x"C0C0BFA4F882A492",
-27624 => x"C0C0BFA4F882A499",
-27623 => x"C0C0BFA4F882A4B0",
-27622 => x"C0C0BFA4F882A4A4",
-27621 => x"C0C0BFA4F882A4F9",
-27620 => x"C0C0BFA4F882A4C0",
-27619 => x"C0C0BFA4F882F990",
-27618 => x"C0C0BFA4F882F980",
-27617 => x"C0C0BFA4F882F9F8",
-27616 => x"C0C0BFA4F882F982",
-27615 => x"C0C0BFA4F882F992",
-27614 => x"C0C0BFA4F882F999",
-27613 => x"C0C0BFA4F882F9B0",
-27612 => x"C0C0BFA4F882F9A4",
-27611 => x"C0C0BFA4F882F9F9",
-27610 => x"C0C0BFA4F882F9C0",
-27609 => x"C0C0BFA4F882C090",
-27608 => x"C0C0BFA4F882C080",
-27607 => x"C0C0BFA4F882C0F8",
-27606 => x"C0C0BFA4F882C082",
-27605 => x"C0C0BFA4F882C092",
-27604 => x"C0C0BFA4F882C099",
-27603 => x"C0C0BFA4F882C0B0",
-27602 => x"C0C0BFA4F882C0A4",
-27601 => x"C0C0BFA4F882C0F9",
-27600 => x"C0C0BFA4F882C0C0",
-27599 => x"C0C0BFA4F8929090",
-27598 => x"C0C0BFA4F8929080",
-27597 => x"C0C0BFA4F89290F8",
-27596 => x"C0C0BFA4F8929082",
-27595 => x"C0C0BFA4F8929092",
-27594 => x"C0C0BFA4F8929099",
-27593 => x"C0C0BFA4F89290B0",
-27592 => x"C0C0BFA4F89290A4",
-27591 => x"C0C0BFA4F89290F9",
-27590 => x"C0C0BFA4F89290C0",
-27589 => x"C0C0BFA4F8928090",
-27588 => x"C0C0BFA4F8928080",
-27587 => x"C0C0BFA4F89280F8",
-27586 => x"C0C0BFA4F8928082",
-27585 => x"C0C0BFA4F8928092",
-27584 => x"C0C0BFA4F8928099",
-27583 => x"C0C0BFA4F89280B0",
-27582 => x"C0C0BFA4F89280A4",
-27581 => x"C0C0BFA4F89280F9",
-27580 => x"C0C0BFA4F89280C0",
-27579 => x"C0C0BFA4F892F890",
-27578 => x"C0C0BFA4F892F880",
-27577 => x"C0C0BFA4F892F8F8",
-27576 => x"C0C0BFA4F892F882",
-27575 => x"C0C0BFA4F892F892",
-27574 => x"C0C0BFA4F892F899",
-27573 => x"C0C0BFA4F892F8B0",
-27572 => x"C0C0BFA4F892F8A4",
-27571 => x"C0C0BFA4F892F8F9",
-27570 => x"C0C0BFA4F892F8C0",
-27569 => x"C0C0BFA4F8928290",
-27568 => x"C0C0BFA4F8928280",
-27567 => x"C0C0BFA4F89282F8",
-27566 => x"C0C0BFA4F8928282",
-27565 => x"C0C0BFA4F8928292",
-27564 => x"C0C0BFA4F8928299",
-27563 => x"C0C0BFA4F89282B0",
-27562 => x"C0C0BFA4F89282A4",
-27561 => x"C0C0BFA4F89282F9",
-27560 => x"C0C0BFA4F89282C0",
-27559 => x"C0C0BFA4F8929290",
-27558 => x"C0C0BFA4F8929280",
-27557 => x"C0C0BFA4F89292F8",
-27556 => x"C0C0BFA4F8929282",
-27555 => x"C0C0BFA4F8929292",
-27554 => x"C0C0BFA4F8929299",
-27553 => x"C0C0BFA4F89292B0",
-27552 => x"C0C0BFA4F89292A4",
-27551 => x"C0C0BFA4F89292F9",
-27550 => x"C0C0BFA4F89292C0",
-27549 => x"C0C0BFA4F8929990",
-27548 => x"C0C0BFA4F8929980",
-27547 => x"C0C0BFA4F89299F8",
-27546 => x"C0C0BFA4F8929982",
-27545 => x"C0C0BFA4F8929992",
-27544 => x"C0C0BFA4F8929999",
-27543 => x"C0C0BFA4F89299B0",
-27542 => x"C0C0BFA4F89299A4",
-27541 => x"C0C0BFA4F89299F9",
-27540 => x"C0C0BFA4F89299C0",
-27539 => x"C0C0BFA4F892B090",
-27538 => x"C0C0BFA4F892B080",
-27537 => x"C0C0BFA4F892B0F8",
-27536 => x"C0C0BFA4F892B082",
-27535 => x"C0C0BFA4F892B092",
-27534 => x"C0C0BFA4F892B099",
-27533 => x"C0C0BFA4F892B0B0",
-27532 => x"C0C0BFA4F892B0A4",
-27531 => x"C0C0BFA4F892B0F9",
-27530 => x"C0C0BFA4F892B0C0",
-27529 => x"C0C0BFA4F892A490",
-27528 => x"C0C0BFA4F892A480",
-27527 => x"C0C0BFA4F892A4F8",
-27526 => x"C0C0BFA4F892A482",
-27525 => x"C0C0BFA4F892A492",
-27524 => x"C0C0BFA4F892A499",
-27523 => x"C0C0BFA4F892A4B0",
-27522 => x"C0C0BFA4F892A4A4",
-27521 => x"C0C0BFA4F892A4F9",
-27520 => x"C0C0BFA4F892A4C0",
-27519 => x"C0C0BFA4F892F990",
-27518 => x"C0C0BFA4F892F980",
-27517 => x"C0C0BFA4F892F9F8",
-27516 => x"C0C0BFA4F892F982",
-27515 => x"C0C0BFA4F892F992",
-27514 => x"C0C0BFA4F892F999",
-27513 => x"C0C0BFA4F892F9B0",
-27512 => x"C0C0BFA4F892F9A4",
-27511 => x"C0C0BFA4F892F9F9",
-27510 => x"C0C0BFA4F892F9C0",
-27509 => x"C0C0BFA4F892C090",
-27508 => x"C0C0BFA4F892C080",
-27507 => x"C0C0BFA4F892C0F8",
-27506 => x"C0C0BFA4F892C082",
-27505 => x"C0C0BFA4F892C092",
-27504 => x"C0C0BFA4F892C099",
-27503 => x"C0C0BFA4F892C0B0",
-27502 => x"C0C0BFA4F892C0A4",
-27501 => x"C0C0BFA4F892C0F9",
-27500 => x"C0C0BFA4F892C0C0",
-27499 => x"C0C0BFA4F8999090",
-27498 => x"C0C0BFA4F8999080",
-27497 => x"C0C0BFA4F89990F8",
-27496 => x"C0C0BFA4F8999082",
-27495 => x"C0C0BFA4F8999092",
-27494 => x"C0C0BFA4F8999099",
-27493 => x"C0C0BFA4F89990B0",
-27492 => x"C0C0BFA4F89990A4",
-27491 => x"C0C0BFA4F89990F9",
-27490 => x"C0C0BFA4F89990C0",
-27489 => x"C0C0BFA4F8998090",
-27488 => x"C0C0BFA4F8998080",
-27487 => x"C0C0BFA4F89980F8",
-27486 => x"C0C0BFA4F8998082",
-27485 => x"C0C0BFA4F8998092",
-27484 => x"C0C0BFA4F8998099",
-27483 => x"C0C0BFA4F89980B0",
-27482 => x"C0C0BFA4F89980A4",
-27481 => x"C0C0BFA4F89980F9",
-27480 => x"C0C0BFA4F89980C0",
-27479 => x"C0C0BFA4F899F890",
-27478 => x"C0C0BFA4F899F880",
-27477 => x"C0C0BFA4F899F8F8",
-27476 => x"C0C0BFA4F899F882",
-27475 => x"C0C0BFA4F899F892",
-27474 => x"C0C0BFA4F899F899",
-27473 => x"C0C0BFA4F899F8B0",
-27472 => x"C0C0BFA4F899F8A4",
-27471 => x"C0C0BFA4F899F8F9",
-27470 => x"C0C0BFA4F899F8C0",
-27469 => x"C0C0BFA4F8998290",
-27468 => x"C0C0BFA4F8998280",
-27467 => x"C0C0BFA4F89982F8",
-27466 => x"C0C0BFA4F8998282",
-27465 => x"C0C0BFA4F8998292",
-27464 => x"C0C0BFA4F8998299",
-27463 => x"C0C0BFA4F89982B0",
-27462 => x"C0C0BFA4F89982A4",
-27461 => x"C0C0BFA4F89982F9",
-27460 => x"C0C0BFA4F89982C0",
-27459 => x"C0C0BFA4F8999290",
-27458 => x"C0C0BFA4F8999280",
-27457 => x"C0C0BFA4F89992F8",
-27456 => x"C0C0BFA4F8999282",
-27455 => x"C0C0BFA4F8999292",
-27454 => x"C0C0BFA4F8999299",
-27453 => x"C0C0BFA4F89992B0",
-27452 => x"C0C0BFA4F89992A4",
-27451 => x"C0C0BFA4F89992F9",
-27450 => x"C0C0BFA4F89992C0",
-27449 => x"C0C0BFA4F8999990",
-27448 => x"C0C0BFA4F8999980",
-27447 => x"C0C0BFA4F89999F8",
-27446 => x"C0C0BFA4F8999982",
-27445 => x"C0C0BFA4F8999992",
-27444 => x"C0C0BFA4F8999999",
-27443 => x"C0C0BFA4F89999B0",
-27442 => x"C0C0BFA4F89999A4",
-27441 => x"C0C0BFA4F89999F9",
-27440 => x"C0C0BFA4F89999C0",
-27439 => x"C0C0BFA4F899B090",
-27438 => x"C0C0BFA4F899B080",
-27437 => x"C0C0BFA4F899B0F8",
-27436 => x"C0C0BFA4F899B082",
-27435 => x"C0C0BFA4F899B092",
-27434 => x"C0C0BFA4F899B099",
-27433 => x"C0C0BFA4F899B0B0",
-27432 => x"C0C0BFA4F899B0A4",
-27431 => x"C0C0BFA4F899B0F9",
-27430 => x"C0C0BFA4F899B0C0",
-27429 => x"C0C0BFA4F899A490",
-27428 => x"C0C0BFA4F899A480",
-27427 => x"C0C0BFA4F899A4F8",
-27426 => x"C0C0BFA4F899A482",
-27425 => x"C0C0BFA4F899A492",
-27424 => x"C0C0BFA4F899A499",
-27423 => x"C0C0BFA4F899A4B0",
-27422 => x"C0C0BFA4F899A4A4",
-27421 => x"C0C0BFA4F899A4F9",
-27420 => x"C0C0BFA4F899A4C0",
-27419 => x"C0C0BFA4F899F990",
-27418 => x"C0C0BFA4F899F980",
-27417 => x"C0C0BFA4F899F9F8",
-27416 => x"C0C0BFA4F899F982",
-27415 => x"C0C0BFA4F899F992",
-27414 => x"C0C0BFA4F899F999",
-27413 => x"C0C0BFA4F899F9B0",
-27412 => x"C0C0BFA4F899F9A4",
-27411 => x"C0C0BFA4F899F9F9",
-27410 => x"C0C0BFA4F899F9C0",
-27409 => x"C0C0BFA4F899C090",
-27408 => x"C0C0BFA4F899C080",
-27407 => x"C0C0BFA4F899C0F8",
-27406 => x"C0C0BFA4F899C082",
-27405 => x"C0C0BFA4F899C092",
-27404 => x"C0C0BFA4F899C099",
-27403 => x"C0C0BFA4F899C0B0",
-27402 => x"C0C0BFA4F899C0A4",
-27401 => x"C0C0BFA4F899C0F9",
-27400 => x"C0C0BFA4F899C0C0",
-27399 => x"C0C0BFA4F8B09090",
-27398 => x"C0C0BFA4F8B09080",
-27397 => x"C0C0BFA4F8B090F8",
-27396 => x"C0C0BFA4F8B09082",
-27395 => x"C0C0BFA4F8B09092",
-27394 => x"C0C0BFA4F8B09099",
-27393 => x"C0C0BFA4F8B090B0",
-27392 => x"C0C0BFA4F8B090A4",
-27391 => x"C0C0BFA4F8B090F9",
-27390 => x"C0C0BFA4F8B090C0",
-27389 => x"C0C0BFA4F8B08090",
-27388 => x"C0C0BFA4F8B08080",
-27387 => x"C0C0BFA4F8B080F8",
-27386 => x"C0C0BFA4F8B08082",
-27385 => x"C0C0BFA4F8B08092",
-27384 => x"C0C0BFA4F8B08099",
-27383 => x"C0C0BFA4F8B080B0",
-27382 => x"C0C0BFA4F8B080A4",
-27381 => x"C0C0BFA4F8B080F9",
-27380 => x"C0C0BFA4F8B080C0",
-27379 => x"C0C0BFA4F8B0F890",
-27378 => x"C0C0BFA4F8B0F880",
-27377 => x"C0C0BFA4F8B0F8F8",
-27376 => x"C0C0BFA4F8B0F882",
-27375 => x"C0C0BFA4F8B0F892",
-27374 => x"C0C0BFA4F8B0F899",
-27373 => x"C0C0BFA4F8B0F8B0",
-27372 => x"C0C0BFA4F8B0F8A4",
-27371 => x"C0C0BFA4F8B0F8F9",
-27370 => x"C0C0BFA4F8B0F8C0",
-27369 => x"C0C0BFA4F8B08290",
-27368 => x"C0C0BFA4F8B08280",
-27367 => x"C0C0BFA4F8B082F8",
-27366 => x"C0C0BFA4F8B08282",
-27365 => x"C0C0BFA4F8B08292",
-27364 => x"C0C0BFA4F8B08299",
-27363 => x"C0C0BFA4F8B082B0",
-27362 => x"C0C0BFA4F8B082A4",
-27361 => x"C0C0BFA4F8B082F9",
-27360 => x"C0C0BFA4F8B082C0",
-27359 => x"C0C0BFA4F8B09290",
-27358 => x"C0C0BFA4F8B09280",
-27357 => x"C0C0BFA4F8B092F8",
-27356 => x"C0C0BFA4F8B09282",
-27355 => x"C0C0BFA4F8B09292",
-27354 => x"C0C0BFA4F8B09299",
-27353 => x"C0C0BFA4F8B092B0",
-27352 => x"C0C0BFA4F8B092A4",
-27351 => x"C0C0BFA4F8B092F9",
-27350 => x"C0C0BFA4F8B092C0",
-27349 => x"C0C0BFA4F8B09990",
-27348 => x"C0C0BFA4F8B09980",
-27347 => x"C0C0BFA4F8B099F8",
-27346 => x"C0C0BFA4F8B09982",
-27345 => x"C0C0BFA4F8B09992",
-27344 => x"C0C0BFA4F8B09999",
-27343 => x"C0C0BFA4F8B099B0",
-27342 => x"C0C0BFA4F8B099A4",
-27341 => x"C0C0BFA4F8B099F9",
-27340 => x"C0C0BFA4F8B099C0",
-27339 => x"C0C0BFA4F8B0B090",
-27338 => x"C0C0BFA4F8B0B080",
-27337 => x"C0C0BFA4F8B0B0F8",
-27336 => x"C0C0BFA4F8B0B082",
-27335 => x"C0C0BFA4F8B0B092",
-27334 => x"C0C0BFA4F8B0B099",
-27333 => x"C0C0BFA4F8B0B0B0",
-27332 => x"C0C0BFA4F8B0B0A4",
-27331 => x"C0C0BFA4F8B0B0F9",
-27330 => x"C0C0BFA4F8B0B0C0",
-27329 => x"C0C0BFA4F8B0A490",
-27328 => x"C0C0BFA4F8B0A480",
-27327 => x"C0C0BFA4F8B0A4F8",
-27326 => x"C0C0BFA4F8B0A482",
-27325 => x"C0C0BFA4F8B0A492",
-27324 => x"C0C0BFA4F8B0A499",
-27323 => x"C0C0BFA4F8B0A4B0",
-27322 => x"C0C0BFA4F8B0A4A4",
-27321 => x"C0C0BFA4F8B0A4F9",
-27320 => x"C0C0BFA4F8B0A4C0",
-27319 => x"C0C0BFA4F8B0F990",
-27318 => x"C0C0BFA4F8B0F980",
-27317 => x"C0C0BFA4F8B0F9F8",
-27316 => x"C0C0BFA4F8B0F982",
-27315 => x"C0C0BFA4F8B0F992",
-27314 => x"C0C0BFA4F8B0F999",
-27313 => x"C0C0BFA4F8B0F9B0",
-27312 => x"C0C0BFA4F8B0F9A4",
-27311 => x"C0C0BFA4F8B0F9F9",
-27310 => x"C0C0BFA4F8B0F9C0",
-27309 => x"C0C0BFA4F8B0C090",
-27308 => x"C0C0BFA4F8B0C080",
-27307 => x"C0C0BFA4F8B0C0F8",
-27306 => x"C0C0BFA4F8B0C082",
-27305 => x"C0C0BFA4F8B0C092",
-27304 => x"C0C0BFA4F8B0C099",
-27303 => x"C0C0BFA4F8B0C0B0",
-27302 => x"C0C0BFA4F8B0C0A4",
-27301 => x"C0C0BFA4F8B0C0F9",
-27300 => x"C0C0BFA4F8B0C0C0",
-27299 => x"C0C0BFA4F8A49090",
-27298 => x"C0C0BFA4F8A49080",
-27297 => x"C0C0BFA4F8A490F8",
-27296 => x"C0C0BFA4F8A49082",
-27295 => x"C0C0BFA4F8A49092",
-27294 => x"C0C0BFA4F8A49099",
-27293 => x"C0C0BFA4F8A490B0",
-27292 => x"C0C0BFA4F8A490A4",
-27291 => x"C0C0BFA4F8A490F9",
-27290 => x"C0C0BFA4F8A490C0",
-27289 => x"C0C0BFA4F8A48090",
-27288 => x"C0C0BFA4F8A48080",
-27287 => x"C0C0BFA4F8A480F8",
-27286 => x"C0C0BFA4F8A48082",
-27285 => x"C0C0BFA4F8A48092",
-27284 => x"C0C0BFA4F8A48099",
-27283 => x"C0C0BFA4F8A480B0",
-27282 => x"C0C0BFA4F8A480A4",
-27281 => x"C0C0BFA4F8A480F9",
-27280 => x"C0C0BFA4F8A480C0",
-27279 => x"C0C0BFA4F8A4F890",
-27278 => x"C0C0BFA4F8A4F880",
-27277 => x"C0C0BFA4F8A4F8F8",
-27276 => x"C0C0BFA4F8A4F882",
-27275 => x"C0C0BFA4F8A4F892",
-27274 => x"C0C0BFA4F8A4F899",
-27273 => x"C0C0BFA4F8A4F8B0",
-27272 => x"C0C0BFA4F8A4F8A4",
-27271 => x"C0C0BFA4F8A4F8F9",
-27270 => x"C0C0BFA4F8A4F8C0",
-27269 => x"C0C0BFA4F8A48290",
-27268 => x"C0C0BFA4F8A48280",
-27267 => x"C0C0BFA4F8A482F8",
-27266 => x"C0C0BFA4F8A48282",
-27265 => x"C0C0BFA4F8A48292",
-27264 => x"C0C0BFA4F8A48299",
-27263 => x"C0C0BFA4F8A482B0",
-27262 => x"C0C0BFA4F8A482A4",
-27261 => x"C0C0BFA4F8A482F9",
-27260 => x"C0C0BFA4F8A482C0",
-27259 => x"C0C0BFA4F8A49290",
-27258 => x"C0C0BFA4F8A49280",
-27257 => x"C0C0BFA4F8A492F8",
-27256 => x"C0C0BFA4F8A49282",
-27255 => x"C0C0BFA4F8A49292",
-27254 => x"C0C0BFA4F8A49299",
-27253 => x"C0C0BFA4F8A492B0",
-27252 => x"C0C0BFA4F8A492A4",
-27251 => x"C0C0BFA4F8A492F9",
-27250 => x"C0C0BFA4F8A492C0",
-27249 => x"C0C0BFA4F8A49990",
-27248 => x"C0C0BFA4F8A49980",
-27247 => x"C0C0BFA4F8A499F8",
-27246 => x"C0C0BFA4F8A49982",
-27245 => x"C0C0BFA4F8A49992",
-27244 => x"C0C0BFA4F8A49999",
-27243 => x"C0C0BFA4F8A499B0",
-27242 => x"C0C0BFA4F8A499A4",
-27241 => x"C0C0BFA4F8A499F9",
-27240 => x"C0C0BFA4F8A499C0",
-27239 => x"C0C0BFA4F8A4B090",
-27238 => x"C0C0BFA4F8A4B080",
-27237 => x"C0C0BFA4F8A4B0F8",
-27236 => x"C0C0BFA4F8A4B082",
-27235 => x"C0C0BFA4F8A4B092",
-27234 => x"C0C0BFA4F8A4B099",
-27233 => x"C0C0BFA4F8A4B0B0",
-27232 => x"C0C0BFA4F8A4B0A4",
-27231 => x"C0C0BFA4F8A4B0F9",
-27230 => x"C0C0BFA4F8A4B0C0",
-27229 => x"C0C0BFA4F8A4A490",
-27228 => x"C0C0BFA4F8A4A480",
-27227 => x"C0C0BFA4F8A4A4F8",
-27226 => x"C0C0BFA4F8A4A482",
-27225 => x"C0C0BFA4F8A4A492",
-27224 => x"C0C0BFA4F8A4A499",
-27223 => x"C0C0BFA4F8A4A4B0",
-27222 => x"C0C0BFA4F8A4A4A4",
-27221 => x"C0C0BFA4F8A4A4F9",
-27220 => x"C0C0BFA4F8A4A4C0",
-27219 => x"C0C0BFA4F8A4F990",
-27218 => x"C0C0BFA4F8A4F980",
-27217 => x"C0C0BFA4F8A4F9F8",
-27216 => x"C0C0BFA4F8A4F982",
-27215 => x"C0C0BFA4F8A4F992",
-27214 => x"C0C0BFA4F8A4F999",
-27213 => x"C0C0BFA4F8A4F9B0",
-27212 => x"C0C0BFA4F8A4F9A4",
-27211 => x"C0C0BFA4F8A4F9F9",
-27210 => x"C0C0BFA4F8A4F9C0",
-27209 => x"C0C0BFA4F8A4C090",
-27208 => x"C0C0BFA4F8A4C080",
-27207 => x"C0C0BFA4F8A4C0F8",
-27206 => x"C0C0BFA4F8A4C082",
-27205 => x"C0C0BFA4F8A4C092",
-27204 => x"C0C0BFA4F8A4C099",
-27203 => x"C0C0BFA4F8A4C0B0",
-27202 => x"C0C0BFA4F8A4C0A4",
-27201 => x"C0C0BFA4F8A4C0F9",
-27200 => x"C0C0BFA4F8A4C0C0",
-27199 => x"C0C0BFA4F8F99090",
-27198 => x"C0C0BFA4F8F99080",
-27197 => x"C0C0BFA4F8F990F8",
-27196 => x"C0C0BFA4F8F99082",
-27195 => x"C0C0BFA4F8F99092",
-27194 => x"C0C0BFA4F8F99099",
-27193 => x"C0C0BFA4F8F990B0",
-27192 => x"C0C0BFA4F8F990A4",
-27191 => x"C0C0BFA4F8F990F9",
-27190 => x"C0C0BFA4F8F990C0",
-27189 => x"C0C0BFA4F8F98090",
-27188 => x"C0C0BFA4F8F98080",
-27187 => x"C0C0BFA4F8F980F8",
-27186 => x"C0C0BFA4F8F98082",
-27185 => x"C0C0BFA4F8F98092",
-27184 => x"C0C0BFA4F8F98099",
-27183 => x"C0C0BFA4F8F980B0",
-27182 => x"C0C0BFA4F8F980A4",
-27181 => x"C0C0BFA4F8F980F9",
-27180 => x"C0C0BFA4F8F980C0",
-27179 => x"C0C0BFA4F8F9F890",
-27178 => x"C0C0BFA4F8F9F880",
-27177 => x"C0C0BFA4F8F9F8F8",
-27176 => x"C0C0BFA4F8F9F882",
-27175 => x"C0C0BFA4F8F9F892",
-27174 => x"C0C0BFA4F8F9F899",
-27173 => x"C0C0BFA4F8F9F8B0",
-27172 => x"C0C0BFA4F8F9F8A4",
-27171 => x"C0C0BFA4F8F9F8F9",
-27170 => x"C0C0BFA4F8F9F8C0",
-27169 => x"C0C0BFA4F8F98290",
-27168 => x"C0C0BFA4F8F98280",
-27167 => x"C0C0BFA4F8F982F8",
-27166 => x"C0C0BFA4F8F98282",
-27165 => x"C0C0BFA4F8F98292",
-27164 => x"C0C0BFA4F8F98299",
-27163 => x"C0C0BFA4F8F982B0",
-27162 => x"C0C0BFA4F8F982A4",
-27161 => x"C0C0BFA4F8F982F9",
-27160 => x"C0C0BFA4F8F982C0",
-27159 => x"C0C0BFA4F8F99290",
-27158 => x"C0C0BFA4F8F99280",
-27157 => x"C0C0BFA4F8F992F8",
-27156 => x"C0C0BFA4F8F99282",
-27155 => x"C0C0BFA4F8F99292",
-27154 => x"C0C0BFA4F8F99299",
-27153 => x"C0C0BFA4F8F992B0",
-27152 => x"C0C0BFA4F8F992A4",
-27151 => x"C0C0BFA4F8F992F9",
-27150 => x"C0C0BFA4F8F992C0",
-27149 => x"C0C0BFA4F8F99990",
-27148 => x"C0C0BFA4F8F99980",
-27147 => x"C0C0BFA4F8F999F8",
-27146 => x"C0C0BFA4F8F99982",
-27145 => x"C0C0BFA4F8F99992",
-27144 => x"C0C0BFA4F8F99999",
-27143 => x"C0C0BFA4F8F999B0",
-27142 => x"C0C0BFA4F8F999A4",
-27141 => x"C0C0BFA4F8F999F9",
-27140 => x"C0C0BFA4F8F999C0",
-27139 => x"C0C0BFA4F8F9B090",
-27138 => x"C0C0BFA4F8F9B080",
-27137 => x"C0C0BFA4F8F9B0F8",
-27136 => x"C0C0BFA4F8F9B082",
-27135 => x"C0C0BFA4F8F9B092",
-27134 => x"C0C0BFA4F8F9B099",
-27133 => x"C0C0BFA4F8F9B0B0",
-27132 => x"C0C0BFA4F8F9B0A4",
-27131 => x"C0C0BFA4F8F9B0F9",
-27130 => x"C0C0BFA4F8F9B0C0",
-27129 => x"C0C0BFA4F8F9A490",
-27128 => x"C0C0BFA4F8F9A480",
-27127 => x"C0C0BFA4F8F9A4F8",
-27126 => x"C0C0BFA4F8F9A482",
-27125 => x"C0C0BFA4F8F9A492",
-27124 => x"C0C0BFA4F8F9A499",
-27123 => x"C0C0BFA4F8F9A4B0",
-27122 => x"C0C0BFA4F8F9A4A4",
-27121 => x"C0C0BFA4F8F9A4F9",
-27120 => x"C0C0BFA4F8F9A4C0",
-27119 => x"C0C0BFA4F8F9F990",
-27118 => x"C0C0BFA4F8F9F980",
-27117 => x"C0C0BFA4F8F9F9F8",
-27116 => x"C0C0BFA4F8F9F982",
-27115 => x"C0C0BFA4F8F9F992",
-27114 => x"C0C0BFA4F8F9F999",
-27113 => x"C0C0BFA4F8F9F9B0",
-27112 => x"C0C0BFA4F8F9F9A4",
-27111 => x"C0C0BFA4F8F9F9F9",
-27110 => x"C0C0BFA4F8F9F9C0",
-27109 => x"C0C0BFA4F8F9C090",
-27108 => x"C0C0BFA4F8F9C080",
-27107 => x"C0C0BFA4F8F9C0F8",
-27106 => x"C0C0BFA4F8F9C082",
-27105 => x"C0C0BFA4F8F9C092",
-27104 => x"C0C0BFA4F8F9C099",
-27103 => x"C0C0BFA4F8F9C0B0",
-27102 => x"C0C0BFA4F8F9C0A4",
-27101 => x"C0C0BFA4F8F9C0F9",
-27100 => x"C0C0BFA4F8F9C0C0",
-27099 => x"C0C0BFA4F8C09090",
-27098 => x"C0C0BFA4F8C09080",
-27097 => x"C0C0BFA4F8C090F8",
-27096 => x"C0C0BFA4F8C09082",
-27095 => x"C0C0BFA4F8C09092",
-27094 => x"C0C0BFA4F8C09099",
-27093 => x"C0C0BFA4F8C090B0",
-27092 => x"C0C0BFA4F8C090A4",
-27091 => x"C0C0BFA4F8C090F9",
-27090 => x"C0C0BFA4F8C090C0",
-27089 => x"C0C0BFA4F8C08090",
-27088 => x"C0C0BFA4F8C08080",
-27087 => x"C0C0BFA4F8C080F8",
-27086 => x"C0C0BFA4F8C08082",
-27085 => x"C0C0BFA4F8C08092",
-27084 => x"C0C0BFA4F8C08099",
-27083 => x"C0C0BFA4F8C080B0",
-27082 => x"C0C0BFA4F8C080A4",
-27081 => x"C0C0BFA4F8C080F9",
-27080 => x"C0C0BFA4F8C080C0",
-27079 => x"C0C0BFA4F8C0F890",
-27078 => x"C0C0BFA4F8C0F880",
-27077 => x"C0C0BFA4F8C0F8F8",
-27076 => x"C0C0BFA4F8C0F882",
-27075 => x"C0C0BFA4F8C0F892",
-27074 => x"C0C0BFA4F8C0F899",
-27073 => x"C0C0BFA4F8C0F8B0",
-27072 => x"C0C0BFA4F8C0F8A4",
-27071 => x"C0C0BFA4F8C0F8F9",
-27070 => x"C0C0BFA4F8C0F8C0",
-27069 => x"C0C0BFA4F8C08290",
-27068 => x"C0C0BFA4F8C08280",
-27067 => x"C0C0BFA4F8C082F8",
-27066 => x"C0C0BFA4F8C08282",
-27065 => x"C0C0BFA4F8C08292",
-27064 => x"C0C0BFA4F8C08299",
-27063 => x"C0C0BFA4F8C082B0",
-27062 => x"C0C0BFA4F8C082A4",
-27061 => x"C0C0BFA4F8C082F9",
-27060 => x"C0C0BFA4F8C082C0",
-27059 => x"C0C0BFA4F8C09290",
-27058 => x"C0C0BFA4F8C09280",
-27057 => x"C0C0BFA4F8C092F8",
-27056 => x"C0C0BFA4F8C09282",
-27055 => x"C0C0BFA4F8C09292",
-27054 => x"C0C0BFA4F8C09299",
-27053 => x"C0C0BFA4F8C092B0",
-27052 => x"C0C0BFA4F8C092A4",
-27051 => x"C0C0BFA4F8C092F9",
-27050 => x"C0C0BFA4F8C092C0",
-27049 => x"C0C0BFA4F8C09990",
-27048 => x"C0C0BFA4F8C09980",
-27047 => x"C0C0BFA4F8C099F8",
-27046 => x"C0C0BFA4F8C09982",
-27045 => x"C0C0BFA4F8C09992",
-27044 => x"C0C0BFA4F8C09999",
-27043 => x"C0C0BFA4F8C099B0",
-27042 => x"C0C0BFA4F8C099A4",
-27041 => x"C0C0BFA4F8C099F9",
-27040 => x"C0C0BFA4F8C099C0",
-27039 => x"C0C0BFA4F8C0B090",
-27038 => x"C0C0BFA4F8C0B080",
-27037 => x"C0C0BFA4F8C0B0F8",
-27036 => x"C0C0BFA4F8C0B082",
-27035 => x"C0C0BFA4F8C0B092",
-27034 => x"C0C0BFA4F8C0B099",
-27033 => x"C0C0BFA4F8C0B0B0",
-27032 => x"C0C0BFA4F8C0B0A4",
-27031 => x"C0C0BFA4F8C0B0F9",
-27030 => x"C0C0BFA4F8C0B0C0",
-27029 => x"C0C0BFA4F8C0A490",
-27028 => x"C0C0BFA4F8C0A480",
-27027 => x"C0C0BFA4F8C0A4F8",
-27026 => x"C0C0BFA4F8C0A482",
-27025 => x"C0C0BFA4F8C0A492",
-27024 => x"C0C0BFA4F8C0A499",
-27023 => x"C0C0BFA4F8C0A4B0",
-27022 => x"C0C0BFA4F8C0A4A4",
-27021 => x"C0C0BFA4F8C0A4F9",
-27020 => x"C0C0BFA4F8C0A4C0",
-27019 => x"C0C0BFA4F8C0F990",
-27018 => x"C0C0BFA4F8C0F980",
-27017 => x"C0C0BFA4F8C0F9F8",
-27016 => x"C0C0BFA4F8C0F982",
-27015 => x"C0C0BFA4F8C0F992",
-27014 => x"C0C0BFA4F8C0F999",
-27013 => x"C0C0BFA4F8C0F9B0",
-27012 => x"C0C0BFA4F8C0F9A4",
-27011 => x"C0C0BFA4F8C0F9F9",
-27010 => x"C0C0BFA4F8C0F9C0",
-27009 => x"C0C0BFA4F8C0C090",
-27008 => x"C0C0BFA4F8C0C080",
-27007 => x"C0C0BFA4F8C0C0F8",
-27006 => x"C0C0BFA4F8C0C082",
-27005 => x"C0C0BFA4F8C0C092",
-27004 => x"C0C0BFA4F8C0C099",
-27003 => x"C0C0BFA4F8C0C0B0",
-27002 => x"C0C0BFA4F8C0C0A4",
-27001 => x"C0C0BFA4F8C0C0F9",
-27000 => x"C0C0BFA4F8C0C0C0",
-26999 => x"C0C0BFA482909090",
-26998 => x"C0C0BFA482909080",
-26997 => x"C0C0BFA4829090F8",
-26996 => x"C0C0BFA482909082",
-26995 => x"C0C0BFA482909092",
-26994 => x"C0C0BFA482909099",
-26993 => x"C0C0BFA4829090B0",
-26992 => x"C0C0BFA4829090A4",
-26991 => x"C0C0BFA4829090F9",
-26990 => x"C0C0BFA4829090C0",
-26989 => x"C0C0BFA482908090",
-26988 => x"C0C0BFA482908080",
-26987 => x"C0C0BFA4829080F8",
-26986 => x"C0C0BFA482908082",
-26985 => x"C0C0BFA482908092",
-26984 => x"C0C0BFA482908099",
-26983 => x"C0C0BFA4829080B0",
-26982 => x"C0C0BFA4829080A4",
-26981 => x"C0C0BFA4829080F9",
-26980 => x"C0C0BFA4829080C0",
-26979 => x"C0C0BFA48290F890",
-26978 => x"C0C0BFA48290F880",
-26977 => x"C0C0BFA48290F8F8",
-26976 => x"C0C0BFA48290F882",
-26975 => x"C0C0BFA48290F892",
-26974 => x"C0C0BFA48290F899",
-26973 => x"C0C0BFA48290F8B0",
-26972 => x"C0C0BFA48290F8A4",
-26971 => x"C0C0BFA48290F8F9",
-26970 => x"C0C0BFA48290F8C0",
-26969 => x"C0C0BFA482908290",
-26968 => x"C0C0BFA482908280",
-26967 => x"C0C0BFA4829082F8",
-26966 => x"C0C0BFA482908282",
-26965 => x"C0C0BFA482908292",
-26964 => x"C0C0BFA482908299",
-26963 => x"C0C0BFA4829082B0",
-26962 => x"C0C0BFA4829082A4",
-26961 => x"C0C0BFA4829082F9",
-26960 => x"C0C0BFA4829082C0",
-26959 => x"C0C0BFA482909290",
-26958 => x"C0C0BFA482909280",
-26957 => x"C0C0BFA4829092F8",
-26956 => x"C0C0BFA482909282",
-26955 => x"C0C0BFA482909292",
-26954 => x"C0C0BFA482909299",
-26953 => x"C0C0BFA4829092B0",
-26952 => x"C0C0BFA4829092A4",
-26951 => x"C0C0BFA4829092F9",
-26950 => x"C0C0BFA4829092C0",
-26949 => x"C0C0BFA482909990",
-26948 => x"C0C0BFA482909980",
-26947 => x"C0C0BFA4829099F8",
-26946 => x"C0C0BFA482909982",
-26945 => x"C0C0BFA482909992",
-26944 => x"C0C0BFA482909999",
-26943 => x"C0C0BFA4829099B0",
-26942 => x"C0C0BFA4829099A4",
-26941 => x"C0C0BFA4829099F9",
-26940 => x"C0C0BFA4829099C0",
-26939 => x"C0C0BFA48290B090",
-26938 => x"C0C0BFA48290B080",
-26937 => x"C0C0BFA48290B0F8",
-26936 => x"C0C0BFA48290B082",
-26935 => x"C0C0BFA48290B092",
-26934 => x"C0C0BFA48290B099",
-26933 => x"C0C0BFA48290B0B0",
-26932 => x"C0C0BFA48290B0A4",
-26931 => x"C0C0BFA48290B0F9",
-26930 => x"C0C0BFA48290B0C0",
-26929 => x"C0C0BFA48290A490",
-26928 => x"C0C0BFA48290A480",
-26927 => x"C0C0BFA48290A4F8",
-26926 => x"C0C0BFA48290A482",
-26925 => x"C0C0BFA48290A492",
-26924 => x"C0C0BFA48290A499",
-26923 => x"C0C0BFA48290A4B0",
-26922 => x"C0C0BFA48290A4A4",
-26921 => x"C0C0BFA48290A4F9",
-26920 => x"C0C0BFA48290A4C0",
-26919 => x"C0C0BFA48290F990",
-26918 => x"C0C0BFA48290F980",
-26917 => x"C0C0BFA48290F9F8",
-26916 => x"C0C0BFA48290F982",
-26915 => x"C0C0BFA48290F992",
-26914 => x"C0C0BFA48290F999",
-26913 => x"C0C0BFA48290F9B0",
-26912 => x"C0C0BFA48290F9A4",
-26911 => x"C0C0BFA48290F9F9",
-26910 => x"C0C0BFA48290F9C0",
-26909 => x"C0C0BFA48290C090",
-26908 => x"C0C0BFA48290C080",
-26907 => x"C0C0BFA48290C0F8",
-26906 => x"C0C0BFA48290C082",
-26905 => x"C0C0BFA48290C092",
-26904 => x"C0C0BFA48290C099",
-26903 => x"C0C0BFA48290C0B0",
-26902 => x"C0C0BFA48290C0A4",
-26901 => x"C0C0BFA48290C0F9",
-26900 => x"C0C0BFA48290C0C0",
-26899 => x"C0C0BFA482809090",
-26898 => x"C0C0BFA482809080",
-26897 => x"C0C0BFA4828090F8",
-26896 => x"C0C0BFA482809082",
-26895 => x"C0C0BFA482809092",
-26894 => x"C0C0BFA482809099",
-26893 => x"C0C0BFA4828090B0",
-26892 => x"C0C0BFA4828090A4",
-26891 => x"C0C0BFA4828090F9",
-26890 => x"C0C0BFA4828090C0",
-26889 => x"C0C0BFA482808090",
-26888 => x"C0C0BFA482808080",
-26887 => x"C0C0BFA4828080F8",
-26886 => x"C0C0BFA482808082",
-26885 => x"C0C0BFA482808092",
-26884 => x"C0C0BFA482808099",
-26883 => x"C0C0BFA4828080B0",
-26882 => x"C0C0BFA4828080A4",
-26881 => x"C0C0BFA4828080F9",
-26880 => x"C0C0BFA4828080C0",
-26879 => x"C0C0BFA48280F890",
-26878 => x"C0C0BFA48280F880",
-26877 => x"C0C0BFA48280F8F8",
-26876 => x"C0C0BFA48280F882",
-26875 => x"C0C0BFA48280F892",
-26874 => x"C0C0BFA48280F899",
-26873 => x"C0C0BFA48280F8B0",
-26872 => x"C0C0BFA48280F8A4",
-26871 => x"C0C0BFA48280F8F9",
-26870 => x"C0C0BFA48280F8C0",
-26869 => x"C0C0BFA482808290",
-26868 => x"C0C0BFA482808280",
-26867 => x"C0C0BFA4828082F8",
-26866 => x"C0C0BFA482808282",
-26865 => x"C0C0BFA482808292",
-26864 => x"C0C0BFA482808299",
-26863 => x"C0C0BFA4828082B0",
-26862 => x"C0C0BFA4828082A4",
-26861 => x"C0C0BFA4828082F9",
-26860 => x"C0C0BFA4828082C0",
-26859 => x"C0C0BFA482809290",
-26858 => x"C0C0BFA482809280",
-26857 => x"C0C0BFA4828092F8",
-26856 => x"C0C0BFA482809282",
-26855 => x"C0C0BFA482809292",
-26854 => x"C0C0BFA482809299",
-26853 => x"C0C0BFA4828092B0",
-26852 => x"C0C0BFA4828092A4",
-26851 => x"C0C0BFA4828092F9",
-26850 => x"C0C0BFA4828092C0",
-26849 => x"C0C0BFA482809990",
-26848 => x"C0C0BFA482809980",
-26847 => x"C0C0BFA4828099F8",
-26846 => x"C0C0BFA482809982",
-26845 => x"C0C0BFA482809992",
-26844 => x"C0C0BFA482809999",
-26843 => x"C0C0BFA4828099B0",
-26842 => x"C0C0BFA4828099A4",
-26841 => x"C0C0BFA4828099F9",
-26840 => x"C0C0BFA4828099C0",
-26839 => x"C0C0BFA48280B090",
-26838 => x"C0C0BFA48280B080",
-26837 => x"C0C0BFA48280B0F8",
-26836 => x"C0C0BFA48280B082",
-26835 => x"C0C0BFA48280B092",
-26834 => x"C0C0BFA48280B099",
-26833 => x"C0C0BFA48280B0B0",
-26832 => x"C0C0BFA48280B0A4",
-26831 => x"C0C0BFA48280B0F9",
-26830 => x"C0C0BFA48280B0C0",
-26829 => x"C0C0BFA48280A490",
-26828 => x"C0C0BFA48280A480",
-26827 => x"C0C0BFA48280A4F8",
-26826 => x"C0C0BFA48280A482",
-26825 => x"C0C0BFA48280A492",
-26824 => x"C0C0BFA48280A499",
-26823 => x"C0C0BFA48280A4B0",
-26822 => x"C0C0BFA48280A4A4",
-26821 => x"C0C0BFA48280A4F9",
-26820 => x"C0C0BFA48280A4C0",
-26819 => x"C0C0BFA48280F990",
-26818 => x"C0C0BFA48280F980",
-26817 => x"C0C0BFA48280F9F8",
-26816 => x"C0C0BFA48280F982",
-26815 => x"C0C0BFA48280F992",
-26814 => x"C0C0BFA48280F999",
-26813 => x"C0C0BFA48280F9B0",
-26812 => x"C0C0BFA48280F9A4",
-26811 => x"C0C0BFA48280F9F9",
-26810 => x"C0C0BFA48280F9C0",
-26809 => x"C0C0BFA48280C090",
-26808 => x"C0C0BFA48280C080",
-26807 => x"C0C0BFA48280C0F8",
-26806 => x"C0C0BFA48280C082",
-26805 => x"C0C0BFA48280C092",
-26804 => x"C0C0BFA48280C099",
-26803 => x"C0C0BFA48280C0B0",
-26802 => x"C0C0BFA48280C0A4",
-26801 => x"C0C0BFA48280C0F9",
-26800 => x"C0C0BFA48280C0C0",
-26799 => x"C0C0BFA482F89090",
-26798 => x"C0C0BFA482F89080",
-26797 => x"C0C0BFA482F890F8",
-26796 => x"C0C0BFA482F89082",
-26795 => x"C0C0BFA482F89092",
-26794 => x"C0C0BFA482F89099",
-26793 => x"C0C0BFA482F890B0",
-26792 => x"C0C0BFA482F890A4",
-26791 => x"C0C0BFA482F890F9",
-26790 => x"C0C0BFA482F890C0",
-26789 => x"C0C0BFA482F88090",
-26788 => x"C0C0BFA482F88080",
-26787 => x"C0C0BFA482F880F8",
-26786 => x"C0C0BFA482F88082",
-26785 => x"C0C0BFA482F88092",
-26784 => x"C0C0BFA482F88099",
-26783 => x"C0C0BFA482F880B0",
-26782 => x"C0C0BFA482F880A4",
-26781 => x"C0C0BFA482F880F9",
-26780 => x"C0C0BFA482F880C0",
-26779 => x"C0C0BFA482F8F890",
-26778 => x"C0C0BFA482F8F880",
-26777 => x"C0C0BFA482F8F8F8",
-26776 => x"C0C0BFA482F8F882",
-26775 => x"C0C0BFA482F8F892",
-26774 => x"C0C0BFA482F8F899",
-26773 => x"C0C0BFA482F8F8B0",
-26772 => x"C0C0BFA482F8F8A4",
-26771 => x"C0C0BFA482F8F8F9",
-26770 => x"C0C0BFA482F8F8C0",
-26769 => x"C0C0BFA482F88290",
-26768 => x"C0C0BFA482F88280",
-26767 => x"C0C0BFA482F882F8",
-26766 => x"C0C0BFA482F88282",
-26765 => x"C0C0BFA482F88292",
-26764 => x"C0C0BFA482F88299",
-26763 => x"C0C0BFA482F882B0",
-26762 => x"C0C0BFA482F882A4",
-26761 => x"C0C0BFA482F882F9",
-26760 => x"C0C0BFA482F882C0",
-26759 => x"C0C0BFA482F89290",
-26758 => x"C0C0BFA482F89280",
-26757 => x"C0C0BFA482F892F8",
-26756 => x"C0C0BFA482F89282",
-26755 => x"C0C0BFA482F89292",
-26754 => x"C0C0BFA482F89299",
-26753 => x"C0C0BFA482F892B0",
-26752 => x"C0C0BFA482F892A4",
-26751 => x"C0C0BFA482F892F9",
-26750 => x"C0C0BFA482F892C0",
-26749 => x"C0C0BFA482F89990",
-26748 => x"C0C0BFA482F89980",
-26747 => x"C0C0BFA482F899F8",
-26746 => x"C0C0BFA482F89982",
-26745 => x"C0C0BFA482F89992",
-26744 => x"C0C0BFA482F89999",
-26743 => x"C0C0BFA482F899B0",
-26742 => x"C0C0BFA482F899A4",
-26741 => x"C0C0BFA482F899F9",
-26740 => x"C0C0BFA482F899C0",
-26739 => x"C0C0BFA482F8B090",
-26738 => x"C0C0BFA482F8B080",
-26737 => x"C0C0BFA482F8B0F8",
-26736 => x"C0C0BFA482F8B082",
-26735 => x"C0C0BFA482F8B092",
-26734 => x"C0C0BFA482F8B099",
-26733 => x"C0C0BFA482F8B0B0",
-26732 => x"C0C0BFA482F8B0A4",
-26731 => x"C0C0BFA482F8B0F9",
-26730 => x"C0C0BFA482F8B0C0",
-26729 => x"C0C0BFA482F8A490",
-26728 => x"C0C0BFA482F8A480",
-26727 => x"C0C0BFA482F8A4F8",
-26726 => x"C0C0BFA482F8A482",
-26725 => x"C0C0BFA482F8A492",
-26724 => x"C0C0BFA482F8A499",
-26723 => x"C0C0BFA482F8A4B0",
-26722 => x"C0C0BFA482F8A4A4",
-26721 => x"C0C0BFA482F8A4F9",
-26720 => x"C0C0BFA482F8A4C0",
-26719 => x"C0C0BFA482F8F990",
-26718 => x"C0C0BFA482F8F980",
-26717 => x"C0C0BFA482F8F9F8",
-26716 => x"C0C0BFA482F8F982",
-26715 => x"C0C0BFA482F8F992",
-26714 => x"C0C0BFA482F8F999",
-26713 => x"C0C0BFA482F8F9B0",
-26712 => x"C0C0BFA482F8F9A4",
-26711 => x"C0C0BFA482F8F9F9",
-26710 => x"C0C0BFA482F8F9C0",
-26709 => x"C0C0BFA482F8C090",
-26708 => x"C0C0BFA482F8C080",
-26707 => x"C0C0BFA482F8C0F8",
-26706 => x"C0C0BFA482F8C082",
-26705 => x"C0C0BFA482F8C092",
-26704 => x"C0C0BFA482F8C099",
-26703 => x"C0C0BFA482F8C0B0",
-26702 => x"C0C0BFA482F8C0A4",
-26701 => x"C0C0BFA482F8C0F9",
-26700 => x"C0C0BFA482F8C0C0",
-26699 => x"C0C0BFA482829090",
-26698 => x"C0C0BFA482829080",
-26697 => x"C0C0BFA4828290F8",
-26696 => x"C0C0BFA482829082",
-26695 => x"C0C0BFA482829092",
-26694 => x"C0C0BFA482829099",
-26693 => x"C0C0BFA4828290B0",
-26692 => x"C0C0BFA4828290A4",
-26691 => x"C0C0BFA4828290F9",
-26690 => x"C0C0BFA4828290C0",
-26689 => x"C0C0BFA482828090",
-26688 => x"C0C0BFA482828080",
-26687 => x"C0C0BFA4828280F8",
-26686 => x"C0C0BFA482828082",
-26685 => x"C0C0BFA482828092",
-26684 => x"C0C0BFA482828099",
-26683 => x"C0C0BFA4828280B0",
-26682 => x"C0C0BFA4828280A4",
-26681 => x"C0C0BFA4828280F9",
-26680 => x"C0C0BFA4828280C0",
-26679 => x"C0C0BFA48282F890",
-26678 => x"C0C0BFA48282F880",
-26677 => x"C0C0BFA48282F8F8",
-26676 => x"C0C0BFA48282F882",
-26675 => x"C0C0BFA48282F892",
-26674 => x"C0C0BFA48282F899",
-26673 => x"C0C0BFA48282F8B0",
-26672 => x"C0C0BFA48282F8A4",
-26671 => x"C0C0BFA48282F8F9",
-26670 => x"C0C0BFA48282F8C0",
-26669 => x"C0C0BFA482828290",
-26668 => x"C0C0BFA482828280",
-26667 => x"C0C0BFA4828282F8",
-26666 => x"C0C0BFA482828282",
-26665 => x"C0C0BFA482828292",
-26664 => x"C0C0BFA482828299",
-26663 => x"C0C0BFA4828282B0",
-26662 => x"C0C0BFA4828282A4",
-26661 => x"C0C0BFA4828282F9",
-26660 => x"C0C0BFA4828282C0",
-26659 => x"C0C0BFA482829290",
-26658 => x"C0C0BFA482829280",
-26657 => x"C0C0BFA4828292F8",
-26656 => x"C0C0BFA482829282",
-26655 => x"C0C0BFA482829292",
-26654 => x"C0C0BFA482829299",
-26653 => x"C0C0BFA4828292B0",
-26652 => x"C0C0BFA4828292A4",
-26651 => x"C0C0BFA4828292F9",
-26650 => x"C0C0BFA4828292C0",
-26649 => x"C0C0BFA482829990",
-26648 => x"C0C0BFA482829980",
-26647 => x"C0C0BFA4828299F8",
-26646 => x"C0C0BFA482829982",
-26645 => x"C0C0BFA482829992",
-26644 => x"C0C0BFA482829999",
-26643 => x"C0C0BFA4828299B0",
-26642 => x"C0C0BFA4828299A4",
-26641 => x"C0C0BFA4828299F9",
-26640 => x"C0C0BFA4828299C0",
-26639 => x"C0C0BFA48282B090",
-26638 => x"C0C0BFA48282B080",
-26637 => x"C0C0BFA48282B0F8",
-26636 => x"C0C0BFA48282B082",
-26635 => x"C0C0BFA48282B092",
-26634 => x"C0C0BFA48282B099",
-26633 => x"C0C0BFA48282B0B0",
-26632 => x"C0C0BFA48282B0A4",
-26631 => x"C0C0BFA48282B0F9",
-26630 => x"C0C0BFA48282B0C0",
-26629 => x"C0C0BFA48282A490",
-26628 => x"C0C0BFA48282A480",
-26627 => x"C0C0BFA48282A4F8",
-26626 => x"C0C0BFA48282A482",
-26625 => x"C0C0BFA48282A492",
-26624 => x"C0C0BFA48282A499",
-26623 => x"C0C0BFA48282A4B0",
-26622 => x"C0C0BFA48282A4A4",
-26621 => x"C0C0BFA48282A4F9",
-26620 => x"C0C0BFA48282A4C0",
-26619 => x"C0C0BFA48282F990",
-26618 => x"C0C0BFA48282F980",
-26617 => x"C0C0BFA48282F9F8",
-26616 => x"C0C0BFA48282F982",
-26615 => x"C0C0BFA48282F992",
-26614 => x"C0C0BFA48282F999",
-26613 => x"C0C0BFA48282F9B0",
-26612 => x"C0C0BFA48282F9A4",
-26611 => x"C0C0BFA48282F9F9",
-26610 => x"C0C0BFA48282F9C0",
-26609 => x"C0C0BFA48282C090",
-26608 => x"C0C0BFA48282C080",
-26607 => x"C0C0BFA48282C0F8",
-26606 => x"C0C0BFA48282C082",
-26605 => x"C0C0BFA48282C092",
-26604 => x"C0C0BFA48282C099",
-26603 => x"C0C0BFA48282C0B0",
-26602 => x"C0C0BFA48282C0A4",
-26601 => x"C0C0BFA48282C0F9",
-26600 => x"C0C0BFA48282C0C0",
-26599 => x"C0C0BFA482929090",
-26598 => x"C0C0BFA482929080",
-26597 => x"C0C0BFA4829290F8",
-26596 => x"C0C0BFA482929082",
-26595 => x"C0C0BFA482929092",
-26594 => x"C0C0BFA482929099",
-26593 => x"C0C0BFA4829290B0",
-26592 => x"C0C0BFA4829290A4",
-26591 => x"C0C0BFA4829290F9",
-26590 => x"C0C0BFA4829290C0",
-26589 => x"C0C0BFA482928090",
-26588 => x"C0C0BFA482928080",
-26587 => x"C0C0BFA4829280F8",
-26586 => x"C0C0BFA482928082",
-26585 => x"C0C0BFA482928092",
-26584 => x"C0C0BFA482928099",
-26583 => x"C0C0BFA4829280B0",
-26582 => x"C0C0BFA4829280A4",
-26581 => x"C0C0BFA4829280F9",
-26580 => x"C0C0BFA4829280C0",
-26579 => x"C0C0BFA48292F890",
-26578 => x"C0C0BFA48292F880",
-26577 => x"C0C0BFA48292F8F8",
-26576 => x"C0C0BFA48292F882",
-26575 => x"C0C0BFA48292F892",
-26574 => x"C0C0BFA48292F899",
-26573 => x"C0C0BFA48292F8B0",
-26572 => x"C0C0BFA48292F8A4",
-26571 => x"C0C0BFA48292F8F9",
-26570 => x"C0C0BFA48292F8C0",
-26569 => x"C0C0BFA482928290",
-26568 => x"C0C0BFA482928280",
-26567 => x"C0C0BFA4829282F8",
-26566 => x"C0C0BFA482928282",
-26565 => x"C0C0BFA482928292",
-26564 => x"C0C0BFA482928299",
-26563 => x"C0C0BFA4829282B0",
-26562 => x"C0C0BFA4829282A4",
-26561 => x"C0C0BFA4829282F9",
-26560 => x"C0C0BFA4829282C0",
-26559 => x"C0C0BFA482929290",
-26558 => x"C0C0BFA482929280",
-26557 => x"C0C0BFA4829292F8",
-26556 => x"C0C0BFA482929282",
-26555 => x"C0C0BFA482929292",
-26554 => x"C0C0BFA482929299",
-26553 => x"C0C0BFA4829292B0",
-26552 => x"C0C0BFA4829292A4",
-26551 => x"C0C0BFA4829292F9",
-26550 => x"C0C0BFA4829292C0",
-26549 => x"C0C0BFA482929990",
-26548 => x"C0C0BFA482929980",
-26547 => x"C0C0BFA4829299F8",
-26546 => x"C0C0BFA482929982",
-26545 => x"C0C0BFA482929992",
-26544 => x"C0C0BFA482929999",
-26543 => x"C0C0BFA4829299B0",
-26542 => x"C0C0BFA4829299A4",
-26541 => x"C0C0BFA4829299F9",
-26540 => x"C0C0BFA4829299C0",
-26539 => x"C0C0BFA48292B090",
-26538 => x"C0C0BFA48292B080",
-26537 => x"C0C0BFA48292B0F8",
-26536 => x"C0C0BFA48292B082",
-26535 => x"C0C0BFA48292B092",
-26534 => x"C0C0BFA48292B099",
-26533 => x"C0C0BFA48292B0B0",
-26532 => x"C0C0BFA48292B0A4",
-26531 => x"C0C0BFA48292B0F9",
-26530 => x"C0C0BFA48292B0C0",
-26529 => x"C0C0BFA48292A490",
-26528 => x"C0C0BFA48292A480",
-26527 => x"C0C0BFA48292A4F8",
-26526 => x"C0C0BFA48292A482",
-26525 => x"C0C0BFA48292A492",
-26524 => x"C0C0BFA48292A499",
-26523 => x"C0C0BFA48292A4B0",
-26522 => x"C0C0BFA48292A4A4",
-26521 => x"C0C0BFA48292A4F9",
-26520 => x"C0C0BFA48292A4C0",
-26519 => x"C0C0BFA48292F990",
-26518 => x"C0C0BFA48292F980",
-26517 => x"C0C0BFA48292F9F8",
-26516 => x"C0C0BFA48292F982",
-26515 => x"C0C0BFA48292F992",
-26514 => x"C0C0BFA48292F999",
-26513 => x"C0C0BFA48292F9B0",
-26512 => x"C0C0BFA48292F9A4",
-26511 => x"C0C0BFA48292F9F9",
-26510 => x"C0C0BFA48292F9C0",
-26509 => x"C0C0BFA48292C090",
-26508 => x"C0C0BFA48292C080",
-26507 => x"C0C0BFA48292C0F8",
-26506 => x"C0C0BFA48292C082",
-26505 => x"C0C0BFA48292C092",
-26504 => x"C0C0BFA48292C099",
-26503 => x"C0C0BFA48292C0B0",
-26502 => x"C0C0BFA48292C0A4",
-26501 => x"C0C0BFA48292C0F9",
-26500 => x"C0C0BFA48292C0C0",
-26499 => x"C0C0BFA482999090",
-26498 => x"C0C0BFA482999080",
-26497 => x"C0C0BFA4829990F8",
-26496 => x"C0C0BFA482999082",
-26495 => x"C0C0BFA482999092",
-26494 => x"C0C0BFA482999099",
-26493 => x"C0C0BFA4829990B0",
-26492 => x"C0C0BFA4829990A4",
-26491 => x"C0C0BFA4829990F9",
-26490 => x"C0C0BFA4829990C0",
-26489 => x"C0C0BFA482998090",
-26488 => x"C0C0BFA482998080",
-26487 => x"C0C0BFA4829980F8",
-26486 => x"C0C0BFA482998082",
-26485 => x"C0C0BFA482998092",
-26484 => x"C0C0BFA482998099",
-26483 => x"C0C0BFA4829980B0",
-26482 => x"C0C0BFA4829980A4",
-26481 => x"C0C0BFA4829980F9",
-26480 => x"C0C0BFA4829980C0",
-26479 => x"C0C0BFA48299F890",
-26478 => x"C0C0BFA48299F880",
-26477 => x"C0C0BFA48299F8F8",
-26476 => x"C0C0BFA48299F882",
-26475 => x"C0C0BFA48299F892",
-26474 => x"C0C0BFA48299F899",
-26473 => x"C0C0BFA48299F8B0",
-26472 => x"C0C0BFA48299F8A4",
-26471 => x"C0C0BFA48299F8F9",
-26470 => x"C0C0BFA48299F8C0",
-26469 => x"C0C0BFA482998290",
-26468 => x"C0C0BFA482998280",
-26467 => x"C0C0BFA4829982F8",
-26466 => x"C0C0BFA482998282",
-26465 => x"C0C0BFA482998292",
-26464 => x"C0C0BFA482998299",
-26463 => x"C0C0BFA4829982B0",
-26462 => x"C0C0BFA4829982A4",
-26461 => x"C0C0BFA4829982F9",
-26460 => x"C0C0BFA4829982C0",
-26459 => x"C0C0BFA482999290",
-26458 => x"C0C0BFA482999280",
-26457 => x"C0C0BFA4829992F8",
-26456 => x"C0C0BFA482999282",
-26455 => x"C0C0BFA482999292",
-26454 => x"C0C0BFA482999299",
-26453 => x"C0C0BFA4829992B0",
-26452 => x"C0C0BFA4829992A4",
-26451 => x"C0C0BFA4829992F9",
-26450 => x"C0C0BFA4829992C0",
-26449 => x"C0C0BFA482999990",
-26448 => x"C0C0BFA482999980",
-26447 => x"C0C0BFA4829999F8",
-26446 => x"C0C0BFA482999982",
-26445 => x"C0C0BFA482999992",
-26444 => x"C0C0BFA482999999",
-26443 => x"C0C0BFA4829999B0",
-26442 => x"C0C0BFA4829999A4",
-26441 => x"C0C0BFA4829999F9",
-26440 => x"C0C0BFA4829999C0",
-26439 => x"C0C0BFA48299B090",
-26438 => x"C0C0BFA48299B080",
-26437 => x"C0C0BFA48299B0F8",
-26436 => x"C0C0BFA48299B082",
-26435 => x"C0C0BFA48299B092",
-26434 => x"C0C0BFA48299B099",
-26433 => x"C0C0BFA48299B0B0",
-26432 => x"C0C0BFA48299B0A4",
-26431 => x"C0C0BFA48299B0F9",
-26430 => x"C0C0BFA48299B0C0",
-26429 => x"C0C0BFA48299A490",
-26428 => x"C0C0BFA48299A480",
-26427 => x"C0C0BFA48299A4F8",
-26426 => x"C0C0BFA48299A482",
-26425 => x"C0C0BFA48299A492",
-26424 => x"C0C0BFA48299A499",
-26423 => x"C0C0BFA48299A4B0",
-26422 => x"C0C0BFA48299A4A4",
-26421 => x"C0C0BFA48299A4F9",
-26420 => x"C0C0BFA48299A4C0",
-26419 => x"C0C0BFA48299F990",
-26418 => x"C0C0BFA48299F980",
-26417 => x"C0C0BFA48299F9F8",
-26416 => x"C0C0BFA48299F982",
-26415 => x"C0C0BFA48299F992",
-26414 => x"C0C0BFA48299F999",
-26413 => x"C0C0BFA48299F9B0",
-26412 => x"C0C0BFA48299F9A4",
-26411 => x"C0C0BFA48299F9F9",
-26410 => x"C0C0BFA48299F9C0",
-26409 => x"C0C0BFA48299C090",
-26408 => x"C0C0BFA48299C080",
-26407 => x"C0C0BFA48299C0F8",
-26406 => x"C0C0BFA48299C082",
-26405 => x"C0C0BFA48299C092",
-26404 => x"C0C0BFA48299C099",
-26403 => x"C0C0BFA48299C0B0",
-26402 => x"C0C0BFA48299C0A4",
-26401 => x"C0C0BFA48299C0F9",
-26400 => x"C0C0BFA48299C0C0",
-26399 => x"C0C0BFA482B09090",
-26398 => x"C0C0BFA482B09080",
-26397 => x"C0C0BFA482B090F8",
-26396 => x"C0C0BFA482B09082",
-26395 => x"C0C0BFA482B09092",
-26394 => x"C0C0BFA482B09099",
-26393 => x"C0C0BFA482B090B0",
-26392 => x"C0C0BFA482B090A4",
-26391 => x"C0C0BFA482B090F9",
-26390 => x"C0C0BFA482B090C0",
-26389 => x"C0C0BFA482B08090",
-26388 => x"C0C0BFA482B08080",
-26387 => x"C0C0BFA482B080F8",
-26386 => x"C0C0BFA482B08082",
-26385 => x"C0C0BFA482B08092",
-26384 => x"C0C0BFA482B08099",
-26383 => x"C0C0BFA482B080B0",
-26382 => x"C0C0BFA482B080A4",
-26381 => x"C0C0BFA482B080F9",
-26380 => x"C0C0BFA482B080C0",
-26379 => x"C0C0BFA482B0F890",
-26378 => x"C0C0BFA482B0F880",
-26377 => x"C0C0BFA482B0F8F8",
-26376 => x"C0C0BFA482B0F882",
-26375 => x"C0C0BFA482B0F892",
-26374 => x"C0C0BFA482B0F899",
-26373 => x"C0C0BFA482B0F8B0",
-26372 => x"C0C0BFA482B0F8A4",
-26371 => x"C0C0BFA482B0F8F9",
-26370 => x"C0C0BFA482B0F8C0",
-26369 => x"C0C0BFA482B08290",
-26368 => x"C0C0BFA482B08280",
-26367 => x"C0C0BFA482B082F8",
-26366 => x"C0C0BFA482B08282",
-26365 => x"C0C0BFA482B08292",
-26364 => x"C0C0BFA482B08299",
-26363 => x"C0C0BFA482B082B0",
-26362 => x"C0C0BFA482B082A4",
-26361 => x"C0C0BFA482B082F9",
-26360 => x"C0C0BFA482B082C0",
-26359 => x"C0C0BFA482B09290",
-26358 => x"C0C0BFA482B09280",
-26357 => x"C0C0BFA482B092F8",
-26356 => x"C0C0BFA482B09282",
-26355 => x"C0C0BFA482B09292",
-26354 => x"C0C0BFA482B09299",
-26353 => x"C0C0BFA482B092B0",
-26352 => x"C0C0BFA482B092A4",
-26351 => x"C0C0BFA482B092F9",
-26350 => x"C0C0BFA482B092C0",
-26349 => x"C0C0BFA482B09990",
-26348 => x"C0C0BFA482B09980",
-26347 => x"C0C0BFA482B099F8",
-26346 => x"C0C0BFA482B09982",
-26345 => x"C0C0BFA482B09992",
-26344 => x"C0C0BFA482B09999",
-26343 => x"C0C0BFA482B099B0",
-26342 => x"C0C0BFA482B099A4",
-26341 => x"C0C0BFA482B099F9",
-26340 => x"C0C0BFA482B099C0",
-26339 => x"C0C0BFA482B0B090",
-26338 => x"C0C0BFA482B0B080",
-26337 => x"C0C0BFA482B0B0F8",
-26336 => x"C0C0BFA482B0B082",
-26335 => x"C0C0BFA482B0B092",
-26334 => x"C0C0BFA482B0B099",
-26333 => x"C0C0BFA482B0B0B0",
-26332 => x"C0C0BFA482B0B0A4",
-26331 => x"C0C0BFA482B0B0F9",
-26330 => x"C0C0BFA482B0B0C0",
-26329 => x"C0C0BFA482B0A490",
-26328 => x"C0C0BFA482B0A480",
-26327 => x"C0C0BFA482B0A4F8",
-26326 => x"C0C0BFA482B0A482",
-26325 => x"C0C0BFA482B0A492",
-26324 => x"C0C0BFA482B0A499",
-26323 => x"C0C0BFA482B0A4B0",
-26322 => x"C0C0BFA482B0A4A4",
-26321 => x"C0C0BFA482B0A4F9",
-26320 => x"C0C0BFA482B0A4C0",
-26319 => x"C0C0BFA482B0F990",
-26318 => x"C0C0BFA482B0F980",
-26317 => x"C0C0BFA482B0F9F8",
-26316 => x"C0C0BFA482B0F982",
-26315 => x"C0C0BFA482B0F992",
-26314 => x"C0C0BFA482B0F999",
-26313 => x"C0C0BFA482B0F9B0",
-26312 => x"C0C0BFA482B0F9A4",
-26311 => x"C0C0BFA482B0F9F9",
-26310 => x"C0C0BFA482B0F9C0",
-26309 => x"C0C0BFA482B0C090",
-26308 => x"C0C0BFA482B0C080",
-26307 => x"C0C0BFA482B0C0F8",
-26306 => x"C0C0BFA482B0C082",
-26305 => x"C0C0BFA482B0C092",
-26304 => x"C0C0BFA482B0C099",
-26303 => x"C0C0BFA482B0C0B0",
-26302 => x"C0C0BFA482B0C0A4",
-26301 => x"C0C0BFA482B0C0F9",
-26300 => x"C0C0BFA482B0C0C0",
-26299 => x"C0C0BFA482A49090",
-26298 => x"C0C0BFA482A49080",
-26297 => x"C0C0BFA482A490F8",
-26296 => x"C0C0BFA482A49082",
-26295 => x"C0C0BFA482A49092",
-26294 => x"C0C0BFA482A49099",
-26293 => x"C0C0BFA482A490B0",
-26292 => x"C0C0BFA482A490A4",
-26291 => x"C0C0BFA482A490F9",
-26290 => x"C0C0BFA482A490C0",
-26289 => x"C0C0BFA482A48090",
-26288 => x"C0C0BFA482A48080",
-26287 => x"C0C0BFA482A480F8",
-26286 => x"C0C0BFA482A48082",
-26285 => x"C0C0BFA482A48092",
-26284 => x"C0C0BFA482A48099",
-26283 => x"C0C0BFA482A480B0",
-26282 => x"C0C0BFA482A480A4",
-26281 => x"C0C0BFA482A480F9",
-26280 => x"C0C0BFA482A480C0",
-26279 => x"C0C0BFA482A4F890",
-26278 => x"C0C0BFA482A4F880",
-26277 => x"C0C0BFA482A4F8F8",
-26276 => x"C0C0BFA482A4F882",
-26275 => x"C0C0BFA482A4F892",
-26274 => x"C0C0BFA482A4F899",
-26273 => x"C0C0BFA482A4F8B0",
-26272 => x"C0C0BFA482A4F8A4",
-26271 => x"C0C0BFA482A4F8F9",
-26270 => x"C0C0BFA482A4F8C0",
-26269 => x"C0C0BFA482A48290",
-26268 => x"C0C0BFA482A48280",
-26267 => x"C0C0BFA482A482F8",
-26266 => x"C0C0BFA482A48282",
-26265 => x"C0C0BFA482A48292",
-26264 => x"C0C0BFA482A48299",
-26263 => x"C0C0BFA482A482B0",
-26262 => x"C0C0BFA482A482A4",
-26261 => x"C0C0BFA482A482F9",
-26260 => x"C0C0BFA482A482C0",
-26259 => x"C0C0BFA482A49290",
-26258 => x"C0C0BFA482A49280",
-26257 => x"C0C0BFA482A492F8",
-26256 => x"C0C0BFA482A49282",
-26255 => x"C0C0BFA482A49292",
-26254 => x"C0C0BFA482A49299",
-26253 => x"C0C0BFA482A492B0",
-26252 => x"C0C0BFA482A492A4",
-26251 => x"C0C0BFA482A492F9",
-26250 => x"C0C0BFA482A492C0",
-26249 => x"C0C0BFA482A49990",
-26248 => x"C0C0BFA482A49980",
-26247 => x"C0C0BFA482A499F8",
-26246 => x"C0C0BFA482A49982",
-26245 => x"C0C0BFA482A49992",
-26244 => x"C0C0BFA482A49999",
-26243 => x"C0C0BFA482A499B0",
-26242 => x"C0C0BFA482A499A4",
-26241 => x"C0C0BFA482A499F9",
-26240 => x"C0C0BFA482A499C0",
-26239 => x"C0C0BFA482A4B090",
-26238 => x"C0C0BFA482A4B080",
-26237 => x"C0C0BFA482A4B0F8",
-26236 => x"C0C0BFA482A4B082",
-26235 => x"C0C0BFA482A4B092",
-26234 => x"C0C0BFA482A4B099",
-26233 => x"C0C0BFA482A4B0B0",
-26232 => x"C0C0BFA482A4B0A4",
-26231 => x"C0C0BFA482A4B0F9",
-26230 => x"C0C0BFA482A4B0C0",
-26229 => x"C0C0BFA482A4A490",
-26228 => x"C0C0BFA482A4A480",
-26227 => x"C0C0BFA482A4A4F8",
-26226 => x"C0C0BFA482A4A482",
-26225 => x"C0C0BFA482A4A492",
-26224 => x"C0C0BFA482A4A499",
-26223 => x"C0C0BFA482A4A4B0",
-26222 => x"C0C0BFA482A4A4A4",
-26221 => x"C0C0BFA482A4A4F9",
-26220 => x"C0C0BFA482A4A4C0",
-26219 => x"C0C0BFA482A4F990",
-26218 => x"C0C0BFA482A4F980",
-26217 => x"C0C0BFA482A4F9F8",
-26216 => x"C0C0BFA482A4F982",
-26215 => x"C0C0BFA482A4F992",
-26214 => x"C0C0BFA482A4F999",
-26213 => x"C0C0BFA482A4F9B0",
-26212 => x"C0C0BFA482A4F9A4",
-26211 => x"C0C0BFA482A4F9F9",
-26210 => x"C0C0BFA482A4F9C0",
-26209 => x"C0C0BFA482A4C090",
-26208 => x"C0C0BFA482A4C080",
-26207 => x"C0C0BFA482A4C0F8",
-26206 => x"C0C0BFA482A4C082",
-26205 => x"C0C0BFA482A4C092",
-26204 => x"C0C0BFA482A4C099",
-26203 => x"C0C0BFA482A4C0B0",
-26202 => x"C0C0BFA482A4C0A4",
-26201 => x"C0C0BFA482A4C0F9",
-26200 => x"C0C0BFA482A4C0C0",
-26199 => x"C0C0BFA482F99090",
-26198 => x"C0C0BFA482F99080",
-26197 => x"C0C0BFA482F990F8",
-26196 => x"C0C0BFA482F99082",
-26195 => x"C0C0BFA482F99092",
-26194 => x"C0C0BFA482F99099",
-26193 => x"C0C0BFA482F990B0",
-26192 => x"C0C0BFA482F990A4",
-26191 => x"C0C0BFA482F990F9",
-26190 => x"C0C0BFA482F990C0",
-26189 => x"C0C0BFA482F98090",
-26188 => x"C0C0BFA482F98080",
-26187 => x"C0C0BFA482F980F8",
-26186 => x"C0C0BFA482F98082",
-26185 => x"C0C0BFA482F98092",
-26184 => x"C0C0BFA482F98099",
-26183 => x"C0C0BFA482F980B0",
-26182 => x"C0C0BFA482F980A4",
-26181 => x"C0C0BFA482F980F9",
-26180 => x"C0C0BFA482F980C0",
-26179 => x"C0C0BFA482F9F890",
-26178 => x"C0C0BFA482F9F880",
-26177 => x"C0C0BFA482F9F8F8",
-26176 => x"C0C0BFA482F9F882",
-26175 => x"C0C0BFA482F9F892",
-26174 => x"C0C0BFA482F9F899",
-26173 => x"C0C0BFA482F9F8B0",
-26172 => x"C0C0BFA482F9F8A4",
-26171 => x"C0C0BFA482F9F8F9",
-26170 => x"C0C0BFA482F9F8C0",
-26169 => x"C0C0BFA482F98290",
-26168 => x"C0C0BFA482F98280",
-26167 => x"C0C0BFA482F982F8",
-26166 => x"C0C0BFA482F98282",
-26165 => x"C0C0BFA482F98292",
-26164 => x"C0C0BFA482F98299",
-26163 => x"C0C0BFA482F982B0",
-26162 => x"C0C0BFA482F982A4",
-26161 => x"C0C0BFA482F982F9",
-26160 => x"C0C0BFA482F982C0",
-26159 => x"C0C0BFA482F99290",
-26158 => x"C0C0BFA482F99280",
-26157 => x"C0C0BFA482F992F8",
-26156 => x"C0C0BFA482F99282",
-26155 => x"C0C0BFA482F99292",
-26154 => x"C0C0BFA482F99299",
-26153 => x"C0C0BFA482F992B0",
-26152 => x"C0C0BFA482F992A4",
-26151 => x"C0C0BFA482F992F9",
-26150 => x"C0C0BFA482F992C0",
-26149 => x"C0C0BFA482F99990",
-26148 => x"C0C0BFA482F99980",
-26147 => x"C0C0BFA482F999F8",
-26146 => x"C0C0BFA482F99982",
-26145 => x"C0C0BFA482F99992",
-26144 => x"C0C0BFA482F99999",
-26143 => x"C0C0BFA482F999B0",
-26142 => x"C0C0BFA482F999A4",
-26141 => x"C0C0BFA482F999F9",
-26140 => x"C0C0BFA482F999C0",
-26139 => x"C0C0BFA482F9B090",
-26138 => x"C0C0BFA482F9B080",
-26137 => x"C0C0BFA482F9B0F8",
-26136 => x"C0C0BFA482F9B082",
-26135 => x"C0C0BFA482F9B092",
-26134 => x"C0C0BFA482F9B099",
-26133 => x"C0C0BFA482F9B0B0",
-26132 => x"C0C0BFA482F9B0A4",
-26131 => x"C0C0BFA482F9B0F9",
-26130 => x"C0C0BFA482F9B0C0",
-26129 => x"C0C0BFA482F9A490",
-26128 => x"C0C0BFA482F9A480",
-26127 => x"C0C0BFA482F9A4F8",
-26126 => x"C0C0BFA482F9A482",
-26125 => x"C0C0BFA482F9A492",
-26124 => x"C0C0BFA482F9A499",
-26123 => x"C0C0BFA482F9A4B0",
-26122 => x"C0C0BFA482F9A4A4",
-26121 => x"C0C0BFA482F9A4F9",
-26120 => x"C0C0BFA482F9A4C0",
-26119 => x"C0C0BFA482F9F990",
-26118 => x"C0C0BFA482F9F980",
-26117 => x"C0C0BFA482F9F9F8",
-26116 => x"C0C0BFA482F9F982",
-26115 => x"C0C0BFA482F9F992",
-26114 => x"C0C0BFA482F9F999",
-26113 => x"C0C0BFA482F9F9B0",
-26112 => x"C0C0BFA482F9F9A4",
-26111 => x"C0C0BFA482F9F9F9",
-26110 => x"C0C0BFA482F9F9C0",
-26109 => x"C0C0BFA482F9C090",
-26108 => x"C0C0BFA482F9C080",
-26107 => x"C0C0BFA482F9C0F8",
-26106 => x"C0C0BFA482F9C082",
-26105 => x"C0C0BFA482F9C092",
-26104 => x"C0C0BFA482F9C099",
-26103 => x"C0C0BFA482F9C0B0",
-26102 => x"C0C0BFA482F9C0A4",
-26101 => x"C0C0BFA482F9C0F9",
-26100 => x"C0C0BFA482F9C0C0",
-26099 => x"C0C0BFA482C09090",
-26098 => x"C0C0BFA482C09080",
-26097 => x"C0C0BFA482C090F8",
-26096 => x"C0C0BFA482C09082",
-26095 => x"C0C0BFA482C09092",
-26094 => x"C0C0BFA482C09099",
-26093 => x"C0C0BFA482C090B0",
-26092 => x"C0C0BFA482C090A4",
-26091 => x"C0C0BFA482C090F9",
-26090 => x"C0C0BFA482C090C0",
-26089 => x"C0C0BFA482C08090",
-26088 => x"C0C0BFA482C08080",
-26087 => x"C0C0BFA482C080F8",
-26086 => x"C0C0BFA482C08082",
-26085 => x"C0C0BFA482C08092",
-26084 => x"C0C0BFA482C08099",
-26083 => x"C0C0BFA482C080B0",
-26082 => x"C0C0BFA482C080A4",
-26081 => x"C0C0BFA482C080F9",
-26080 => x"C0C0BFA482C080C0",
-26079 => x"C0C0BFA482C0F890",
-26078 => x"C0C0BFA482C0F880",
-26077 => x"C0C0BFA482C0F8F8",
-26076 => x"C0C0BFA482C0F882",
-26075 => x"C0C0BFA482C0F892",
-26074 => x"C0C0BFA482C0F899",
-26073 => x"C0C0BFA482C0F8B0",
-26072 => x"C0C0BFA482C0F8A4",
-26071 => x"C0C0BFA482C0F8F9",
-26070 => x"C0C0BFA482C0F8C0",
-26069 => x"C0C0BFA482C08290",
-26068 => x"C0C0BFA482C08280",
-26067 => x"C0C0BFA482C082F8",
-26066 => x"C0C0BFA482C08282",
-26065 => x"C0C0BFA482C08292",
-26064 => x"C0C0BFA482C08299",
-26063 => x"C0C0BFA482C082B0",
-26062 => x"C0C0BFA482C082A4",
-26061 => x"C0C0BFA482C082F9",
-26060 => x"C0C0BFA482C082C0",
-26059 => x"C0C0BFA482C09290",
-26058 => x"C0C0BFA482C09280",
-26057 => x"C0C0BFA482C092F8",
-26056 => x"C0C0BFA482C09282",
-26055 => x"C0C0BFA482C09292",
-26054 => x"C0C0BFA482C09299",
-26053 => x"C0C0BFA482C092B0",
-26052 => x"C0C0BFA482C092A4",
-26051 => x"C0C0BFA482C092F9",
-26050 => x"C0C0BFA482C092C0",
-26049 => x"C0C0BFA482C09990",
-26048 => x"C0C0BFA482C09980",
-26047 => x"C0C0BFA482C099F8",
-26046 => x"C0C0BFA482C09982",
-26045 => x"C0C0BFA482C09992",
-26044 => x"C0C0BFA482C09999",
-26043 => x"C0C0BFA482C099B0",
-26042 => x"C0C0BFA482C099A4",
-26041 => x"C0C0BFA482C099F9",
-26040 => x"C0C0BFA482C099C0",
-26039 => x"C0C0BFA482C0B090",
-26038 => x"C0C0BFA482C0B080",
-26037 => x"C0C0BFA482C0B0F8",
-26036 => x"C0C0BFA482C0B082",
-26035 => x"C0C0BFA482C0B092",
-26034 => x"C0C0BFA482C0B099",
-26033 => x"C0C0BFA482C0B0B0",
-26032 => x"C0C0BFA482C0B0A4",
-26031 => x"C0C0BFA482C0B0F9",
-26030 => x"C0C0BFA482C0B0C0",
-26029 => x"C0C0BFA482C0A490",
-26028 => x"C0C0BFA482C0A480",
-26027 => x"C0C0BFA482C0A4F8",
-26026 => x"C0C0BFA482C0A482",
-26025 => x"C0C0BFA482C0A492",
-26024 => x"C0C0BFA482C0A499",
-26023 => x"C0C0BFA482C0A4B0",
-26022 => x"C0C0BFA482C0A4A4",
-26021 => x"C0C0BFA482C0A4F9",
-26020 => x"C0C0BFA482C0A4C0",
-26019 => x"C0C0BFA482C0F990",
-26018 => x"C0C0BFA482C0F980",
-26017 => x"C0C0BFA482C0F9F8",
-26016 => x"C0C0BFA482C0F982",
-26015 => x"C0C0BFA482C0F992",
-26014 => x"C0C0BFA482C0F999",
-26013 => x"C0C0BFA482C0F9B0",
-26012 => x"C0C0BFA482C0F9A4",
-26011 => x"C0C0BFA482C0F9F9",
-26010 => x"C0C0BFA482C0F9C0",
-26009 => x"C0C0BFA482C0C090",
-26008 => x"C0C0BFA482C0C080",
-26007 => x"C0C0BFA482C0C0F8",
-26006 => x"C0C0BFA482C0C082",
-26005 => x"C0C0BFA482C0C092",
-26004 => x"C0C0BFA482C0C099",
-26003 => x"C0C0BFA482C0C0B0",
-26002 => x"C0C0BFA482C0C0A4",
-26001 => x"C0C0BFA482C0C0F9",
-26000 => x"C0C0BFA482C0C0C0",
-25999 => x"C0C0BFA492909090",
-25998 => x"C0C0BFA492909080",
-25997 => x"C0C0BFA4929090F8",
-25996 => x"C0C0BFA492909082",
-25995 => x"C0C0BFA492909092",
-25994 => x"C0C0BFA492909099",
-25993 => x"C0C0BFA4929090B0",
-25992 => x"C0C0BFA4929090A4",
-25991 => x"C0C0BFA4929090F9",
-25990 => x"C0C0BFA4929090C0",
-25989 => x"C0C0BFA492908090",
-25988 => x"C0C0BFA492908080",
-25987 => x"C0C0BFA4929080F8",
-25986 => x"C0C0BFA492908082",
-25985 => x"C0C0BFA492908092",
-25984 => x"C0C0BFA492908099",
-25983 => x"C0C0BFA4929080B0",
-25982 => x"C0C0BFA4929080A4",
-25981 => x"C0C0BFA4929080F9",
-25980 => x"C0C0BFA4929080C0",
-25979 => x"C0C0BFA49290F890",
-25978 => x"C0C0BFA49290F880",
-25977 => x"C0C0BFA49290F8F8",
-25976 => x"C0C0BFA49290F882",
-25975 => x"C0C0BFA49290F892",
-25974 => x"C0C0BFA49290F899",
-25973 => x"C0C0BFA49290F8B0",
-25972 => x"C0C0BFA49290F8A4",
-25971 => x"C0C0BFA49290F8F9",
-25970 => x"C0C0BFA49290F8C0",
-25969 => x"C0C0BFA492908290",
-25968 => x"C0C0BFA492908280",
-25967 => x"C0C0BFA4929082F8",
-25966 => x"C0C0BFA492908282",
-25965 => x"C0C0BFA492908292",
-25964 => x"C0C0BFA492908299",
-25963 => x"C0C0BFA4929082B0",
-25962 => x"C0C0BFA4929082A4",
-25961 => x"C0C0BFA4929082F9",
-25960 => x"C0C0BFA4929082C0",
-25959 => x"C0C0BFA492909290",
-25958 => x"C0C0BFA492909280",
-25957 => x"C0C0BFA4929092F8",
-25956 => x"C0C0BFA492909282",
-25955 => x"C0C0BFA492909292",
-25954 => x"C0C0BFA492909299",
-25953 => x"C0C0BFA4929092B0",
-25952 => x"C0C0BFA4929092A4",
-25951 => x"C0C0BFA4929092F9",
-25950 => x"C0C0BFA4929092C0",
-25949 => x"C0C0BFA492909990",
-25948 => x"C0C0BFA492909980",
-25947 => x"C0C0BFA4929099F8",
-25946 => x"C0C0BFA492909982",
-25945 => x"C0C0BFA492909992",
-25944 => x"C0C0BFA492909999",
-25943 => x"C0C0BFA4929099B0",
-25942 => x"C0C0BFA4929099A4",
-25941 => x"C0C0BFA4929099F9",
-25940 => x"C0C0BFA4929099C0",
-25939 => x"C0C0BFA49290B090",
-25938 => x"C0C0BFA49290B080",
-25937 => x"C0C0BFA49290B0F8",
-25936 => x"C0C0BFA49290B082",
-25935 => x"C0C0BFA49290B092",
-25934 => x"C0C0BFA49290B099",
-25933 => x"C0C0BFA49290B0B0",
-25932 => x"C0C0BFA49290B0A4",
-25931 => x"C0C0BFA49290B0F9",
-25930 => x"C0C0BFA49290B0C0",
-25929 => x"C0C0BFA49290A490",
-25928 => x"C0C0BFA49290A480",
-25927 => x"C0C0BFA49290A4F8",
-25926 => x"C0C0BFA49290A482",
-25925 => x"C0C0BFA49290A492",
-25924 => x"C0C0BFA49290A499",
-25923 => x"C0C0BFA49290A4B0",
-25922 => x"C0C0BFA49290A4A4",
-25921 => x"C0C0BFA49290A4F9",
-25920 => x"C0C0BFA49290A4C0",
-25919 => x"C0C0BFA49290F990",
-25918 => x"C0C0BFA49290F980",
-25917 => x"C0C0BFA49290F9F8",
-25916 => x"C0C0BFA49290F982",
-25915 => x"C0C0BFA49290F992",
-25914 => x"C0C0BFA49290F999",
-25913 => x"C0C0BFA49290F9B0",
-25912 => x"C0C0BFA49290F9A4",
-25911 => x"C0C0BFA49290F9F9",
-25910 => x"C0C0BFA49290F9C0",
-25909 => x"C0C0BFA49290C090",
-25908 => x"C0C0BFA49290C080",
-25907 => x"C0C0BFA49290C0F8",
-25906 => x"C0C0BFA49290C082",
-25905 => x"C0C0BFA49290C092",
-25904 => x"C0C0BFA49290C099",
-25903 => x"C0C0BFA49290C0B0",
-25902 => x"C0C0BFA49290C0A4",
-25901 => x"C0C0BFA49290C0F9",
-25900 => x"C0C0BFA49290C0C0",
-25899 => x"C0C0BFA492809090",
-25898 => x"C0C0BFA492809080",
-25897 => x"C0C0BFA4928090F8",
-25896 => x"C0C0BFA492809082",
-25895 => x"C0C0BFA492809092",
-25894 => x"C0C0BFA492809099",
-25893 => x"C0C0BFA4928090B0",
-25892 => x"C0C0BFA4928090A4",
-25891 => x"C0C0BFA4928090F9",
-25890 => x"C0C0BFA4928090C0",
-25889 => x"C0C0BFA492808090",
-25888 => x"C0C0BFA492808080",
-25887 => x"C0C0BFA4928080F8",
-25886 => x"C0C0BFA492808082",
-25885 => x"C0C0BFA492808092",
-25884 => x"C0C0BFA492808099",
-25883 => x"C0C0BFA4928080B0",
-25882 => x"C0C0BFA4928080A4",
-25881 => x"C0C0BFA4928080F9",
-25880 => x"C0C0BFA4928080C0",
-25879 => x"C0C0BFA49280F890",
-25878 => x"C0C0BFA49280F880",
-25877 => x"C0C0BFA49280F8F8",
-25876 => x"C0C0BFA49280F882",
-25875 => x"C0C0BFA49280F892",
-25874 => x"C0C0BFA49280F899",
-25873 => x"C0C0BFA49280F8B0",
-25872 => x"C0C0BFA49280F8A4",
-25871 => x"C0C0BFA49280F8F9",
-25870 => x"C0C0BFA49280F8C0",
-25869 => x"C0C0BFA492808290",
-25868 => x"C0C0BFA492808280",
-25867 => x"C0C0BFA4928082F8",
-25866 => x"C0C0BFA492808282",
-25865 => x"C0C0BFA492808292",
-25864 => x"C0C0BFA492808299",
-25863 => x"C0C0BFA4928082B0",
-25862 => x"C0C0BFA4928082A4",
-25861 => x"C0C0BFA4928082F9",
-25860 => x"C0C0BFA4928082C0",
-25859 => x"C0C0BFA492809290",
-25858 => x"C0C0BFA492809280",
-25857 => x"C0C0BFA4928092F8",
-25856 => x"C0C0BFA492809282",
-25855 => x"C0C0BFA492809292",
-25854 => x"C0C0BFA492809299",
-25853 => x"C0C0BFA4928092B0",
-25852 => x"C0C0BFA4928092A4",
-25851 => x"C0C0BFA4928092F9",
-25850 => x"C0C0BFA4928092C0",
-25849 => x"C0C0BFA492809990",
-25848 => x"C0C0BFA492809980",
-25847 => x"C0C0BFA4928099F8",
-25846 => x"C0C0BFA492809982",
-25845 => x"C0C0BFA492809992",
-25844 => x"C0C0BFA492809999",
-25843 => x"C0C0BFA4928099B0",
-25842 => x"C0C0BFA4928099A4",
-25841 => x"C0C0BFA4928099F9",
-25840 => x"C0C0BFA4928099C0",
-25839 => x"C0C0BFA49280B090",
-25838 => x"C0C0BFA49280B080",
-25837 => x"C0C0BFA49280B0F8",
-25836 => x"C0C0BFA49280B082",
-25835 => x"C0C0BFA49280B092",
-25834 => x"C0C0BFA49280B099",
-25833 => x"C0C0BFA49280B0B0",
-25832 => x"C0C0BFA49280B0A4",
-25831 => x"C0C0BFA49280B0F9",
-25830 => x"C0C0BFA49280B0C0",
-25829 => x"C0C0BFA49280A490",
-25828 => x"C0C0BFA49280A480",
-25827 => x"C0C0BFA49280A4F8",
-25826 => x"C0C0BFA49280A482",
-25825 => x"C0C0BFA49280A492",
-25824 => x"C0C0BFA49280A499",
-25823 => x"C0C0BFA49280A4B0",
-25822 => x"C0C0BFA49280A4A4",
-25821 => x"C0C0BFA49280A4F9",
-25820 => x"C0C0BFA49280A4C0",
-25819 => x"C0C0BFA49280F990",
-25818 => x"C0C0BFA49280F980",
-25817 => x"C0C0BFA49280F9F8",
-25816 => x"C0C0BFA49280F982",
-25815 => x"C0C0BFA49280F992",
-25814 => x"C0C0BFA49280F999",
-25813 => x"C0C0BFA49280F9B0",
-25812 => x"C0C0BFA49280F9A4",
-25811 => x"C0C0BFA49280F9F9",
-25810 => x"C0C0BFA49280F9C0",
-25809 => x"C0C0BFA49280C090",
-25808 => x"C0C0BFA49280C080",
-25807 => x"C0C0BFA49280C0F8",
-25806 => x"C0C0BFA49280C082",
-25805 => x"C0C0BFA49280C092",
-25804 => x"C0C0BFA49280C099",
-25803 => x"C0C0BFA49280C0B0",
-25802 => x"C0C0BFA49280C0A4",
-25801 => x"C0C0BFA49280C0F9",
-25800 => x"C0C0BFA49280C0C0",
-25799 => x"C0C0BFA492F89090",
-25798 => x"C0C0BFA492F89080",
-25797 => x"C0C0BFA492F890F8",
-25796 => x"C0C0BFA492F89082",
-25795 => x"C0C0BFA492F89092",
-25794 => x"C0C0BFA492F89099",
-25793 => x"C0C0BFA492F890B0",
-25792 => x"C0C0BFA492F890A4",
-25791 => x"C0C0BFA492F890F9",
-25790 => x"C0C0BFA492F890C0",
-25789 => x"C0C0BFA492F88090",
-25788 => x"C0C0BFA492F88080",
-25787 => x"C0C0BFA492F880F8",
-25786 => x"C0C0BFA492F88082",
-25785 => x"C0C0BFA492F88092",
-25784 => x"C0C0BFA492F88099",
-25783 => x"C0C0BFA492F880B0",
-25782 => x"C0C0BFA492F880A4",
-25781 => x"C0C0BFA492F880F9",
-25780 => x"C0C0BFA492F880C0",
-25779 => x"C0C0BFA492F8F890",
-25778 => x"C0C0BFA492F8F880",
-25777 => x"C0C0BFA492F8F8F8",
-25776 => x"C0C0BFA492F8F882",
-25775 => x"C0C0BFA492F8F892",
-25774 => x"C0C0BFA492F8F899",
-25773 => x"C0C0BFA492F8F8B0",
-25772 => x"C0C0BFA492F8F8A4",
-25771 => x"C0C0BFA492F8F8F9",
-25770 => x"C0C0BFA492F8F8C0",
-25769 => x"C0C0BFA492F88290",
-25768 => x"C0C0BFA492F88280",
-25767 => x"C0C0BFA492F882F8",
-25766 => x"C0C0BFA492F88282",
-25765 => x"C0C0BFA492F88292",
-25764 => x"C0C0BFA492F88299",
-25763 => x"C0C0BFA492F882B0",
-25762 => x"C0C0BFA492F882A4",
-25761 => x"C0C0BFA492F882F9",
-25760 => x"C0C0BFA492F882C0",
-25759 => x"C0C0BFA492F89290",
-25758 => x"C0C0BFA492F89280",
-25757 => x"C0C0BFA492F892F8",
-25756 => x"C0C0BFA492F89282",
-25755 => x"C0C0BFA492F89292",
-25754 => x"C0C0BFA492F89299",
-25753 => x"C0C0BFA492F892B0",
-25752 => x"C0C0BFA492F892A4",
-25751 => x"C0C0BFA492F892F9",
-25750 => x"C0C0BFA492F892C0",
-25749 => x"C0C0BFA492F89990",
-25748 => x"C0C0BFA492F89980",
-25747 => x"C0C0BFA492F899F8",
-25746 => x"C0C0BFA492F89982",
-25745 => x"C0C0BFA492F89992",
-25744 => x"C0C0BFA492F89999",
-25743 => x"C0C0BFA492F899B0",
-25742 => x"C0C0BFA492F899A4",
-25741 => x"C0C0BFA492F899F9",
-25740 => x"C0C0BFA492F899C0",
-25739 => x"C0C0BFA492F8B090",
-25738 => x"C0C0BFA492F8B080",
-25737 => x"C0C0BFA492F8B0F8",
-25736 => x"C0C0BFA492F8B082",
-25735 => x"C0C0BFA492F8B092",
-25734 => x"C0C0BFA492F8B099",
-25733 => x"C0C0BFA492F8B0B0",
-25732 => x"C0C0BFA492F8B0A4",
-25731 => x"C0C0BFA492F8B0F9",
-25730 => x"C0C0BFA492F8B0C0",
-25729 => x"C0C0BFA492F8A490",
-25728 => x"C0C0BFA492F8A480",
-25727 => x"C0C0BFA492F8A4F8",
-25726 => x"C0C0BFA492F8A482",
-25725 => x"C0C0BFA492F8A492",
-25724 => x"C0C0BFA492F8A499",
-25723 => x"C0C0BFA492F8A4B0",
-25722 => x"C0C0BFA492F8A4A4",
-25721 => x"C0C0BFA492F8A4F9",
-25720 => x"C0C0BFA492F8A4C0",
-25719 => x"C0C0BFA492F8F990",
-25718 => x"C0C0BFA492F8F980",
-25717 => x"C0C0BFA492F8F9F8",
-25716 => x"C0C0BFA492F8F982",
-25715 => x"C0C0BFA492F8F992",
-25714 => x"C0C0BFA492F8F999",
-25713 => x"C0C0BFA492F8F9B0",
-25712 => x"C0C0BFA492F8F9A4",
-25711 => x"C0C0BFA492F8F9F9",
-25710 => x"C0C0BFA492F8F9C0",
-25709 => x"C0C0BFA492F8C090",
-25708 => x"C0C0BFA492F8C080",
-25707 => x"C0C0BFA492F8C0F8",
-25706 => x"C0C0BFA492F8C082",
-25705 => x"C0C0BFA492F8C092",
-25704 => x"C0C0BFA492F8C099",
-25703 => x"C0C0BFA492F8C0B0",
-25702 => x"C0C0BFA492F8C0A4",
-25701 => x"C0C0BFA492F8C0F9",
-25700 => x"C0C0BFA492F8C0C0",
-25699 => x"C0C0BFA492829090",
-25698 => x"C0C0BFA492829080",
-25697 => x"C0C0BFA4928290F8",
-25696 => x"C0C0BFA492829082",
-25695 => x"C0C0BFA492829092",
-25694 => x"C0C0BFA492829099",
-25693 => x"C0C0BFA4928290B0",
-25692 => x"C0C0BFA4928290A4",
-25691 => x"C0C0BFA4928290F9",
-25690 => x"C0C0BFA4928290C0",
-25689 => x"C0C0BFA492828090",
-25688 => x"C0C0BFA492828080",
-25687 => x"C0C0BFA4928280F8",
-25686 => x"C0C0BFA492828082",
-25685 => x"C0C0BFA492828092",
-25684 => x"C0C0BFA492828099",
-25683 => x"C0C0BFA4928280B0",
-25682 => x"C0C0BFA4928280A4",
-25681 => x"C0C0BFA4928280F9",
-25680 => x"C0C0BFA4928280C0",
-25679 => x"C0C0BFA49282F890",
-25678 => x"C0C0BFA49282F880",
-25677 => x"C0C0BFA49282F8F8",
-25676 => x"C0C0BFA49282F882",
-25675 => x"C0C0BFA49282F892",
-25674 => x"C0C0BFA49282F899",
-25673 => x"C0C0BFA49282F8B0",
-25672 => x"C0C0BFA49282F8A4",
-25671 => x"C0C0BFA49282F8F9",
-25670 => x"C0C0BFA49282F8C0",
-25669 => x"C0C0BFA492828290",
-25668 => x"C0C0BFA492828280",
-25667 => x"C0C0BFA4928282F8",
-25666 => x"C0C0BFA492828282",
-25665 => x"C0C0BFA492828292",
-25664 => x"C0C0BFA492828299",
-25663 => x"C0C0BFA4928282B0",
-25662 => x"C0C0BFA4928282A4",
-25661 => x"C0C0BFA4928282F9",
-25660 => x"C0C0BFA4928282C0",
-25659 => x"C0C0BFA492829290",
-25658 => x"C0C0BFA492829280",
-25657 => x"C0C0BFA4928292F8",
-25656 => x"C0C0BFA492829282",
-25655 => x"C0C0BFA492829292",
-25654 => x"C0C0BFA492829299",
-25653 => x"C0C0BFA4928292B0",
-25652 => x"C0C0BFA4928292A4",
-25651 => x"C0C0BFA4928292F9",
-25650 => x"C0C0BFA4928292C0",
-25649 => x"C0C0BFA492829990",
-25648 => x"C0C0BFA492829980",
-25647 => x"C0C0BFA4928299F8",
-25646 => x"C0C0BFA492829982",
-25645 => x"C0C0BFA492829992",
-25644 => x"C0C0BFA492829999",
-25643 => x"C0C0BFA4928299B0",
-25642 => x"C0C0BFA4928299A4",
-25641 => x"C0C0BFA4928299F9",
-25640 => x"C0C0BFA4928299C0",
-25639 => x"C0C0BFA49282B090",
-25638 => x"C0C0BFA49282B080",
-25637 => x"C0C0BFA49282B0F8",
-25636 => x"C0C0BFA49282B082",
-25635 => x"C0C0BFA49282B092",
-25634 => x"C0C0BFA49282B099",
-25633 => x"C0C0BFA49282B0B0",
-25632 => x"C0C0BFA49282B0A4",
-25631 => x"C0C0BFA49282B0F9",
-25630 => x"C0C0BFA49282B0C0",
-25629 => x"C0C0BFA49282A490",
-25628 => x"C0C0BFA49282A480",
-25627 => x"C0C0BFA49282A4F8",
-25626 => x"C0C0BFA49282A482",
-25625 => x"C0C0BFA49282A492",
-25624 => x"C0C0BFA49282A499",
-25623 => x"C0C0BFA49282A4B0",
-25622 => x"C0C0BFA49282A4A4",
-25621 => x"C0C0BFA49282A4F9",
-25620 => x"C0C0BFA49282A4C0",
-25619 => x"C0C0BFA49282F990",
-25618 => x"C0C0BFA49282F980",
-25617 => x"C0C0BFA49282F9F8",
-25616 => x"C0C0BFA49282F982",
-25615 => x"C0C0BFA49282F992",
-25614 => x"C0C0BFA49282F999",
-25613 => x"C0C0BFA49282F9B0",
-25612 => x"C0C0BFA49282F9A4",
-25611 => x"C0C0BFA49282F9F9",
-25610 => x"C0C0BFA49282F9C0",
-25609 => x"C0C0BFA49282C090",
-25608 => x"C0C0BFA49282C080",
-25607 => x"C0C0BFA49282C0F8",
-25606 => x"C0C0BFA49282C082",
-25605 => x"C0C0BFA49282C092",
-25604 => x"C0C0BFA49282C099",
-25603 => x"C0C0BFA49282C0B0",
-25602 => x"C0C0BFA49282C0A4",
-25601 => x"C0C0BFA49282C0F9",
-25600 => x"C0C0BFA49282C0C0",
-25599 => x"C0C0BFA492929090",
-25598 => x"C0C0BFA492929080",
-25597 => x"C0C0BFA4929290F8",
-25596 => x"C0C0BFA492929082",
-25595 => x"C0C0BFA492929092",
-25594 => x"C0C0BFA492929099",
-25593 => x"C0C0BFA4929290B0",
-25592 => x"C0C0BFA4929290A4",
-25591 => x"C0C0BFA4929290F9",
-25590 => x"C0C0BFA4929290C0",
-25589 => x"C0C0BFA492928090",
-25588 => x"C0C0BFA492928080",
-25587 => x"C0C0BFA4929280F8",
-25586 => x"C0C0BFA492928082",
-25585 => x"C0C0BFA492928092",
-25584 => x"C0C0BFA492928099",
-25583 => x"C0C0BFA4929280B0",
-25582 => x"C0C0BFA4929280A4",
-25581 => x"C0C0BFA4929280F9",
-25580 => x"C0C0BFA4929280C0",
-25579 => x"C0C0BFA49292F890",
-25578 => x"C0C0BFA49292F880",
-25577 => x"C0C0BFA49292F8F8",
-25576 => x"C0C0BFA49292F882",
-25575 => x"C0C0BFA49292F892",
-25574 => x"C0C0BFA49292F899",
-25573 => x"C0C0BFA49292F8B0",
-25572 => x"C0C0BFA49292F8A4",
-25571 => x"C0C0BFA49292F8F9",
-25570 => x"C0C0BFA49292F8C0",
-25569 => x"C0C0BFA492928290",
-25568 => x"C0C0BFA492928280",
-25567 => x"C0C0BFA4929282F8",
-25566 => x"C0C0BFA492928282",
-25565 => x"C0C0BFA492928292",
-25564 => x"C0C0BFA492928299",
-25563 => x"C0C0BFA4929282B0",
-25562 => x"C0C0BFA4929282A4",
-25561 => x"C0C0BFA4929282F9",
-25560 => x"C0C0BFA4929282C0",
-25559 => x"C0C0BFA492929290",
-25558 => x"C0C0BFA492929280",
-25557 => x"C0C0BFA4929292F8",
-25556 => x"C0C0BFA492929282",
-25555 => x"C0C0BFA492929292",
-25554 => x"C0C0BFA492929299",
-25553 => x"C0C0BFA4929292B0",
-25552 => x"C0C0BFA4929292A4",
-25551 => x"C0C0BFA4929292F9",
-25550 => x"C0C0BFA4929292C0",
-25549 => x"C0C0BFA492929990",
-25548 => x"C0C0BFA492929980",
-25547 => x"C0C0BFA4929299F8",
-25546 => x"C0C0BFA492929982",
-25545 => x"C0C0BFA492929992",
-25544 => x"C0C0BFA492929999",
-25543 => x"C0C0BFA4929299B0",
-25542 => x"C0C0BFA4929299A4",
-25541 => x"C0C0BFA4929299F9",
-25540 => x"C0C0BFA4929299C0",
-25539 => x"C0C0BFA49292B090",
-25538 => x"C0C0BFA49292B080",
-25537 => x"C0C0BFA49292B0F8",
-25536 => x"C0C0BFA49292B082",
-25535 => x"C0C0BFA49292B092",
-25534 => x"C0C0BFA49292B099",
-25533 => x"C0C0BFA49292B0B0",
-25532 => x"C0C0BFA49292B0A4",
-25531 => x"C0C0BFA49292B0F9",
-25530 => x"C0C0BFA49292B0C0",
-25529 => x"C0C0BFA49292A490",
-25528 => x"C0C0BFA49292A480",
-25527 => x"C0C0BFA49292A4F8",
-25526 => x"C0C0BFA49292A482",
-25525 => x"C0C0BFA49292A492",
-25524 => x"C0C0BFA49292A499",
-25523 => x"C0C0BFA49292A4B0",
-25522 => x"C0C0BFA49292A4A4",
-25521 => x"C0C0BFA49292A4F9",
-25520 => x"C0C0BFA49292A4C0",
-25519 => x"C0C0BFA49292F990",
-25518 => x"C0C0BFA49292F980",
-25517 => x"C0C0BFA49292F9F8",
-25516 => x"C0C0BFA49292F982",
-25515 => x"C0C0BFA49292F992",
-25514 => x"C0C0BFA49292F999",
-25513 => x"C0C0BFA49292F9B0",
-25512 => x"C0C0BFA49292F9A4",
-25511 => x"C0C0BFA49292F9F9",
-25510 => x"C0C0BFA49292F9C0",
-25509 => x"C0C0BFA49292C090",
-25508 => x"C0C0BFA49292C080",
-25507 => x"C0C0BFA49292C0F8",
-25506 => x"C0C0BFA49292C082",
-25505 => x"C0C0BFA49292C092",
-25504 => x"C0C0BFA49292C099",
-25503 => x"C0C0BFA49292C0B0",
-25502 => x"C0C0BFA49292C0A4",
-25501 => x"C0C0BFA49292C0F9",
-25500 => x"C0C0BFA49292C0C0",
-25499 => x"C0C0BFA492999090",
-25498 => x"C0C0BFA492999080",
-25497 => x"C0C0BFA4929990F8",
-25496 => x"C0C0BFA492999082",
-25495 => x"C0C0BFA492999092",
-25494 => x"C0C0BFA492999099",
-25493 => x"C0C0BFA4929990B0",
-25492 => x"C0C0BFA4929990A4",
-25491 => x"C0C0BFA4929990F9",
-25490 => x"C0C0BFA4929990C0",
-25489 => x"C0C0BFA492998090",
-25488 => x"C0C0BFA492998080",
-25487 => x"C0C0BFA4929980F8",
-25486 => x"C0C0BFA492998082",
-25485 => x"C0C0BFA492998092",
-25484 => x"C0C0BFA492998099",
-25483 => x"C0C0BFA4929980B0",
-25482 => x"C0C0BFA4929980A4",
-25481 => x"C0C0BFA4929980F9",
-25480 => x"C0C0BFA4929980C0",
-25479 => x"C0C0BFA49299F890",
-25478 => x"C0C0BFA49299F880",
-25477 => x"C0C0BFA49299F8F8",
-25476 => x"C0C0BFA49299F882",
-25475 => x"C0C0BFA49299F892",
-25474 => x"C0C0BFA49299F899",
-25473 => x"C0C0BFA49299F8B0",
-25472 => x"C0C0BFA49299F8A4",
-25471 => x"C0C0BFA49299F8F9",
-25470 => x"C0C0BFA49299F8C0",
-25469 => x"C0C0BFA492998290",
-25468 => x"C0C0BFA492998280",
-25467 => x"C0C0BFA4929982F8",
-25466 => x"C0C0BFA492998282",
-25465 => x"C0C0BFA492998292",
-25464 => x"C0C0BFA492998299",
-25463 => x"C0C0BFA4929982B0",
-25462 => x"C0C0BFA4929982A4",
-25461 => x"C0C0BFA4929982F9",
-25460 => x"C0C0BFA4929982C0",
-25459 => x"C0C0BFA492999290",
-25458 => x"C0C0BFA492999280",
-25457 => x"C0C0BFA4929992F8",
-25456 => x"C0C0BFA492999282",
-25455 => x"C0C0BFA492999292",
-25454 => x"C0C0BFA492999299",
-25453 => x"C0C0BFA4929992B0",
-25452 => x"C0C0BFA4929992A4",
-25451 => x"C0C0BFA4929992F9",
-25450 => x"C0C0BFA4929992C0",
-25449 => x"C0C0BFA492999990",
-25448 => x"C0C0BFA492999980",
-25447 => x"C0C0BFA4929999F8",
-25446 => x"C0C0BFA492999982",
-25445 => x"C0C0BFA492999992",
-25444 => x"C0C0BFA492999999",
-25443 => x"C0C0BFA4929999B0",
-25442 => x"C0C0BFA4929999A4",
-25441 => x"C0C0BFA4929999F9",
-25440 => x"C0C0BFA4929999C0",
-25439 => x"C0C0BFA49299B090",
-25438 => x"C0C0BFA49299B080",
-25437 => x"C0C0BFA49299B0F8",
-25436 => x"C0C0BFA49299B082",
-25435 => x"C0C0BFA49299B092",
-25434 => x"C0C0BFA49299B099",
-25433 => x"C0C0BFA49299B0B0",
-25432 => x"C0C0BFA49299B0A4",
-25431 => x"C0C0BFA49299B0F9",
-25430 => x"C0C0BFA49299B0C0",
-25429 => x"C0C0BFA49299A490",
-25428 => x"C0C0BFA49299A480",
-25427 => x"C0C0BFA49299A4F8",
-25426 => x"C0C0BFA49299A482",
-25425 => x"C0C0BFA49299A492",
-25424 => x"C0C0BFA49299A499",
-25423 => x"C0C0BFA49299A4B0",
-25422 => x"C0C0BFA49299A4A4",
-25421 => x"C0C0BFA49299A4F9",
-25420 => x"C0C0BFA49299A4C0",
-25419 => x"C0C0BFA49299F990",
-25418 => x"C0C0BFA49299F980",
-25417 => x"C0C0BFA49299F9F8",
-25416 => x"C0C0BFA49299F982",
-25415 => x"C0C0BFA49299F992",
-25414 => x"C0C0BFA49299F999",
-25413 => x"C0C0BFA49299F9B0",
-25412 => x"C0C0BFA49299F9A4",
-25411 => x"C0C0BFA49299F9F9",
-25410 => x"C0C0BFA49299F9C0",
-25409 => x"C0C0BFA49299C090",
-25408 => x"C0C0BFA49299C080",
-25407 => x"C0C0BFA49299C0F8",
-25406 => x"C0C0BFA49299C082",
-25405 => x"C0C0BFA49299C092",
-25404 => x"C0C0BFA49299C099",
-25403 => x"C0C0BFA49299C0B0",
-25402 => x"C0C0BFA49299C0A4",
-25401 => x"C0C0BFA49299C0F9",
-25400 => x"C0C0BFA49299C0C0",
-25399 => x"C0C0BFA492B09090",
-25398 => x"C0C0BFA492B09080",
-25397 => x"C0C0BFA492B090F8",
-25396 => x"C0C0BFA492B09082",
-25395 => x"C0C0BFA492B09092",
-25394 => x"C0C0BFA492B09099",
-25393 => x"C0C0BFA492B090B0",
-25392 => x"C0C0BFA492B090A4",
-25391 => x"C0C0BFA492B090F9",
-25390 => x"C0C0BFA492B090C0",
-25389 => x"C0C0BFA492B08090",
-25388 => x"C0C0BFA492B08080",
-25387 => x"C0C0BFA492B080F8",
-25386 => x"C0C0BFA492B08082",
-25385 => x"C0C0BFA492B08092",
-25384 => x"C0C0BFA492B08099",
-25383 => x"C0C0BFA492B080B0",
-25382 => x"C0C0BFA492B080A4",
-25381 => x"C0C0BFA492B080F9",
-25380 => x"C0C0BFA492B080C0",
-25379 => x"C0C0BFA492B0F890",
-25378 => x"C0C0BFA492B0F880",
-25377 => x"C0C0BFA492B0F8F8",
-25376 => x"C0C0BFA492B0F882",
-25375 => x"C0C0BFA492B0F892",
-25374 => x"C0C0BFA492B0F899",
-25373 => x"C0C0BFA492B0F8B0",
-25372 => x"C0C0BFA492B0F8A4",
-25371 => x"C0C0BFA492B0F8F9",
-25370 => x"C0C0BFA492B0F8C0",
-25369 => x"C0C0BFA492B08290",
-25368 => x"C0C0BFA492B08280",
-25367 => x"C0C0BFA492B082F8",
-25366 => x"C0C0BFA492B08282",
-25365 => x"C0C0BFA492B08292",
-25364 => x"C0C0BFA492B08299",
-25363 => x"C0C0BFA492B082B0",
-25362 => x"C0C0BFA492B082A4",
-25361 => x"C0C0BFA492B082F9",
-25360 => x"C0C0BFA492B082C0",
-25359 => x"C0C0BFA492B09290",
-25358 => x"C0C0BFA492B09280",
-25357 => x"C0C0BFA492B092F8",
-25356 => x"C0C0BFA492B09282",
-25355 => x"C0C0BFA492B09292",
-25354 => x"C0C0BFA492B09299",
-25353 => x"C0C0BFA492B092B0",
-25352 => x"C0C0BFA492B092A4",
-25351 => x"C0C0BFA492B092F9",
-25350 => x"C0C0BFA492B092C0",
-25349 => x"C0C0BFA492B09990",
-25348 => x"C0C0BFA492B09980",
-25347 => x"C0C0BFA492B099F8",
-25346 => x"C0C0BFA492B09982",
-25345 => x"C0C0BFA492B09992",
-25344 => x"C0C0BFA492B09999",
-25343 => x"C0C0BFA492B099B0",
-25342 => x"C0C0BFA492B099A4",
-25341 => x"C0C0BFA492B099F9",
-25340 => x"C0C0BFA492B099C0",
-25339 => x"C0C0BFA492B0B090",
-25338 => x"C0C0BFA492B0B080",
-25337 => x"C0C0BFA492B0B0F8",
-25336 => x"C0C0BFA492B0B082",
-25335 => x"C0C0BFA492B0B092",
-25334 => x"C0C0BFA492B0B099",
-25333 => x"C0C0BFA492B0B0B0",
-25332 => x"C0C0BFA492B0B0A4",
-25331 => x"C0C0BFA492B0B0F9",
-25330 => x"C0C0BFA492B0B0C0",
-25329 => x"C0C0BFA492B0A490",
-25328 => x"C0C0BFA492B0A480",
-25327 => x"C0C0BFA492B0A4F8",
-25326 => x"C0C0BFA492B0A482",
-25325 => x"C0C0BFA492B0A492",
-25324 => x"C0C0BFA492B0A499",
-25323 => x"C0C0BFA492B0A4B0",
-25322 => x"C0C0BFA492B0A4A4",
-25321 => x"C0C0BFA492B0A4F9",
-25320 => x"C0C0BFA492B0A4C0",
-25319 => x"C0C0BFA492B0F990",
-25318 => x"C0C0BFA492B0F980",
-25317 => x"C0C0BFA492B0F9F8",
-25316 => x"C0C0BFA492B0F982",
-25315 => x"C0C0BFA492B0F992",
-25314 => x"C0C0BFA492B0F999",
-25313 => x"C0C0BFA492B0F9B0",
-25312 => x"C0C0BFA492B0F9A4",
-25311 => x"C0C0BFA492B0F9F9",
-25310 => x"C0C0BFA492B0F9C0",
-25309 => x"C0C0BFA492B0C090",
-25308 => x"C0C0BFA492B0C080",
-25307 => x"C0C0BFA492B0C0F8",
-25306 => x"C0C0BFA492B0C082",
-25305 => x"C0C0BFA492B0C092",
-25304 => x"C0C0BFA492B0C099",
-25303 => x"C0C0BFA492B0C0B0",
-25302 => x"C0C0BFA492B0C0A4",
-25301 => x"C0C0BFA492B0C0F9",
-25300 => x"C0C0BFA492B0C0C0",
-25299 => x"C0C0BFA492A49090",
-25298 => x"C0C0BFA492A49080",
-25297 => x"C0C0BFA492A490F8",
-25296 => x"C0C0BFA492A49082",
-25295 => x"C0C0BFA492A49092",
-25294 => x"C0C0BFA492A49099",
-25293 => x"C0C0BFA492A490B0",
-25292 => x"C0C0BFA492A490A4",
-25291 => x"C0C0BFA492A490F9",
-25290 => x"C0C0BFA492A490C0",
-25289 => x"C0C0BFA492A48090",
-25288 => x"C0C0BFA492A48080",
-25287 => x"C0C0BFA492A480F8",
-25286 => x"C0C0BFA492A48082",
-25285 => x"C0C0BFA492A48092",
-25284 => x"C0C0BFA492A48099",
-25283 => x"C0C0BFA492A480B0",
-25282 => x"C0C0BFA492A480A4",
-25281 => x"C0C0BFA492A480F9",
-25280 => x"C0C0BFA492A480C0",
-25279 => x"C0C0BFA492A4F890",
-25278 => x"C0C0BFA492A4F880",
-25277 => x"C0C0BFA492A4F8F8",
-25276 => x"C0C0BFA492A4F882",
-25275 => x"C0C0BFA492A4F892",
-25274 => x"C0C0BFA492A4F899",
-25273 => x"C0C0BFA492A4F8B0",
-25272 => x"C0C0BFA492A4F8A4",
-25271 => x"C0C0BFA492A4F8F9",
-25270 => x"C0C0BFA492A4F8C0",
-25269 => x"C0C0BFA492A48290",
-25268 => x"C0C0BFA492A48280",
-25267 => x"C0C0BFA492A482F8",
-25266 => x"C0C0BFA492A48282",
-25265 => x"C0C0BFA492A48292",
-25264 => x"C0C0BFA492A48299",
-25263 => x"C0C0BFA492A482B0",
-25262 => x"C0C0BFA492A482A4",
-25261 => x"C0C0BFA492A482F9",
-25260 => x"C0C0BFA492A482C0",
-25259 => x"C0C0BFA492A49290",
-25258 => x"C0C0BFA492A49280",
-25257 => x"C0C0BFA492A492F8",
-25256 => x"C0C0BFA492A49282",
-25255 => x"C0C0BFA492A49292",
-25254 => x"C0C0BFA492A49299",
-25253 => x"C0C0BFA492A492B0",
-25252 => x"C0C0BFA492A492A4",
-25251 => x"C0C0BFA492A492F9",
-25250 => x"C0C0BFA492A492C0",
-25249 => x"C0C0BFA492A49990",
-25248 => x"C0C0BFA492A49980",
-25247 => x"C0C0BFA492A499F8",
-25246 => x"C0C0BFA492A49982",
-25245 => x"C0C0BFA492A49992",
-25244 => x"C0C0BFA492A49999",
-25243 => x"C0C0BFA492A499B0",
-25242 => x"C0C0BFA492A499A4",
-25241 => x"C0C0BFA492A499F9",
-25240 => x"C0C0BFA492A499C0",
-25239 => x"C0C0BFA492A4B090",
-25238 => x"C0C0BFA492A4B080",
-25237 => x"C0C0BFA492A4B0F8",
-25236 => x"C0C0BFA492A4B082",
-25235 => x"C0C0BFA492A4B092",
-25234 => x"C0C0BFA492A4B099",
-25233 => x"C0C0BFA492A4B0B0",
-25232 => x"C0C0BFA492A4B0A4",
-25231 => x"C0C0BFA492A4B0F9",
-25230 => x"C0C0BFA492A4B0C0",
-25229 => x"C0C0BFA492A4A490",
-25228 => x"C0C0BFA492A4A480",
-25227 => x"C0C0BFA492A4A4F8",
-25226 => x"C0C0BFA492A4A482",
-25225 => x"C0C0BFA492A4A492",
-25224 => x"C0C0BFA492A4A499",
-25223 => x"C0C0BFA492A4A4B0",
-25222 => x"C0C0BFA492A4A4A4",
-25221 => x"C0C0BFA492A4A4F9",
-25220 => x"C0C0BFA492A4A4C0",
-25219 => x"C0C0BFA492A4F990",
-25218 => x"C0C0BFA492A4F980",
-25217 => x"C0C0BFA492A4F9F8",
-25216 => x"C0C0BFA492A4F982",
-25215 => x"C0C0BFA492A4F992",
-25214 => x"C0C0BFA492A4F999",
-25213 => x"C0C0BFA492A4F9B0",
-25212 => x"C0C0BFA492A4F9A4",
-25211 => x"C0C0BFA492A4F9F9",
-25210 => x"C0C0BFA492A4F9C0",
-25209 => x"C0C0BFA492A4C090",
-25208 => x"C0C0BFA492A4C080",
-25207 => x"C0C0BFA492A4C0F8",
-25206 => x"C0C0BFA492A4C082",
-25205 => x"C0C0BFA492A4C092",
-25204 => x"C0C0BFA492A4C099",
-25203 => x"C0C0BFA492A4C0B0",
-25202 => x"C0C0BFA492A4C0A4",
-25201 => x"C0C0BFA492A4C0F9",
-25200 => x"C0C0BFA492A4C0C0",
-25199 => x"C0C0BFA492F99090",
-25198 => x"C0C0BFA492F99080",
-25197 => x"C0C0BFA492F990F8",
-25196 => x"C0C0BFA492F99082",
-25195 => x"C0C0BFA492F99092",
-25194 => x"C0C0BFA492F99099",
-25193 => x"C0C0BFA492F990B0",
-25192 => x"C0C0BFA492F990A4",
-25191 => x"C0C0BFA492F990F9",
-25190 => x"C0C0BFA492F990C0",
-25189 => x"C0C0BFA492F98090",
-25188 => x"C0C0BFA492F98080",
-25187 => x"C0C0BFA492F980F8",
-25186 => x"C0C0BFA492F98082",
-25185 => x"C0C0BFA492F98092",
-25184 => x"C0C0BFA492F98099",
-25183 => x"C0C0BFA492F980B0",
-25182 => x"C0C0BFA492F980A4",
-25181 => x"C0C0BFA492F980F9",
-25180 => x"C0C0BFA492F980C0",
-25179 => x"C0C0BFA492F9F890",
-25178 => x"C0C0BFA492F9F880",
-25177 => x"C0C0BFA492F9F8F8",
-25176 => x"C0C0BFA492F9F882",
-25175 => x"C0C0BFA492F9F892",
-25174 => x"C0C0BFA492F9F899",
-25173 => x"C0C0BFA492F9F8B0",
-25172 => x"C0C0BFA492F9F8A4",
-25171 => x"C0C0BFA492F9F8F9",
-25170 => x"C0C0BFA492F9F8C0",
-25169 => x"C0C0BFA492F98290",
-25168 => x"C0C0BFA492F98280",
-25167 => x"C0C0BFA492F982F8",
-25166 => x"C0C0BFA492F98282",
-25165 => x"C0C0BFA492F98292",
-25164 => x"C0C0BFA492F98299",
-25163 => x"C0C0BFA492F982B0",
-25162 => x"C0C0BFA492F982A4",
-25161 => x"C0C0BFA492F982F9",
-25160 => x"C0C0BFA492F982C0",
-25159 => x"C0C0BFA492F99290",
-25158 => x"C0C0BFA492F99280",
-25157 => x"C0C0BFA492F992F8",
-25156 => x"C0C0BFA492F99282",
-25155 => x"C0C0BFA492F99292",
-25154 => x"C0C0BFA492F99299",
-25153 => x"C0C0BFA492F992B0",
-25152 => x"C0C0BFA492F992A4",
-25151 => x"C0C0BFA492F992F9",
-25150 => x"C0C0BFA492F992C0",
-25149 => x"C0C0BFA492F99990",
-25148 => x"C0C0BFA492F99980",
-25147 => x"C0C0BFA492F999F8",
-25146 => x"C0C0BFA492F99982",
-25145 => x"C0C0BFA492F99992",
-25144 => x"C0C0BFA492F99999",
-25143 => x"C0C0BFA492F999B0",
-25142 => x"C0C0BFA492F999A4",
-25141 => x"C0C0BFA492F999F9",
-25140 => x"C0C0BFA492F999C0",
-25139 => x"C0C0BFA492F9B090",
-25138 => x"C0C0BFA492F9B080",
-25137 => x"C0C0BFA492F9B0F8",
-25136 => x"C0C0BFA492F9B082",
-25135 => x"C0C0BFA492F9B092",
-25134 => x"C0C0BFA492F9B099",
-25133 => x"C0C0BFA492F9B0B0",
-25132 => x"C0C0BFA492F9B0A4",
-25131 => x"C0C0BFA492F9B0F9",
-25130 => x"C0C0BFA492F9B0C0",
-25129 => x"C0C0BFA492F9A490",
-25128 => x"C0C0BFA492F9A480",
-25127 => x"C0C0BFA492F9A4F8",
-25126 => x"C0C0BFA492F9A482",
-25125 => x"C0C0BFA492F9A492",
-25124 => x"C0C0BFA492F9A499",
-25123 => x"C0C0BFA492F9A4B0",
-25122 => x"C0C0BFA492F9A4A4",
-25121 => x"C0C0BFA492F9A4F9",
-25120 => x"C0C0BFA492F9A4C0",
-25119 => x"C0C0BFA492F9F990",
-25118 => x"C0C0BFA492F9F980",
-25117 => x"C0C0BFA492F9F9F8",
-25116 => x"C0C0BFA492F9F982",
-25115 => x"C0C0BFA492F9F992",
-25114 => x"C0C0BFA492F9F999",
-25113 => x"C0C0BFA492F9F9B0",
-25112 => x"C0C0BFA492F9F9A4",
-25111 => x"C0C0BFA492F9F9F9",
-25110 => x"C0C0BFA492F9F9C0",
-25109 => x"C0C0BFA492F9C090",
-25108 => x"C0C0BFA492F9C080",
-25107 => x"C0C0BFA492F9C0F8",
-25106 => x"C0C0BFA492F9C082",
-25105 => x"C0C0BFA492F9C092",
-25104 => x"C0C0BFA492F9C099",
-25103 => x"C0C0BFA492F9C0B0",
-25102 => x"C0C0BFA492F9C0A4",
-25101 => x"C0C0BFA492F9C0F9",
-25100 => x"C0C0BFA492F9C0C0",
-25099 => x"C0C0BFA492C09090",
-25098 => x"C0C0BFA492C09080",
-25097 => x"C0C0BFA492C090F8",
-25096 => x"C0C0BFA492C09082",
-25095 => x"C0C0BFA492C09092",
-25094 => x"C0C0BFA492C09099",
-25093 => x"C0C0BFA492C090B0",
-25092 => x"C0C0BFA492C090A4",
-25091 => x"C0C0BFA492C090F9",
-25090 => x"C0C0BFA492C090C0",
-25089 => x"C0C0BFA492C08090",
-25088 => x"C0C0BFA492C08080",
-25087 => x"C0C0BFA492C080F8",
-25086 => x"C0C0BFA492C08082",
-25085 => x"C0C0BFA492C08092",
-25084 => x"C0C0BFA492C08099",
-25083 => x"C0C0BFA492C080B0",
-25082 => x"C0C0BFA492C080A4",
-25081 => x"C0C0BFA492C080F9",
-25080 => x"C0C0BFA492C080C0",
-25079 => x"C0C0BFA492C0F890",
-25078 => x"C0C0BFA492C0F880",
-25077 => x"C0C0BFA492C0F8F8",
-25076 => x"C0C0BFA492C0F882",
-25075 => x"C0C0BFA492C0F892",
-25074 => x"C0C0BFA492C0F899",
-25073 => x"C0C0BFA492C0F8B0",
-25072 => x"C0C0BFA492C0F8A4",
-25071 => x"C0C0BFA492C0F8F9",
-25070 => x"C0C0BFA492C0F8C0",
-25069 => x"C0C0BFA492C08290",
-25068 => x"C0C0BFA492C08280",
-25067 => x"C0C0BFA492C082F8",
-25066 => x"C0C0BFA492C08282",
-25065 => x"C0C0BFA492C08292",
-25064 => x"C0C0BFA492C08299",
-25063 => x"C0C0BFA492C082B0",
-25062 => x"C0C0BFA492C082A4",
-25061 => x"C0C0BFA492C082F9",
-25060 => x"C0C0BFA492C082C0",
-25059 => x"C0C0BFA492C09290",
-25058 => x"C0C0BFA492C09280",
-25057 => x"C0C0BFA492C092F8",
-25056 => x"C0C0BFA492C09282",
-25055 => x"C0C0BFA492C09292",
-25054 => x"C0C0BFA492C09299",
-25053 => x"C0C0BFA492C092B0",
-25052 => x"C0C0BFA492C092A4",
-25051 => x"C0C0BFA492C092F9",
-25050 => x"C0C0BFA492C092C0",
-25049 => x"C0C0BFA492C09990",
-25048 => x"C0C0BFA492C09980",
-25047 => x"C0C0BFA492C099F8",
-25046 => x"C0C0BFA492C09982",
-25045 => x"C0C0BFA492C09992",
-25044 => x"C0C0BFA492C09999",
-25043 => x"C0C0BFA492C099B0",
-25042 => x"C0C0BFA492C099A4",
-25041 => x"C0C0BFA492C099F9",
-25040 => x"C0C0BFA492C099C0",
-25039 => x"C0C0BFA492C0B090",
-25038 => x"C0C0BFA492C0B080",
-25037 => x"C0C0BFA492C0B0F8",
-25036 => x"C0C0BFA492C0B082",
-25035 => x"C0C0BFA492C0B092",
-25034 => x"C0C0BFA492C0B099",
-25033 => x"C0C0BFA492C0B0B0",
-25032 => x"C0C0BFA492C0B0A4",
-25031 => x"C0C0BFA492C0B0F9",
-25030 => x"C0C0BFA492C0B0C0",
-25029 => x"C0C0BFA492C0A490",
-25028 => x"C0C0BFA492C0A480",
-25027 => x"C0C0BFA492C0A4F8",
-25026 => x"C0C0BFA492C0A482",
-25025 => x"C0C0BFA492C0A492",
-25024 => x"C0C0BFA492C0A499",
-25023 => x"C0C0BFA492C0A4B0",
-25022 => x"C0C0BFA492C0A4A4",
-25021 => x"C0C0BFA492C0A4F9",
-25020 => x"C0C0BFA492C0A4C0",
-25019 => x"C0C0BFA492C0F990",
-25018 => x"C0C0BFA492C0F980",
-25017 => x"C0C0BFA492C0F9F8",
-25016 => x"C0C0BFA492C0F982",
-25015 => x"C0C0BFA492C0F992",
-25014 => x"C0C0BFA492C0F999",
-25013 => x"C0C0BFA492C0F9B0",
-25012 => x"C0C0BFA492C0F9A4",
-25011 => x"C0C0BFA492C0F9F9",
-25010 => x"C0C0BFA492C0F9C0",
-25009 => x"C0C0BFA492C0C090",
-25008 => x"C0C0BFA492C0C080",
-25007 => x"C0C0BFA492C0C0F8",
-25006 => x"C0C0BFA492C0C082",
-25005 => x"C0C0BFA492C0C092",
-25004 => x"C0C0BFA492C0C099",
-25003 => x"C0C0BFA492C0C0B0",
-25002 => x"C0C0BFA492C0C0A4",
-25001 => x"C0C0BFA492C0C0F9",
-25000 => x"C0C0BFA492C0C0C0",
-24999 => x"C0C0BFA499909090",
-24998 => x"C0C0BFA499909080",
-24997 => x"C0C0BFA4999090F8",
-24996 => x"C0C0BFA499909082",
-24995 => x"C0C0BFA499909092",
-24994 => x"C0C0BFA499909099",
-24993 => x"C0C0BFA4999090B0",
-24992 => x"C0C0BFA4999090A4",
-24991 => x"C0C0BFA4999090F9",
-24990 => x"C0C0BFA4999090C0",
-24989 => x"C0C0BFA499908090",
-24988 => x"C0C0BFA499908080",
-24987 => x"C0C0BFA4999080F8",
-24986 => x"C0C0BFA499908082",
-24985 => x"C0C0BFA499908092",
-24984 => x"C0C0BFA499908099",
-24983 => x"C0C0BFA4999080B0",
-24982 => x"C0C0BFA4999080A4",
-24981 => x"C0C0BFA4999080F9",
-24980 => x"C0C0BFA4999080C0",
-24979 => x"C0C0BFA49990F890",
-24978 => x"C0C0BFA49990F880",
-24977 => x"C0C0BFA49990F8F8",
-24976 => x"C0C0BFA49990F882",
-24975 => x"C0C0BFA49990F892",
-24974 => x"C0C0BFA49990F899",
-24973 => x"C0C0BFA49990F8B0",
-24972 => x"C0C0BFA49990F8A4",
-24971 => x"C0C0BFA49990F8F9",
-24970 => x"C0C0BFA49990F8C0",
-24969 => x"C0C0BFA499908290",
-24968 => x"C0C0BFA499908280",
-24967 => x"C0C0BFA4999082F8",
-24966 => x"C0C0BFA499908282",
-24965 => x"C0C0BFA499908292",
-24964 => x"C0C0BFA499908299",
-24963 => x"C0C0BFA4999082B0",
-24962 => x"C0C0BFA4999082A4",
-24961 => x"C0C0BFA4999082F9",
-24960 => x"C0C0BFA4999082C0",
-24959 => x"C0C0BFA499909290",
-24958 => x"C0C0BFA499909280",
-24957 => x"C0C0BFA4999092F8",
-24956 => x"C0C0BFA499909282",
-24955 => x"C0C0BFA499909292",
-24954 => x"C0C0BFA499909299",
-24953 => x"C0C0BFA4999092B0",
-24952 => x"C0C0BFA4999092A4",
-24951 => x"C0C0BFA4999092F9",
-24950 => x"C0C0BFA4999092C0",
-24949 => x"C0C0BFA499909990",
-24948 => x"C0C0BFA499909980",
-24947 => x"C0C0BFA4999099F8",
-24946 => x"C0C0BFA499909982",
-24945 => x"C0C0BFA499909992",
-24944 => x"C0C0BFA499909999",
-24943 => x"C0C0BFA4999099B0",
-24942 => x"C0C0BFA4999099A4",
-24941 => x"C0C0BFA4999099F9",
-24940 => x"C0C0BFA4999099C0",
-24939 => x"C0C0BFA49990B090",
-24938 => x"C0C0BFA49990B080",
-24937 => x"C0C0BFA49990B0F8",
-24936 => x"C0C0BFA49990B082",
-24935 => x"C0C0BFA49990B092",
-24934 => x"C0C0BFA49990B099",
-24933 => x"C0C0BFA49990B0B0",
-24932 => x"C0C0BFA49990B0A4",
-24931 => x"C0C0BFA49990B0F9",
-24930 => x"C0C0BFA49990B0C0",
-24929 => x"C0C0BFA49990A490",
-24928 => x"C0C0BFA49990A480",
-24927 => x"C0C0BFA49990A4F8",
-24926 => x"C0C0BFA49990A482",
-24925 => x"C0C0BFA49990A492",
-24924 => x"C0C0BFA49990A499",
-24923 => x"C0C0BFA49990A4B0",
-24922 => x"C0C0BFA49990A4A4",
-24921 => x"C0C0BFA49990A4F9",
-24920 => x"C0C0BFA49990A4C0",
-24919 => x"C0C0BFA49990F990",
-24918 => x"C0C0BFA49990F980",
-24917 => x"C0C0BFA49990F9F8",
-24916 => x"C0C0BFA49990F982",
-24915 => x"C0C0BFA49990F992",
-24914 => x"C0C0BFA49990F999",
-24913 => x"C0C0BFA49990F9B0",
-24912 => x"C0C0BFA49990F9A4",
-24911 => x"C0C0BFA49990F9F9",
-24910 => x"C0C0BFA49990F9C0",
-24909 => x"C0C0BFA49990C090",
-24908 => x"C0C0BFA49990C080",
-24907 => x"C0C0BFA49990C0F8",
-24906 => x"C0C0BFA49990C082",
-24905 => x"C0C0BFA49990C092",
-24904 => x"C0C0BFA49990C099",
-24903 => x"C0C0BFA49990C0B0",
-24902 => x"C0C0BFA49990C0A4",
-24901 => x"C0C0BFA49990C0F9",
-24900 => x"C0C0BFA49990C0C0",
-24899 => x"C0C0BFA499809090",
-24898 => x"C0C0BFA499809080",
-24897 => x"C0C0BFA4998090F8",
-24896 => x"C0C0BFA499809082",
-24895 => x"C0C0BFA499809092",
-24894 => x"C0C0BFA499809099",
-24893 => x"C0C0BFA4998090B0",
-24892 => x"C0C0BFA4998090A4",
-24891 => x"C0C0BFA4998090F9",
-24890 => x"C0C0BFA4998090C0",
-24889 => x"C0C0BFA499808090",
-24888 => x"C0C0BFA499808080",
-24887 => x"C0C0BFA4998080F8",
-24886 => x"C0C0BFA499808082",
-24885 => x"C0C0BFA499808092",
-24884 => x"C0C0BFA499808099",
-24883 => x"C0C0BFA4998080B0",
-24882 => x"C0C0BFA4998080A4",
-24881 => x"C0C0BFA4998080F9",
-24880 => x"C0C0BFA4998080C0",
-24879 => x"C0C0BFA49980F890",
-24878 => x"C0C0BFA49980F880",
-24877 => x"C0C0BFA49980F8F8",
-24876 => x"C0C0BFA49980F882",
-24875 => x"C0C0BFA49980F892",
-24874 => x"C0C0BFA49980F899",
-24873 => x"C0C0BFA49980F8B0",
-24872 => x"C0C0BFA49980F8A4",
-24871 => x"C0C0BFA49980F8F9",
-24870 => x"C0C0BFA49980F8C0",
-24869 => x"C0C0BFA499808290",
-24868 => x"C0C0BFA499808280",
-24867 => x"C0C0BFA4998082F8",
-24866 => x"C0C0BFA499808282",
-24865 => x"C0C0BFA499808292",
-24864 => x"C0C0BFA499808299",
-24863 => x"C0C0BFA4998082B0",
-24862 => x"C0C0BFA4998082A4",
-24861 => x"C0C0BFA4998082F9",
-24860 => x"C0C0BFA4998082C0",
-24859 => x"C0C0BFA499809290",
-24858 => x"C0C0BFA499809280",
-24857 => x"C0C0BFA4998092F8",
-24856 => x"C0C0BFA499809282",
-24855 => x"C0C0BFA499809292",
-24854 => x"C0C0BFA499809299",
-24853 => x"C0C0BFA4998092B0",
-24852 => x"C0C0BFA4998092A4",
-24851 => x"C0C0BFA4998092F9",
-24850 => x"C0C0BFA4998092C0",
-24849 => x"C0C0BFA499809990",
-24848 => x"C0C0BFA499809980",
-24847 => x"C0C0BFA4998099F8",
-24846 => x"C0C0BFA499809982",
-24845 => x"C0C0BFA499809992",
-24844 => x"C0C0BFA499809999",
-24843 => x"C0C0BFA4998099B0",
-24842 => x"C0C0BFA4998099A4",
-24841 => x"C0C0BFA4998099F9",
-24840 => x"C0C0BFA4998099C0",
-24839 => x"C0C0BFA49980B090",
-24838 => x"C0C0BFA49980B080",
-24837 => x"C0C0BFA49980B0F8",
-24836 => x"C0C0BFA49980B082",
-24835 => x"C0C0BFA49980B092",
-24834 => x"C0C0BFA49980B099",
-24833 => x"C0C0BFA49980B0B0",
-24832 => x"C0C0BFA49980B0A4",
-24831 => x"C0C0BFA49980B0F9",
-24830 => x"C0C0BFA49980B0C0",
-24829 => x"C0C0BFA49980A490",
-24828 => x"C0C0BFA49980A480",
-24827 => x"C0C0BFA49980A4F8",
-24826 => x"C0C0BFA49980A482",
-24825 => x"C0C0BFA49980A492",
-24824 => x"C0C0BFA49980A499",
-24823 => x"C0C0BFA49980A4B0",
-24822 => x"C0C0BFA49980A4A4",
-24821 => x"C0C0BFA49980A4F9",
-24820 => x"C0C0BFA49980A4C0",
-24819 => x"C0C0BFA49980F990",
-24818 => x"C0C0BFA49980F980",
-24817 => x"C0C0BFA49980F9F8",
-24816 => x"C0C0BFA49980F982",
-24815 => x"C0C0BFA49980F992",
-24814 => x"C0C0BFA49980F999",
-24813 => x"C0C0BFA49980F9B0",
-24812 => x"C0C0BFA49980F9A4",
-24811 => x"C0C0BFA49980F9F9",
-24810 => x"C0C0BFA49980F9C0",
-24809 => x"C0C0BFA49980C090",
-24808 => x"C0C0BFA49980C080",
-24807 => x"C0C0BFA49980C0F8",
-24806 => x"C0C0BFA49980C082",
-24805 => x"C0C0BFA49980C092",
-24804 => x"C0C0BFA49980C099",
-24803 => x"C0C0BFA49980C0B0",
-24802 => x"C0C0BFA49980C0A4",
-24801 => x"C0C0BFA49980C0F9",
-24800 => x"C0C0BFA49980C0C0",
-24799 => x"C0C0BFA499F89090",
-24798 => x"C0C0BFA499F89080",
-24797 => x"C0C0BFA499F890F8",
-24796 => x"C0C0BFA499F89082",
-24795 => x"C0C0BFA499F89092",
-24794 => x"C0C0BFA499F89099",
-24793 => x"C0C0BFA499F890B0",
-24792 => x"C0C0BFA499F890A4",
-24791 => x"C0C0BFA499F890F9",
-24790 => x"C0C0BFA499F890C0",
-24789 => x"C0C0BFA499F88090",
-24788 => x"C0C0BFA499F88080",
-24787 => x"C0C0BFA499F880F8",
-24786 => x"C0C0BFA499F88082",
-24785 => x"C0C0BFA499F88092",
-24784 => x"C0C0BFA499F88099",
-24783 => x"C0C0BFA499F880B0",
-24782 => x"C0C0BFA499F880A4",
-24781 => x"C0C0BFA499F880F9",
-24780 => x"C0C0BFA499F880C0",
-24779 => x"C0C0BFA499F8F890",
-24778 => x"C0C0BFA499F8F880",
-24777 => x"C0C0BFA499F8F8F8",
-24776 => x"C0C0BFA499F8F882",
-24775 => x"C0C0BFA499F8F892",
-24774 => x"C0C0BFA499F8F899",
-24773 => x"C0C0BFA499F8F8B0",
-24772 => x"C0C0BFA499F8F8A4",
-24771 => x"C0C0BFA499F8F8F9",
-24770 => x"C0C0BFA499F8F8C0",
-24769 => x"C0C0BFA499F88290",
-24768 => x"C0C0BFA499F88280",
-24767 => x"C0C0BFA499F882F8",
-24766 => x"C0C0BFA499F88282",
-24765 => x"C0C0BFA499F88292",
-24764 => x"C0C0BFA499F88299",
-24763 => x"C0C0BFA499F882B0",
-24762 => x"C0C0BFA499F882A4",
-24761 => x"C0C0BFA499F882F9",
-24760 => x"C0C0BFA499F882C0",
-24759 => x"C0C0BFA499F89290",
-24758 => x"C0C0BFA499F89280",
-24757 => x"C0C0BFA499F892F8",
-24756 => x"C0C0BFA499F89282",
-24755 => x"C0C0BFA499F89292",
-24754 => x"C0C0BFA499F89299",
-24753 => x"C0C0BFA499F892B0",
-24752 => x"C0C0BFA499F892A4",
-24751 => x"C0C0BFA499F892F9",
-24750 => x"C0C0BFA499F892C0",
-24749 => x"C0C0BFA499F89990",
-24748 => x"C0C0BFA499F89980",
-24747 => x"C0C0BFA499F899F8",
-24746 => x"C0C0BFA499F89982",
-24745 => x"C0C0BFA499F89992",
-24744 => x"C0C0BFA499F89999",
-24743 => x"C0C0BFA499F899B0",
-24742 => x"C0C0BFA499F899A4",
-24741 => x"C0C0BFA499F899F9",
-24740 => x"C0C0BFA499F899C0",
-24739 => x"C0C0BFA499F8B090",
-24738 => x"C0C0BFA499F8B080",
-24737 => x"C0C0BFA499F8B0F8",
-24736 => x"C0C0BFA499F8B082",
-24735 => x"C0C0BFA499F8B092",
-24734 => x"C0C0BFA499F8B099",
-24733 => x"C0C0BFA499F8B0B0",
-24732 => x"C0C0BFA499F8B0A4",
-24731 => x"C0C0BFA499F8B0F9",
-24730 => x"C0C0BFA499F8B0C0",
-24729 => x"C0C0BFA499F8A490",
-24728 => x"C0C0BFA499F8A480",
-24727 => x"C0C0BFA499F8A4F8",
-24726 => x"C0C0BFA499F8A482",
-24725 => x"C0C0BFA499F8A492",
-24724 => x"C0C0BFA499F8A499",
-24723 => x"C0C0BFA499F8A4B0",
-24722 => x"C0C0BFA499F8A4A4",
-24721 => x"C0C0BFA499F8A4F9",
-24720 => x"C0C0BFA499F8A4C0",
-24719 => x"C0C0BFA499F8F990",
-24718 => x"C0C0BFA499F8F980",
-24717 => x"C0C0BFA499F8F9F8",
-24716 => x"C0C0BFA499F8F982",
-24715 => x"C0C0BFA499F8F992",
-24714 => x"C0C0BFA499F8F999",
-24713 => x"C0C0BFA499F8F9B0",
-24712 => x"C0C0BFA499F8F9A4",
-24711 => x"C0C0BFA499F8F9F9",
-24710 => x"C0C0BFA499F8F9C0",
-24709 => x"C0C0BFA499F8C090",
-24708 => x"C0C0BFA499F8C080",
-24707 => x"C0C0BFA499F8C0F8",
-24706 => x"C0C0BFA499F8C082",
-24705 => x"C0C0BFA499F8C092",
-24704 => x"C0C0BFA499F8C099",
-24703 => x"C0C0BFA499F8C0B0",
-24702 => x"C0C0BFA499F8C0A4",
-24701 => x"C0C0BFA499F8C0F9",
-24700 => x"C0C0BFA499F8C0C0",
-24699 => x"C0C0BFA499829090",
-24698 => x"C0C0BFA499829080",
-24697 => x"C0C0BFA4998290F8",
-24696 => x"C0C0BFA499829082",
-24695 => x"C0C0BFA499829092",
-24694 => x"C0C0BFA499829099",
-24693 => x"C0C0BFA4998290B0",
-24692 => x"C0C0BFA4998290A4",
-24691 => x"C0C0BFA4998290F9",
-24690 => x"C0C0BFA4998290C0",
-24689 => x"C0C0BFA499828090",
-24688 => x"C0C0BFA499828080",
-24687 => x"C0C0BFA4998280F8",
-24686 => x"C0C0BFA499828082",
-24685 => x"C0C0BFA499828092",
-24684 => x"C0C0BFA499828099",
-24683 => x"C0C0BFA4998280B0",
-24682 => x"C0C0BFA4998280A4",
-24681 => x"C0C0BFA4998280F9",
-24680 => x"C0C0BFA4998280C0",
-24679 => x"C0C0BFA49982F890",
-24678 => x"C0C0BFA49982F880",
-24677 => x"C0C0BFA49982F8F8",
-24676 => x"C0C0BFA49982F882",
-24675 => x"C0C0BFA49982F892",
-24674 => x"C0C0BFA49982F899",
-24673 => x"C0C0BFA49982F8B0",
-24672 => x"C0C0BFA49982F8A4",
-24671 => x"C0C0BFA49982F8F9",
-24670 => x"C0C0BFA49982F8C0",
-24669 => x"C0C0BFA499828290",
-24668 => x"C0C0BFA499828280",
-24667 => x"C0C0BFA4998282F8",
-24666 => x"C0C0BFA499828282",
-24665 => x"C0C0BFA499828292",
-24664 => x"C0C0BFA499828299",
-24663 => x"C0C0BFA4998282B0",
-24662 => x"C0C0BFA4998282A4",
-24661 => x"C0C0BFA4998282F9",
-24660 => x"C0C0BFA4998282C0",
-24659 => x"C0C0BFA499829290",
-24658 => x"C0C0BFA499829280",
-24657 => x"C0C0BFA4998292F8",
-24656 => x"C0C0BFA499829282",
-24655 => x"C0C0BFA499829292",
-24654 => x"C0C0BFA499829299",
-24653 => x"C0C0BFA4998292B0",
-24652 => x"C0C0BFA4998292A4",
-24651 => x"C0C0BFA4998292F9",
-24650 => x"C0C0BFA4998292C0",
-24649 => x"C0C0BFA499829990",
-24648 => x"C0C0BFA499829980",
-24647 => x"C0C0BFA4998299F8",
-24646 => x"C0C0BFA499829982",
-24645 => x"C0C0BFA499829992",
-24644 => x"C0C0BFA499829999",
-24643 => x"C0C0BFA4998299B0",
-24642 => x"C0C0BFA4998299A4",
-24641 => x"C0C0BFA4998299F9",
-24640 => x"C0C0BFA4998299C0",
-24639 => x"C0C0BFA49982B090",
-24638 => x"C0C0BFA49982B080",
-24637 => x"C0C0BFA49982B0F8",
-24636 => x"C0C0BFA49982B082",
-24635 => x"C0C0BFA49982B092",
-24634 => x"C0C0BFA49982B099",
-24633 => x"C0C0BFA49982B0B0",
-24632 => x"C0C0BFA49982B0A4",
-24631 => x"C0C0BFA49982B0F9",
-24630 => x"C0C0BFA49982B0C0",
-24629 => x"C0C0BFA49982A490",
-24628 => x"C0C0BFA49982A480",
-24627 => x"C0C0BFA49982A4F8",
-24626 => x"C0C0BFA49982A482",
-24625 => x"C0C0BFA49982A492",
-24624 => x"C0C0BFA49982A499",
-24623 => x"C0C0BFA49982A4B0",
-24622 => x"C0C0BFA49982A4A4",
-24621 => x"C0C0BFA49982A4F9",
-24620 => x"C0C0BFA49982A4C0",
-24619 => x"C0C0BFA49982F990",
-24618 => x"C0C0BFA49982F980",
-24617 => x"C0C0BFA49982F9F8",
-24616 => x"C0C0BFA49982F982",
-24615 => x"C0C0BFA49982F992",
-24614 => x"C0C0BFA49982F999",
-24613 => x"C0C0BFA49982F9B0",
-24612 => x"C0C0BFA49982F9A4",
-24611 => x"C0C0BFA49982F9F9",
-24610 => x"C0C0BFA49982F9C0",
-24609 => x"C0C0BFA49982C090",
-24608 => x"C0C0BFA49982C080",
-24607 => x"C0C0BFA49982C0F8",
-24606 => x"C0C0BFA49982C082",
-24605 => x"C0C0BFA49982C092",
-24604 => x"C0C0BFA49982C099",
-24603 => x"C0C0BFA49982C0B0",
-24602 => x"C0C0BFA49982C0A4",
-24601 => x"C0C0BFA49982C0F9",
-24600 => x"C0C0BFA49982C0C0",
-24599 => x"C0C0BFA499929090",
-24598 => x"C0C0BFA499929080",
-24597 => x"C0C0BFA4999290F8",
-24596 => x"C0C0BFA499929082",
-24595 => x"C0C0BFA499929092",
-24594 => x"C0C0BFA499929099",
-24593 => x"C0C0BFA4999290B0",
-24592 => x"C0C0BFA4999290A4",
-24591 => x"C0C0BFA4999290F9",
-24590 => x"C0C0BFA4999290C0",
-24589 => x"C0C0BFA499928090",
-24588 => x"C0C0BFA499928080",
-24587 => x"C0C0BFA4999280F8",
-24586 => x"C0C0BFA499928082",
-24585 => x"C0C0BFA499928092",
-24584 => x"C0C0BFA499928099",
-24583 => x"C0C0BFA4999280B0",
-24582 => x"C0C0BFA4999280A4",
-24581 => x"C0C0BFA4999280F9",
-24580 => x"C0C0BFA4999280C0",
-24579 => x"C0C0BFA49992F890",
-24578 => x"C0C0BFA49992F880",
-24577 => x"C0C0BFA49992F8F8",
-24576 => x"C0C0BFA49992F882",
-24575 => x"C0C0BFA49992F892",
-24574 => x"C0C0BFA49992F899",
-24573 => x"C0C0BFA49992F8B0",
-24572 => x"C0C0BFA49992F8A4",
-24571 => x"C0C0BFA49992F8F9",
-24570 => x"C0C0BFA49992F8C0",
-24569 => x"C0C0BFA499928290",
-24568 => x"C0C0BFA499928280",
-24567 => x"C0C0BFA4999282F8",
-24566 => x"C0C0BFA499928282",
-24565 => x"C0C0BFA499928292",
-24564 => x"C0C0BFA499928299",
-24563 => x"C0C0BFA4999282B0",
-24562 => x"C0C0BFA4999282A4",
-24561 => x"C0C0BFA4999282F9",
-24560 => x"C0C0BFA4999282C0",
-24559 => x"C0C0BFA499929290",
-24558 => x"C0C0BFA499929280",
-24557 => x"C0C0BFA4999292F8",
-24556 => x"C0C0BFA499929282",
-24555 => x"C0C0BFA499929292",
-24554 => x"C0C0BFA499929299",
-24553 => x"C0C0BFA4999292B0",
-24552 => x"C0C0BFA4999292A4",
-24551 => x"C0C0BFA4999292F9",
-24550 => x"C0C0BFA4999292C0",
-24549 => x"C0C0BFA499929990",
-24548 => x"C0C0BFA499929980",
-24547 => x"C0C0BFA4999299F8",
-24546 => x"C0C0BFA499929982",
-24545 => x"C0C0BFA499929992",
-24544 => x"C0C0BFA499929999",
-24543 => x"C0C0BFA4999299B0",
-24542 => x"C0C0BFA4999299A4",
-24541 => x"C0C0BFA4999299F9",
-24540 => x"C0C0BFA4999299C0",
-24539 => x"C0C0BFA49992B090",
-24538 => x"C0C0BFA49992B080",
-24537 => x"C0C0BFA49992B0F8",
-24536 => x"C0C0BFA49992B082",
-24535 => x"C0C0BFA49992B092",
-24534 => x"C0C0BFA49992B099",
-24533 => x"C0C0BFA49992B0B0",
-24532 => x"C0C0BFA49992B0A4",
-24531 => x"C0C0BFA49992B0F9",
-24530 => x"C0C0BFA49992B0C0",
-24529 => x"C0C0BFA49992A490",
-24528 => x"C0C0BFA49992A480",
-24527 => x"C0C0BFA49992A4F8",
-24526 => x"C0C0BFA49992A482",
-24525 => x"C0C0BFA49992A492",
-24524 => x"C0C0BFA49992A499",
-24523 => x"C0C0BFA49992A4B0",
-24522 => x"C0C0BFA49992A4A4",
-24521 => x"C0C0BFA49992A4F9",
-24520 => x"C0C0BFA49992A4C0",
-24519 => x"C0C0BFA49992F990",
-24518 => x"C0C0BFA49992F980",
-24517 => x"C0C0BFA49992F9F8",
-24516 => x"C0C0BFA49992F982",
-24515 => x"C0C0BFA49992F992",
-24514 => x"C0C0BFA49992F999",
-24513 => x"C0C0BFA49992F9B0",
-24512 => x"C0C0BFA49992F9A4",
-24511 => x"C0C0BFA49992F9F9",
-24510 => x"C0C0BFA49992F9C0",
-24509 => x"C0C0BFA49992C090",
-24508 => x"C0C0BFA49992C080",
-24507 => x"C0C0BFA49992C0F8",
-24506 => x"C0C0BFA49992C082",
-24505 => x"C0C0BFA49992C092",
-24504 => x"C0C0BFA49992C099",
-24503 => x"C0C0BFA49992C0B0",
-24502 => x"C0C0BFA49992C0A4",
-24501 => x"C0C0BFA49992C0F9",
-24500 => x"C0C0BFA49992C0C0",
-24499 => x"C0C0BFA499999090",
-24498 => x"C0C0BFA499999080",
-24497 => x"C0C0BFA4999990F8",
-24496 => x"C0C0BFA499999082",
-24495 => x"C0C0BFA499999092",
-24494 => x"C0C0BFA499999099",
-24493 => x"C0C0BFA4999990B0",
-24492 => x"C0C0BFA4999990A4",
-24491 => x"C0C0BFA4999990F9",
-24490 => x"C0C0BFA4999990C0",
-24489 => x"C0C0BFA499998090",
-24488 => x"C0C0BFA499998080",
-24487 => x"C0C0BFA4999980F8",
-24486 => x"C0C0BFA499998082",
-24485 => x"C0C0BFA499998092",
-24484 => x"C0C0BFA499998099",
-24483 => x"C0C0BFA4999980B0",
-24482 => x"C0C0BFA4999980A4",
-24481 => x"C0C0BFA4999980F9",
-24480 => x"C0C0BFA4999980C0",
-24479 => x"C0C0BFA49999F890",
-24478 => x"C0C0BFA49999F880",
-24477 => x"C0C0BFA49999F8F8",
-24476 => x"C0C0BFA49999F882",
-24475 => x"C0C0BFA49999F892",
-24474 => x"C0C0BFA49999F899",
-24473 => x"C0C0BFA49999F8B0",
-24472 => x"C0C0BFA49999F8A4",
-24471 => x"C0C0BFA49999F8F9",
-24470 => x"C0C0BFA49999F8C0",
-24469 => x"C0C0BFA499998290",
-24468 => x"C0C0BFA499998280",
-24467 => x"C0C0BFA4999982F8",
-24466 => x"C0C0BFA499998282",
-24465 => x"C0C0BFA499998292",
-24464 => x"C0C0BFA499998299",
-24463 => x"C0C0BFA4999982B0",
-24462 => x"C0C0BFA4999982A4",
-24461 => x"C0C0BFA4999982F9",
-24460 => x"C0C0BFA4999982C0",
-24459 => x"C0C0BFA499999290",
-24458 => x"C0C0BFA499999280",
-24457 => x"C0C0BFA4999992F8",
-24456 => x"C0C0BFA499999282",
-24455 => x"C0C0BFA499999292",
-24454 => x"C0C0BFA499999299",
-24453 => x"C0C0BFA4999992B0",
-24452 => x"C0C0BFA4999992A4",
-24451 => x"C0C0BFA4999992F9",
-24450 => x"C0C0BFA4999992C0",
-24449 => x"C0C0BFA499999990",
-24448 => x"C0C0BFA499999980",
-24447 => x"C0C0BFA4999999F8",
-24446 => x"C0C0BFA499999982",
-24445 => x"C0C0BFA499999992",
-24444 => x"C0C0BFA499999999",
-24443 => x"C0C0BFA4999999B0",
-24442 => x"C0C0BFA4999999A4",
-24441 => x"C0C0BFA4999999F9",
-24440 => x"C0C0BFA4999999C0",
-24439 => x"C0C0BFA49999B090",
-24438 => x"C0C0BFA49999B080",
-24437 => x"C0C0BFA49999B0F8",
-24436 => x"C0C0BFA49999B082",
-24435 => x"C0C0BFA49999B092",
-24434 => x"C0C0BFA49999B099",
-24433 => x"C0C0BFA49999B0B0",
-24432 => x"C0C0BFA49999B0A4",
-24431 => x"C0C0BFA49999B0F9",
-24430 => x"C0C0BFA49999B0C0",
-24429 => x"C0C0BFA49999A490",
-24428 => x"C0C0BFA49999A480",
-24427 => x"C0C0BFA49999A4F8",
-24426 => x"C0C0BFA49999A482",
-24425 => x"C0C0BFA49999A492",
-24424 => x"C0C0BFA49999A499",
-24423 => x"C0C0BFA49999A4B0",
-24422 => x"C0C0BFA49999A4A4",
-24421 => x"C0C0BFA49999A4F9",
-24420 => x"C0C0BFA49999A4C0",
-24419 => x"C0C0BFA49999F990",
-24418 => x"C0C0BFA49999F980",
-24417 => x"C0C0BFA49999F9F8",
-24416 => x"C0C0BFA49999F982",
-24415 => x"C0C0BFA49999F992",
-24414 => x"C0C0BFA49999F999",
-24413 => x"C0C0BFA49999F9B0",
-24412 => x"C0C0BFA49999F9A4",
-24411 => x"C0C0BFA49999F9F9",
-24410 => x"C0C0BFA49999F9C0",
-24409 => x"C0C0BFA49999C090",
-24408 => x"C0C0BFA49999C080",
-24407 => x"C0C0BFA49999C0F8",
-24406 => x"C0C0BFA49999C082",
-24405 => x"C0C0BFA49999C092",
-24404 => x"C0C0BFA49999C099",
-24403 => x"C0C0BFA49999C0B0",
-24402 => x"C0C0BFA49999C0A4",
-24401 => x"C0C0BFA49999C0F9",
-24400 => x"C0C0BFA49999C0C0",
-24399 => x"C0C0BFA499B09090",
-24398 => x"C0C0BFA499B09080",
-24397 => x"C0C0BFA499B090F8",
-24396 => x"C0C0BFA499B09082",
-24395 => x"C0C0BFA499B09092",
-24394 => x"C0C0BFA499B09099",
-24393 => x"C0C0BFA499B090B0",
-24392 => x"C0C0BFA499B090A4",
-24391 => x"C0C0BFA499B090F9",
-24390 => x"C0C0BFA499B090C0",
-24389 => x"C0C0BFA499B08090",
-24388 => x"C0C0BFA499B08080",
-24387 => x"C0C0BFA499B080F8",
-24386 => x"C0C0BFA499B08082",
-24385 => x"C0C0BFA499B08092",
-24384 => x"C0C0BFA499B08099",
-24383 => x"C0C0BFA499B080B0",
-24382 => x"C0C0BFA499B080A4",
-24381 => x"C0C0BFA499B080F9",
-24380 => x"C0C0BFA499B080C0",
-24379 => x"C0C0BFA499B0F890",
-24378 => x"C0C0BFA499B0F880",
-24377 => x"C0C0BFA499B0F8F8",
-24376 => x"C0C0BFA499B0F882",
-24375 => x"C0C0BFA499B0F892",
-24374 => x"C0C0BFA499B0F899",
-24373 => x"C0C0BFA499B0F8B0",
-24372 => x"C0C0BFA499B0F8A4",
-24371 => x"C0C0BFA499B0F8F9",
-24370 => x"C0C0BFA499B0F8C0",
-24369 => x"C0C0BFA499B08290",
-24368 => x"C0C0BFA499B08280",
-24367 => x"C0C0BFA499B082F8",
-24366 => x"C0C0BFA499B08282",
-24365 => x"C0C0BFA499B08292",
-24364 => x"C0C0BFA499B08299",
-24363 => x"C0C0BFA499B082B0",
-24362 => x"C0C0BFA499B082A4",
-24361 => x"C0C0BFA499B082F9",
-24360 => x"C0C0BFA499B082C0",
-24359 => x"C0C0BFA499B09290",
-24358 => x"C0C0BFA499B09280",
-24357 => x"C0C0BFA499B092F8",
-24356 => x"C0C0BFA499B09282",
-24355 => x"C0C0BFA499B09292",
-24354 => x"C0C0BFA499B09299",
-24353 => x"C0C0BFA499B092B0",
-24352 => x"C0C0BFA499B092A4",
-24351 => x"C0C0BFA499B092F9",
-24350 => x"C0C0BFA499B092C0",
-24349 => x"C0C0BFA499B09990",
-24348 => x"C0C0BFA499B09980",
-24347 => x"C0C0BFA499B099F8",
-24346 => x"C0C0BFA499B09982",
-24345 => x"C0C0BFA499B09992",
-24344 => x"C0C0BFA499B09999",
-24343 => x"C0C0BFA499B099B0",
-24342 => x"C0C0BFA499B099A4",
-24341 => x"C0C0BFA499B099F9",
-24340 => x"C0C0BFA499B099C0",
-24339 => x"C0C0BFA499B0B090",
-24338 => x"C0C0BFA499B0B080",
-24337 => x"C0C0BFA499B0B0F8",
-24336 => x"C0C0BFA499B0B082",
-24335 => x"C0C0BFA499B0B092",
-24334 => x"C0C0BFA499B0B099",
-24333 => x"C0C0BFA499B0B0B0",
-24332 => x"C0C0BFA499B0B0A4",
-24331 => x"C0C0BFA499B0B0F9",
-24330 => x"C0C0BFA499B0B0C0",
-24329 => x"C0C0BFA499B0A490",
-24328 => x"C0C0BFA499B0A480",
-24327 => x"C0C0BFA499B0A4F8",
-24326 => x"C0C0BFA499B0A482",
-24325 => x"C0C0BFA499B0A492",
-24324 => x"C0C0BFA499B0A499",
-24323 => x"C0C0BFA499B0A4B0",
-24322 => x"C0C0BFA499B0A4A4",
-24321 => x"C0C0BFA499B0A4F9",
-24320 => x"C0C0BFA499B0A4C0",
-24319 => x"C0C0BFA499B0F990",
-24318 => x"C0C0BFA499B0F980",
-24317 => x"C0C0BFA499B0F9F8",
-24316 => x"C0C0BFA499B0F982",
-24315 => x"C0C0BFA499B0F992",
-24314 => x"C0C0BFA499B0F999",
-24313 => x"C0C0BFA499B0F9B0",
-24312 => x"C0C0BFA499B0F9A4",
-24311 => x"C0C0BFA499B0F9F9",
-24310 => x"C0C0BFA499B0F9C0",
-24309 => x"C0C0BFA499B0C090",
-24308 => x"C0C0BFA499B0C080",
-24307 => x"C0C0BFA499B0C0F8",
-24306 => x"C0C0BFA499B0C082",
-24305 => x"C0C0BFA499B0C092",
-24304 => x"C0C0BFA499B0C099",
-24303 => x"C0C0BFA499B0C0B0",
-24302 => x"C0C0BFA499B0C0A4",
-24301 => x"C0C0BFA499B0C0F9",
-24300 => x"C0C0BFA499B0C0C0",
-24299 => x"C0C0BFA499A49090",
-24298 => x"C0C0BFA499A49080",
-24297 => x"C0C0BFA499A490F8",
-24296 => x"C0C0BFA499A49082",
-24295 => x"C0C0BFA499A49092",
-24294 => x"C0C0BFA499A49099",
-24293 => x"C0C0BFA499A490B0",
-24292 => x"C0C0BFA499A490A4",
-24291 => x"C0C0BFA499A490F9",
-24290 => x"C0C0BFA499A490C0",
-24289 => x"C0C0BFA499A48090",
-24288 => x"C0C0BFA499A48080",
-24287 => x"C0C0BFA499A480F8",
-24286 => x"C0C0BFA499A48082",
-24285 => x"C0C0BFA499A48092",
-24284 => x"C0C0BFA499A48099",
-24283 => x"C0C0BFA499A480B0",
-24282 => x"C0C0BFA499A480A4",
-24281 => x"C0C0BFA499A480F9",
-24280 => x"C0C0BFA499A480C0",
-24279 => x"C0C0BFA499A4F890",
-24278 => x"C0C0BFA499A4F880",
-24277 => x"C0C0BFA499A4F8F8",
-24276 => x"C0C0BFA499A4F882",
-24275 => x"C0C0BFA499A4F892",
-24274 => x"C0C0BFA499A4F899",
-24273 => x"C0C0BFA499A4F8B0",
-24272 => x"C0C0BFA499A4F8A4",
-24271 => x"C0C0BFA499A4F8F9",
-24270 => x"C0C0BFA499A4F8C0",
-24269 => x"C0C0BFA499A48290",
-24268 => x"C0C0BFA499A48280",
-24267 => x"C0C0BFA499A482F8",
-24266 => x"C0C0BFA499A48282",
-24265 => x"C0C0BFA499A48292",
-24264 => x"C0C0BFA499A48299",
-24263 => x"C0C0BFA499A482B0",
-24262 => x"C0C0BFA499A482A4",
-24261 => x"C0C0BFA499A482F9",
-24260 => x"C0C0BFA499A482C0",
-24259 => x"C0C0BFA499A49290",
-24258 => x"C0C0BFA499A49280",
-24257 => x"C0C0BFA499A492F8",
-24256 => x"C0C0BFA499A49282",
-24255 => x"C0C0BFA499A49292",
-24254 => x"C0C0BFA499A49299",
-24253 => x"C0C0BFA499A492B0",
-24252 => x"C0C0BFA499A492A4",
-24251 => x"C0C0BFA499A492F9",
-24250 => x"C0C0BFA499A492C0",
-24249 => x"C0C0BFA499A49990",
-24248 => x"C0C0BFA499A49980",
-24247 => x"C0C0BFA499A499F8",
-24246 => x"C0C0BFA499A49982",
-24245 => x"C0C0BFA499A49992",
-24244 => x"C0C0BFA499A49999",
-24243 => x"C0C0BFA499A499B0",
-24242 => x"C0C0BFA499A499A4",
-24241 => x"C0C0BFA499A499F9",
-24240 => x"C0C0BFA499A499C0",
-24239 => x"C0C0BFA499A4B090",
-24238 => x"C0C0BFA499A4B080",
-24237 => x"C0C0BFA499A4B0F8",
-24236 => x"C0C0BFA499A4B082",
-24235 => x"C0C0BFA499A4B092",
-24234 => x"C0C0BFA499A4B099",
-24233 => x"C0C0BFA499A4B0B0",
-24232 => x"C0C0BFA499A4B0A4",
-24231 => x"C0C0BFA499A4B0F9",
-24230 => x"C0C0BFA499A4B0C0",
-24229 => x"C0C0BFA499A4A490",
-24228 => x"C0C0BFA499A4A480",
-24227 => x"C0C0BFA499A4A4F8",
-24226 => x"C0C0BFA499A4A482",
-24225 => x"C0C0BFA499A4A492",
-24224 => x"C0C0BFA499A4A499",
-24223 => x"C0C0BFA499A4A4B0",
-24222 => x"C0C0BFA499A4A4A4",
-24221 => x"C0C0BFA499A4A4F9",
-24220 => x"C0C0BFA499A4A4C0",
-24219 => x"C0C0BFA499A4F990",
-24218 => x"C0C0BFA499A4F980",
-24217 => x"C0C0BFA499A4F9F8",
-24216 => x"C0C0BFA499A4F982",
-24215 => x"C0C0BFA499A4F992",
-24214 => x"C0C0BFA499A4F999",
-24213 => x"C0C0BFA499A4F9B0",
-24212 => x"C0C0BFA499A4F9A4",
-24211 => x"C0C0BFA499A4F9F9",
-24210 => x"C0C0BFA499A4F9C0",
-24209 => x"C0C0BFA499A4C090",
-24208 => x"C0C0BFA499A4C080",
-24207 => x"C0C0BFA499A4C0F8",
-24206 => x"C0C0BFA499A4C082",
-24205 => x"C0C0BFA499A4C092",
-24204 => x"C0C0BFA499A4C099",
-24203 => x"C0C0BFA499A4C0B0",
-24202 => x"C0C0BFA499A4C0A4",
-24201 => x"C0C0BFA499A4C0F9",
-24200 => x"C0C0BFA499A4C0C0",
-24199 => x"C0C0BFA499F99090",
-24198 => x"C0C0BFA499F99080",
-24197 => x"C0C0BFA499F990F8",
-24196 => x"C0C0BFA499F99082",
-24195 => x"C0C0BFA499F99092",
-24194 => x"C0C0BFA499F99099",
-24193 => x"C0C0BFA499F990B0",
-24192 => x"C0C0BFA499F990A4",
-24191 => x"C0C0BFA499F990F9",
-24190 => x"C0C0BFA499F990C0",
-24189 => x"C0C0BFA499F98090",
-24188 => x"C0C0BFA499F98080",
-24187 => x"C0C0BFA499F980F8",
-24186 => x"C0C0BFA499F98082",
-24185 => x"C0C0BFA499F98092",
-24184 => x"C0C0BFA499F98099",
-24183 => x"C0C0BFA499F980B0",
-24182 => x"C0C0BFA499F980A4",
-24181 => x"C0C0BFA499F980F9",
-24180 => x"C0C0BFA499F980C0",
-24179 => x"C0C0BFA499F9F890",
-24178 => x"C0C0BFA499F9F880",
-24177 => x"C0C0BFA499F9F8F8",
-24176 => x"C0C0BFA499F9F882",
-24175 => x"C0C0BFA499F9F892",
-24174 => x"C0C0BFA499F9F899",
-24173 => x"C0C0BFA499F9F8B0",
-24172 => x"C0C0BFA499F9F8A4",
-24171 => x"C0C0BFA499F9F8F9",
-24170 => x"C0C0BFA499F9F8C0",
-24169 => x"C0C0BFA499F98290",
-24168 => x"C0C0BFA499F98280",
-24167 => x"C0C0BFA499F982F8",
-24166 => x"C0C0BFA499F98282",
-24165 => x"C0C0BFA499F98292",
-24164 => x"C0C0BFA499F98299",
-24163 => x"C0C0BFA499F982B0",
-24162 => x"C0C0BFA499F982A4",
-24161 => x"C0C0BFA499F982F9",
-24160 => x"C0C0BFA499F982C0",
-24159 => x"C0C0BFA499F99290",
-24158 => x"C0C0BFA499F99280",
-24157 => x"C0C0BFA499F992F8",
-24156 => x"C0C0BFA499F99282",
-24155 => x"C0C0BFA499F99292",
-24154 => x"C0C0BFA499F99299",
-24153 => x"C0C0BFA499F992B0",
-24152 => x"C0C0BFA499F992A4",
-24151 => x"C0C0BFA499F992F9",
-24150 => x"C0C0BFA499F992C0",
-24149 => x"C0C0BFA499F99990",
-24148 => x"C0C0BFA499F99980",
-24147 => x"C0C0BFA499F999F8",
-24146 => x"C0C0BFA499F99982",
-24145 => x"C0C0BFA499F99992",
-24144 => x"C0C0BFA499F99999",
-24143 => x"C0C0BFA499F999B0",
-24142 => x"C0C0BFA499F999A4",
-24141 => x"C0C0BFA499F999F9",
-24140 => x"C0C0BFA499F999C0",
-24139 => x"C0C0BFA499F9B090",
-24138 => x"C0C0BFA499F9B080",
-24137 => x"C0C0BFA499F9B0F8",
-24136 => x"C0C0BFA499F9B082",
-24135 => x"C0C0BFA499F9B092",
-24134 => x"C0C0BFA499F9B099",
-24133 => x"C0C0BFA499F9B0B0",
-24132 => x"C0C0BFA499F9B0A4",
-24131 => x"C0C0BFA499F9B0F9",
-24130 => x"C0C0BFA499F9B0C0",
-24129 => x"C0C0BFA499F9A490",
-24128 => x"C0C0BFA499F9A480",
-24127 => x"C0C0BFA499F9A4F8",
-24126 => x"C0C0BFA499F9A482",
-24125 => x"C0C0BFA499F9A492",
-24124 => x"C0C0BFA499F9A499",
-24123 => x"C0C0BFA499F9A4B0",
-24122 => x"C0C0BFA499F9A4A4",
-24121 => x"C0C0BFA499F9A4F9",
-24120 => x"C0C0BFA499F9A4C0",
-24119 => x"C0C0BFA499F9F990",
-24118 => x"C0C0BFA499F9F980",
-24117 => x"C0C0BFA499F9F9F8",
-24116 => x"C0C0BFA499F9F982",
-24115 => x"C0C0BFA499F9F992",
-24114 => x"C0C0BFA499F9F999",
-24113 => x"C0C0BFA499F9F9B0",
-24112 => x"C0C0BFA499F9F9A4",
-24111 => x"C0C0BFA499F9F9F9",
-24110 => x"C0C0BFA499F9F9C0",
-24109 => x"C0C0BFA499F9C090",
-24108 => x"C0C0BFA499F9C080",
-24107 => x"C0C0BFA499F9C0F8",
-24106 => x"C0C0BFA499F9C082",
-24105 => x"C0C0BFA499F9C092",
-24104 => x"C0C0BFA499F9C099",
-24103 => x"C0C0BFA499F9C0B0",
-24102 => x"C0C0BFA499F9C0A4",
-24101 => x"C0C0BFA499F9C0F9",
-24100 => x"C0C0BFA499F9C0C0",
-24099 => x"C0C0BFA499C09090",
-24098 => x"C0C0BFA499C09080",
-24097 => x"C0C0BFA499C090F8",
-24096 => x"C0C0BFA499C09082",
-24095 => x"C0C0BFA499C09092",
-24094 => x"C0C0BFA499C09099",
-24093 => x"C0C0BFA499C090B0",
-24092 => x"C0C0BFA499C090A4",
-24091 => x"C0C0BFA499C090F9",
-24090 => x"C0C0BFA499C090C0",
-24089 => x"C0C0BFA499C08090",
-24088 => x"C0C0BFA499C08080",
-24087 => x"C0C0BFA499C080F8",
-24086 => x"C0C0BFA499C08082",
-24085 => x"C0C0BFA499C08092",
-24084 => x"C0C0BFA499C08099",
-24083 => x"C0C0BFA499C080B0",
-24082 => x"C0C0BFA499C080A4",
-24081 => x"C0C0BFA499C080F9",
-24080 => x"C0C0BFA499C080C0",
-24079 => x"C0C0BFA499C0F890",
-24078 => x"C0C0BFA499C0F880",
-24077 => x"C0C0BFA499C0F8F8",
-24076 => x"C0C0BFA499C0F882",
-24075 => x"C0C0BFA499C0F892",
-24074 => x"C0C0BFA499C0F899",
-24073 => x"C0C0BFA499C0F8B0",
-24072 => x"C0C0BFA499C0F8A4",
-24071 => x"C0C0BFA499C0F8F9",
-24070 => x"C0C0BFA499C0F8C0",
-24069 => x"C0C0BFA499C08290",
-24068 => x"C0C0BFA499C08280",
-24067 => x"C0C0BFA499C082F8",
-24066 => x"C0C0BFA499C08282",
-24065 => x"C0C0BFA499C08292",
-24064 => x"C0C0BFA499C08299",
-24063 => x"C0C0BFA499C082B0",
-24062 => x"C0C0BFA499C082A4",
-24061 => x"C0C0BFA499C082F9",
-24060 => x"C0C0BFA499C082C0",
-24059 => x"C0C0BFA499C09290",
-24058 => x"C0C0BFA499C09280",
-24057 => x"C0C0BFA499C092F8",
-24056 => x"C0C0BFA499C09282",
-24055 => x"C0C0BFA499C09292",
-24054 => x"C0C0BFA499C09299",
-24053 => x"C0C0BFA499C092B0",
-24052 => x"C0C0BFA499C092A4",
-24051 => x"C0C0BFA499C092F9",
-24050 => x"C0C0BFA499C092C0",
-24049 => x"C0C0BFA499C09990",
-24048 => x"C0C0BFA499C09980",
-24047 => x"C0C0BFA499C099F8",
-24046 => x"C0C0BFA499C09982",
-24045 => x"C0C0BFA499C09992",
-24044 => x"C0C0BFA499C09999",
-24043 => x"C0C0BFA499C099B0",
-24042 => x"C0C0BFA499C099A4",
-24041 => x"C0C0BFA499C099F9",
-24040 => x"C0C0BFA499C099C0",
-24039 => x"C0C0BFA499C0B090",
-24038 => x"C0C0BFA499C0B080",
-24037 => x"C0C0BFA499C0B0F8",
-24036 => x"C0C0BFA499C0B082",
-24035 => x"C0C0BFA499C0B092",
-24034 => x"C0C0BFA499C0B099",
-24033 => x"C0C0BFA499C0B0B0",
-24032 => x"C0C0BFA499C0B0A4",
-24031 => x"C0C0BFA499C0B0F9",
-24030 => x"C0C0BFA499C0B0C0",
-24029 => x"C0C0BFA499C0A490",
-24028 => x"C0C0BFA499C0A480",
-24027 => x"C0C0BFA499C0A4F8",
-24026 => x"C0C0BFA499C0A482",
-24025 => x"C0C0BFA499C0A492",
-24024 => x"C0C0BFA499C0A499",
-24023 => x"C0C0BFA499C0A4B0",
-24022 => x"C0C0BFA499C0A4A4",
-24021 => x"C0C0BFA499C0A4F9",
-24020 => x"C0C0BFA499C0A4C0",
-24019 => x"C0C0BFA499C0F990",
-24018 => x"C0C0BFA499C0F980",
-24017 => x"C0C0BFA499C0F9F8",
-24016 => x"C0C0BFA499C0F982",
-24015 => x"C0C0BFA499C0F992",
-24014 => x"C0C0BFA499C0F999",
-24013 => x"C0C0BFA499C0F9B0",
-24012 => x"C0C0BFA499C0F9A4",
-24011 => x"C0C0BFA499C0F9F9",
-24010 => x"C0C0BFA499C0F9C0",
-24009 => x"C0C0BFA499C0C090",
-24008 => x"C0C0BFA499C0C080",
-24007 => x"C0C0BFA499C0C0F8",
-24006 => x"C0C0BFA499C0C082",
-24005 => x"C0C0BFA499C0C092",
-24004 => x"C0C0BFA499C0C099",
-24003 => x"C0C0BFA499C0C0B0",
-24002 => x"C0C0BFA499C0C0A4",
-24001 => x"C0C0BFA499C0C0F9",
-24000 => x"C0C0BFA499C0C0C0",
-23999 => x"C0C0BFA4B0909090",
-23998 => x"C0C0BFA4B0909080",
-23997 => x"C0C0BFA4B09090F8",
-23996 => x"C0C0BFA4B0909082",
-23995 => x"C0C0BFA4B0909092",
-23994 => x"C0C0BFA4B0909099",
-23993 => x"C0C0BFA4B09090B0",
-23992 => x"C0C0BFA4B09090A4",
-23991 => x"C0C0BFA4B09090F9",
-23990 => x"C0C0BFA4B09090C0",
-23989 => x"C0C0BFA4B0908090",
-23988 => x"C0C0BFA4B0908080",
-23987 => x"C0C0BFA4B09080F8",
-23986 => x"C0C0BFA4B0908082",
-23985 => x"C0C0BFA4B0908092",
-23984 => x"C0C0BFA4B0908099",
-23983 => x"C0C0BFA4B09080B0",
-23982 => x"C0C0BFA4B09080A4",
-23981 => x"C0C0BFA4B09080F9",
-23980 => x"C0C0BFA4B09080C0",
-23979 => x"C0C0BFA4B090F890",
-23978 => x"C0C0BFA4B090F880",
-23977 => x"C0C0BFA4B090F8F8",
-23976 => x"C0C0BFA4B090F882",
-23975 => x"C0C0BFA4B090F892",
-23974 => x"C0C0BFA4B090F899",
-23973 => x"C0C0BFA4B090F8B0",
-23972 => x"C0C0BFA4B090F8A4",
-23971 => x"C0C0BFA4B090F8F9",
-23970 => x"C0C0BFA4B090F8C0",
-23969 => x"C0C0BFA4B0908290",
-23968 => x"C0C0BFA4B0908280",
-23967 => x"C0C0BFA4B09082F8",
-23966 => x"C0C0BFA4B0908282",
-23965 => x"C0C0BFA4B0908292",
-23964 => x"C0C0BFA4B0908299",
-23963 => x"C0C0BFA4B09082B0",
-23962 => x"C0C0BFA4B09082A4",
-23961 => x"C0C0BFA4B09082F9",
-23960 => x"C0C0BFA4B09082C0",
-23959 => x"C0C0BFA4B0909290",
-23958 => x"C0C0BFA4B0909280",
-23957 => x"C0C0BFA4B09092F8",
-23956 => x"C0C0BFA4B0909282",
-23955 => x"C0C0BFA4B0909292",
-23954 => x"C0C0BFA4B0909299",
-23953 => x"C0C0BFA4B09092B0",
-23952 => x"C0C0BFA4B09092A4",
-23951 => x"C0C0BFA4B09092F9",
-23950 => x"C0C0BFA4B09092C0",
-23949 => x"C0C0BFA4B0909990",
-23948 => x"C0C0BFA4B0909980",
-23947 => x"C0C0BFA4B09099F8",
-23946 => x"C0C0BFA4B0909982",
-23945 => x"C0C0BFA4B0909992",
-23944 => x"C0C0BFA4B0909999",
-23943 => x"C0C0BFA4B09099B0",
-23942 => x"C0C0BFA4B09099A4",
-23941 => x"C0C0BFA4B09099F9",
-23940 => x"C0C0BFA4B09099C0",
-23939 => x"C0C0BFA4B090B090",
-23938 => x"C0C0BFA4B090B080",
-23937 => x"C0C0BFA4B090B0F8",
-23936 => x"C0C0BFA4B090B082",
-23935 => x"C0C0BFA4B090B092",
-23934 => x"C0C0BFA4B090B099",
-23933 => x"C0C0BFA4B090B0B0",
-23932 => x"C0C0BFA4B090B0A4",
-23931 => x"C0C0BFA4B090B0F9",
-23930 => x"C0C0BFA4B090B0C0",
-23929 => x"C0C0BFA4B090A490",
-23928 => x"C0C0BFA4B090A480",
-23927 => x"C0C0BFA4B090A4F8",
-23926 => x"C0C0BFA4B090A482",
-23925 => x"C0C0BFA4B090A492",
-23924 => x"C0C0BFA4B090A499",
-23923 => x"C0C0BFA4B090A4B0",
-23922 => x"C0C0BFA4B090A4A4",
-23921 => x"C0C0BFA4B090A4F9",
-23920 => x"C0C0BFA4B090A4C0",
-23919 => x"C0C0BFA4B090F990",
-23918 => x"C0C0BFA4B090F980",
-23917 => x"C0C0BFA4B090F9F8",
-23916 => x"C0C0BFA4B090F982",
-23915 => x"C0C0BFA4B090F992",
-23914 => x"C0C0BFA4B090F999",
-23913 => x"C0C0BFA4B090F9B0",
-23912 => x"C0C0BFA4B090F9A4",
-23911 => x"C0C0BFA4B090F9F9",
-23910 => x"C0C0BFA4B090F9C0",
-23909 => x"C0C0BFA4B090C090",
-23908 => x"C0C0BFA4B090C080",
-23907 => x"C0C0BFA4B090C0F8",
-23906 => x"C0C0BFA4B090C082",
-23905 => x"C0C0BFA4B090C092",
-23904 => x"C0C0BFA4B090C099",
-23903 => x"C0C0BFA4B090C0B0",
-23902 => x"C0C0BFA4B090C0A4",
-23901 => x"C0C0BFA4B090C0F9",
-23900 => x"C0C0BFA4B090C0C0",
-23899 => x"C0C0BFA4B0809090",
-23898 => x"C0C0BFA4B0809080",
-23897 => x"C0C0BFA4B08090F8",
-23896 => x"C0C0BFA4B0809082",
-23895 => x"C0C0BFA4B0809092",
-23894 => x"C0C0BFA4B0809099",
-23893 => x"C0C0BFA4B08090B0",
-23892 => x"C0C0BFA4B08090A4",
-23891 => x"C0C0BFA4B08090F9",
-23890 => x"C0C0BFA4B08090C0",
-23889 => x"C0C0BFA4B0808090",
-23888 => x"C0C0BFA4B0808080",
-23887 => x"C0C0BFA4B08080F8",
-23886 => x"C0C0BFA4B0808082",
-23885 => x"C0C0BFA4B0808092",
-23884 => x"C0C0BFA4B0808099",
-23883 => x"C0C0BFA4B08080B0",
-23882 => x"C0C0BFA4B08080A4",
-23881 => x"C0C0BFA4B08080F9",
-23880 => x"C0C0BFA4B08080C0",
-23879 => x"C0C0BFA4B080F890",
-23878 => x"C0C0BFA4B080F880",
-23877 => x"C0C0BFA4B080F8F8",
-23876 => x"C0C0BFA4B080F882",
-23875 => x"C0C0BFA4B080F892",
-23874 => x"C0C0BFA4B080F899",
-23873 => x"C0C0BFA4B080F8B0",
-23872 => x"C0C0BFA4B080F8A4",
-23871 => x"C0C0BFA4B080F8F9",
-23870 => x"C0C0BFA4B080F8C0",
-23869 => x"C0C0BFA4B0808290",
-23868 => x"C0C0BFA4B0808280",
-23867 => x"C0C0BFA4B08082F8",
-23866 => x"C0C0BFA4B0808282",
-23865 => x"C0C0BFA4B0808292",
-23864 => x"C0C0BFA4B0808299",
-23863 => x"C0C0BFA4B08082B0",
-23862 => x"C0C0BFA4B08082A4",
-23861 => x"C0C0BFA4B08082F9",
-23860 => x"C0C0BFA4B08082C0",
-23859 => x"C0C0BFA4B0809290",
-23858 => x"C0C0BFA4B0809280",
-23857 => x"C0C0BFA4B08092F8",
-23856 => x"C0C0BFA4B0809282",
-23855 => x"C0C0BFA4B0809292",
-23854 => x"C0C0BFA4B0809299",
-23853 => x"C0C0BFA4B08092B0",
-23852 => x"C0C0BFA4B08092A4",
-23851 => x"C0C0BFA4B08092F9",
-23850 => x"C0C0BFA4B08092C0",
-23849 => x"C0C0BFA4B0809990",
-23848 => x"C0C0BFA4B0809980",
-23847 => x"C0C0BFA4B08099F8",
-23846 => x"C0C0BFA4B0809982",
-23845 => x"C0C0BFA4B0809992",
-23844 => x"C0C0BFA4B0809999",
-23843 => x"C0C0BFA4B08099B0",
-23842 => x"C0C0BFA4B08099A4",
-23841 => x"C0C0BFA4B08099F9",
-23840 => x"C0C0BFA4B08099C0",
-23839 => x"C0C0BFA4B080B090",
-23838 => x"C0C0BFA4B080B080",
-23837 => x"C0C0BFA4B080B0F8",
-23836 => x"C0C0BFA4B080B082",
-23835 => x"C0C0BFA4B080B092",
-23834 => x"C0C0BFA4B080B099",
-23833 => x"C0C0BFA4B080B0B0",
-23832 => x"C0C0BFA4B080B0A4",
-23831 => x"C0C0BFA4B080B0F9",
-23830 => x"C0C0BFA4B080B0C0",
-23829 => x"C0C0BFA4B080A490",
-23828 => x"C0C0BFA4B080A480",
-23827 => x"C0C0BFA4B080A4F8",
-23826 => x"C0C0BFA4B080A482",
-23825 => x"C0C0BFA4B080A492",
-23824 => x"C0C0BFA4B080A499",
-23823 => x"C0C0BFA4B080A4B0",
-23822 => x"C0C0BFA4B080A4A4",
-23821 => x"C0C0BFA4B080A4F9",
-23820 => x"C0C0BFA4B080A4C0",
-23819 => x"C0C0BFA4B080F990",
-23818 => x"C0C0BFA4B080F980",
-23817 => x"C0C0BFA4B080F9F8",
-23816 => x"C0C0BFA4B080F982",
-23815 => x"C0C0BFA4B080F992",
-23814 => x"C0C0BFA4B080F999",
-23813 => x"C0C0BFA4B080F9B0",
-23812 => x"C0C0BFA4B080F9A4",
-23811 => x"C0C0BFA4B080F9F9",
-23810 => x"C0C0BFA4B080F9C0",
-23809 => x"C0C0BFA4B080C090",
-23808 => x"C0C0BFA4B080C080",
-23807 => x"C0C0BFA4B080C0F8",
-23806 => x"C0C0BFA4B080C082",
-23805 => x"C0C0BFA4B080C092",
-23804 => x"C0C0BFA4B080C099",
-23803 => x"C0C0BFA4B080C0B0",
-23802 => x"C0C0BFA4B080C0A4",
-23801 => x"C0C0BFA4B080C0F9",
-23800 => x"C0C0BFA4B080C0C0",
-23799 => x"C0C0BFA4B0F89090",
-23798 => x"C0C0BFA4B0F89080",
-23797 => x"C0C0BFA4B0F890F8",
-23796 => x"C0C0BFA4B0F89082",
-23795 => x"C0C0BFA4B0F89092",
-23794 => x"C0C0BFA4B0F89099",
-23793 => x"C0C0BFA4B0F890B0",
-23792 => x"C0C0BFA4B0F890A4",
-23791 => x"C0C0BFA4B0F890F9",
-23790 => x"C0C0BFA4B0F890C0",
-23789 => x"C0C0BFA4B0F88090",
-23788 => x"C0C0BFA4B0F88080",
-23787 => x"C0C0BFA4B0F880F8",
-23786 => x"C0C0BFA4B0F88082",
-23785 => x"C0C0BFA4B0F88092",
-23784 => x"C0C0BFA4B0F88099",
-23783 => x"C0C0BFA4B0F880B0",
-23782 => x"C0C0BFA4B0F880A4",
-23781 => x"C0C0BFA4B0F880F9",
-23780 => x"C0C0BFA4B0F880C0",
-23779 => x"C0C0BFA4B0F8F890",
-23778 => x"C0C0BFA4B0F8F880",
-23777 => x"C0C0BFA4B0F8F8F8",
-23776 => x"C0C0BFA4B0F8F882",
-23775 => x"C0C0BFA4B0F8F892",
-23774 => x"C0C0BFA4B0F8F899",
-23773 => x"C0C0BFA4B0F8F8B0",
-23772 => x"C0C0BFA4B0F8F8A4",
-23771 => x"C0C0BFA4B0F8F8F9",
-23770 => x"C0C0BFA4B0F8F8C0",
-23769 => x"C0C0BFA4B0F88290",
-23768 => x"C0C0BFA4B0F88280",
-23767 => x"C0C0BFA4B0F882F8",
-23766 => x"C0C0BFA4B0F88282",
-23765 => x"C0C0BFA4B0F88292",
-23764 => x"C0C0BFA4B0F88299",
-23763 => x"C0C0BFA4B0F882B0",
-23762 => x"C0C0BFA4B0F882A4",
-23761 => x"C0C0BFA4B0F882F9",
-23760 => x"C0C0BFA4B0F882C0",
-23759 => x"C0C0BFA4B0F89290",
-23758 => x"C0C0BFA4B0F89280",
-23757 => x"C0C0BFA4B0F892F8",
-23756 => x"C0C0BFA4B0F89282",
-23755 => x"C0C0BFA4B0F89292",
-23754 => x"C0C0BFA4B0F89299",
-23753 => x"C0C0BFA4B0F892B0",
-23752 => x"C0C0BFA4B0F892A4",
-23751 => x"C0C0BFA4B0F892F9",
-23750 => x"C0C0BFA4B0F892C0",
-23749 => x"C0C0BFA4B0F89990",
-23748 => x"C0C0BFA4B0F89980",
-23747 => x"C0C0BFA4B0F899F8",
-23746 => x"C0C0BFA4B0F89982",
-23745 => x"C0C0BFA4B0F89992",
-23744 => x"C0C0BFA4B0F89999",
-23743 => x"C0C0BFA4B0F899B0",
-23742 => x"C0C0BFA4B0F899A4",
-23741 => x"C0C0BFA4B0F899F9",
-23740 => x"C0C0BFA4B0F899C0",
-23739 => x"C0C0BFA4B0F8B090",
-23738 => x"C0C0BFA4B0F8B080",
-23737 => x"C0C0BFA4B0F8B0F8",
-23736 => x"C0C0BFA4B0F8B082",
-23735 => x"C0C0BFA4B0F8B092",
-23734 => x"C0C0BFA4B0F8B099",
-23733 => x"C0C0BFA4B0F8B0B0",
-23732 => x"C0C0BFA4B0F8B0A4",
-23731 => x"C0C0BFA4B0F8B0F9",
-23730 => x"C0C0BFA4B0F8B0C0",
-23729 => x"C0C0BFA4B0F8A490",
-23728 => x"C0C0BFA4B0F8A480",
-23727 => x"C0C0BFA4B0F8A4F8",
-23726 => x"C0C0BFA4B0F8A482",
-23725 => x"C0C0BFA4B0F8A492",
-23724 => x"C0C0BFA4B0F8A499",
-23723 => x"C0C0BFA4B0F8A4B0",
-23722 => x"C0C0BFA4B0F8A4A4",
-23721 => x"C0C0BFA4B0F8A4F9",
-23720 => x"C0C0BFA4B0F8A4C0",
-23719 => x"C0C0BFA4B0F8F990",
-23718 => x"C0C0BFA4B0F8F980",
-23717 => x"C0C0BFA4B0F8F9F8",
-23716 => x"C0C0BFA4B0F8F982",
-23715 => x"C0C0BFA4B0F8F992",
-23714 => x"C0C0BFA4B0F8F999",
-23713 => x"C0C0BFA4B0F8F9B0",
-23712 => x"C0C0BFA4B0F8F9A4",
-23711 => x"C0C0BFA4B0F8F9F9",
-23710 => x"C0C0BFA4B0F8F9C0",
-23709 => x"C0C0BFA4B0F8C090",
-23708 => x"C0C0BFA4B0F8C080",
-23707 => x"C0C0BFA4B0F8C0F8",
-23706 => x"C0C0BFA4B0F8C082",
-23705 => x"C0C0BFA4B0F8C092",
-23704 => x"C0C0BFA4B0F8C099",
-23703 => x"C0C0BFA4B0F8C0B0",
-23702 => x"C0C0BFA4B0F8C0A4",
-23701 => x"C0C0BFA4B0F8C0F9",
-23700 => x"C0C0BFA4B0F8C0C0",
-23699 => x"C0C0BFA4B0829090",
-23698 => x"C0C0BFA4B0829080",
-23697 => x"C0C0BFA4B08290F8",
-23696 => x"C0C0BFA4B0829082",
-23695 => x"C0C0BFA4B0829092",
-23694 => x"C0C0BFA4B0829099",
-23693 => x"C0C0BFA4B08290B0",
-23692 => x"C0C0BFA4B08290A4",
-23691 => x"C0C0BFA4B08290F9",
-23690 => x"C0C0BFA4B08290C0",
-23689 => x"C0C0BFA4B0828090",
-23688 => x"C0C0BFA4B0828080",
-23687 => x"C0C0BFA4B08280F8",
-23686 => x"C0C0BFA4B0828082",
-23685 => x"C0C0BFA4B0828092",
-23684 => x"C0C0BFA4B0828099",
-23683 => x"C0C0BFA4B08280B0",
-23682 => x"C0C0BFA4B08280A4",
-23681 => x"C0C0BFA4B08280F9",
-23680 => x"C0C0BFA4B08280C0",
-23679 => x"C0C0BFA4B082F890",
-23678 => x"C0C0BFA4B082F880",
-23677 => x"C0C0BFA4B082F8F8",
-23676 => x"C0C0BFA4B082F882",
-23675 => x"C0C0BFA4B082F892",
-23674 => x"C0C0BFA4B082F899",
-23673 => x"C0C0BFA4B082F8B0",
-23672 => x"C0C0BFA4B082F8A4",
-23671 => x"C0C0BFA4B082F8F9",
-23670 => x"C0C0BFA4B082F8C0",
-23669 => x"C0C0BFA4B0828290",
-23668 => x"C0C0BFA4B0828280",
-23667 => x"C0C0BFA4B08282F8",
-23666 => x"C0C0BFA4B0828282",
-23665 => x"C0C0BFA4B0828292",
-23664 => x"C0C0BFA4B0828299",
-23663 => x"C0C0BFA4B08282B0",
-23662 => x"C0C0BFA4B08282A4",
-23661 => x"C0C0BFA4B08282F9",
-23660 => x"C0C0BFA4B08282C0",
-23659 => x"C0C0BFA4B0829290",
-23658 => x"C0C0BFA4B0829280",
-23657 => x"C0C0BFA4B08292F8",
-23656 => x"C0C0BFA4B0829282",
-23655 => x"C0C0BFA4B0829292",
-23654 => x"C0C0BFA4B0829299",
-23653 => x"C0C0BFA4B08292B0",
-23652 => x"C0C0BFA4B08292A4",
-23651 => x"C0C0BFA4B08292F9",
-23650 => x"C0C0BFA4B08292C0",
-23649 => x"C0C0BFA4B0829990",
-23648 => x"C0C0BFA4B0829980",
-23647 => x"C0C0BFA4B08299F8",
-23646 => x"C0C0BFA4B0829982",
-23645 => x"C0C0BFA4B0829992",
-23644 => x"C0C0BFA4B0829999",
-23643 => x"C0C0BFA4B08299B0",
-23642 => x"C0C0BFA4B08299A4",
-23641 => x"C0C0BFA4B08299F9",
-23640 => x"C0C0BFA4B08299C0",
-23639 => x"C0C0BFA4B082B090",
-23638 => x"C0C0BFA4B082B080",
-23637 => x"C0C0BFA4B082B0F8",
-23636 => x"C0C0BFA4B082B082",
-23635 => x"C0C0BFA4B082B092",
-23634 => x"C0C0BFA4B082B099",
-23633 => x"C0C0BFA4B082B0B0",
-23632 => x"C0C0BFA4B082B0A4",
-23631 => x"C0C0BFA4B082B0F9",
-23630 => x"C0C0BFA4B082B0C0",
-23629 => x"C0C0BFA4B082A490",
-23628 => x"C0C0BFA4B082A480",
-23627 => x"C0C0BFA4B082A4F8",
-23626 => x"C0C0BFA4B082A482",
-23625 => x"C0C0BFA4B082A492",
-23624 => x"C0C0BFA4B082A499",
-23623 => x"C0C0BFA4B082A4B0",
-23622 => x"C0C0BFA4B082A4A4",
-23621 => x"C0C0BFA4B082A4F9",
-23620 => x"C0C0BFA4B082A4C0",
-23619 => x"C0C0BFA4B082F990",
-23618 => x"C0C0BFA4B082F980",
-23617 => x"C0C0BFA4B082F9F8",
-23616 => x"C0C0BFA4B082F982",
-23615 => x"C0C0BFA4B082F992",
-23614 => x"C0C0BFA4B082F999",
-23613 => x"C0C0BFA4B082F9B0",
-23612 => x"C0C0BFA4B082F9A4",
-23611 => x"C0C0BFA4B082F9F9",
-23610 => x"C0C0BFA4B082F9C0",
-23609 => x"C0C0BFA4B082C090",
-23608 => x"C0C0BFA4B082C080",
-23607 => x"C0C0BFA4B082C0F8",
-23606 => x"C0C0BFA4B082C082",
-23605 => x"C0C0BFA4B082C092",
-23604 => x"C0C0BFA4B082C099",
-23603 => x"C0C0BFA4B082C0B0",
-23602 => x"C0C0BFA4B082C0A4",
-23601 => x"C0C0BFA4B082C0F9",
-23600 => x"C0C0BFA4B082C0C0",
-23599 => x"C0C0BFA4B0929090",
-23598 => x"C0C0BFA4B0929080",
-23597 => x"C0C0BFA4B09290F8",
-23596 => x"C0C0BFA4B0929082",
-23595 => x"C0C0BFA4B0929092",
-23594 => x"C0C0BFA4B0929099",
-23593 => x"C0C0BFA4B09290B0",
-23592 => x"C0C0BFA4B09290A4",
-23591 => x"C0C0BFA4B09290F9",
-23590 => x"C0C0BFA4B09290C0",
-23589 => x"C0C0BFA4B0928090",
-23588 => x"C0C0BFA4B0928080",
-23587 => x"C0C0BFA4B09280F8",
-23586 => x"C0C0BFA4B0928082",
-23585 => x"C0C0BFA4B0928092",
-23584 => x"C0C0BFA4B0928099",
-23583 => x"C0C0BFA4B09280B0",
-23582 => x"C0C0BFA4B09280A4",
-23581 => x"C0C0BFA4B09280F9",
-23580 => x"C0C0BFA4B09280C0",
-23579 => x"C0C0BFA4B092F890",
-23578 => x"C0C0BFA4B092F880",
-23577 => x"C0C0BFA4B092F8F8",
-23576 => x"C0C0BFA4B092F882",
-23575 => x"C0C0BFA4B092F892",
-23574 => x"C0C0BFA4B092F899",
-23573 => x"C0C0BFA4B092F8B0",
-23572 => x"C0C0BFA4B092F8A4",
-23571 => x"C0C0BFA4B092F8F9",
-23570 => x"C0C0BFA4B092F8C0",
-23569 => x"C0C0BFA4B0928290",
-23568 => x"C0C0BFA4B0928280",
-23567 => x"C0C0BFA4B09282F8",
-23566 => x"C0C0BFA4B0928282",
-23565 => x"C0C0BFA4B0928292",
-23564 => x"C0C0BFA4B0928299",
-23563 => x"C0C0BFA4B09282B0",
-23562 => x"C0C0BFA4B09282A4",
-23561 => x"C0C0BFA4B09282F9",
-23560 => x"C0C0BFA4B09282C0",
-23559 => x"C0C0BFA4B0929290",
-23558 => x"C0C0BFA4B0929280",
-23557 => x"C0C0BFA4B09292F8",
-23556 => x"C0C0BFA4B0929282",
-23555 => x"C0C0BFA4B0929292",
-23554 => x"C0C0BFA4B0929299",
-23553 => x"C0C0BFA4B09292B0",
-23552 => x"C0C0BFA4B09292A4",
-23551 => x"C0C0BFA4B09292F9",
-23550 => x"C0C0BFA4B09292C0",
-23549 => x"C0C0BFA4B0929990",
-23548 => x"C0C0BFA4B0929980",
-23547 => x"C0C0BFA4B09299F8",
-23546 => x"C0C0BFA4B0929982",
-23545 => x"C0C0BFA4B0929992",
-23544 => x"C0C0BFA4B0929999",
-23543 => x"C0C0BFA4B09299B0",
-23542 => x"C0C0BFA4B09299A4",
-23541 => x"C0C0BFA4B09299F9",
-23540 => x"C0C0BFA4B09299C0",
-23539 => x"C0C0BFA4B092B090",
-23538 => x"C0C0BFA4B092B080",
-23537 => x"C0C0BFA4B092B0F8",
-23536 => x"C0C0BFA4B092B082",
-23535 => x"C0C0BFA4B092B092",
-23534 => x"C0C0BFA4B092B099",
-23533 => x"C0C0BFA4B092B0B0",
-23532 => x"C0C0BFA4B092B0A4",
-23531 => x"C0C0BFA4B092B0F9",
-23530 => x"C0C0BFA4B092B0C0",
-23529 => x"C0C0BFA4B092A490",
-23528 => x"C0C0BFA4B092A480",
-23527 => x"C0C0BFA4B092A4F8",
-23526 => x"C0C0BFA4B092A482",
-23525 => x"C0C0BFA4B092A492",
-23524 => x"C0C0BFA4B092A499",
-23523 => x"C0C0BFA4B092A4B0",
-23522 => x"C0C0BFA4B092A4A4",
-23521 => x"C0C0BFA4B092A4F9",
-23520 => x"C0C0BFA4B092A4C0",
-23519 => x"C0C0BFA4B092F990",
-23518 => x"C0C0BFA4B092F980",
-23517 => x"C0C0BFA4B092F9F8",
-23516 => x"C0C0BFA4B092F982",
-23515 => x"C0C0BFA4B092F992",
-23514 => x"C0C0BFA4B092F999",
-23513 => x"C0C0BFA4B092F9B0",
-23512 => x"C0C0BFA4B092F9A4",
-23511 => x"C0C0BFA4B092F9F9",
-23510 => x"C0C0BFA4B092F9C0",
-23509 => x"C0C0BFA4B092C090",
-23508 => x"C0C0BFA4B092C080",
-23507 => x"C0C0BFA4B092C0F8",
-23506 => x"C0C0BFA4B092C082",
-23505 => x"C0C0BFA4B092C092",
-23504 => x"C0C0BFA4B092C099",
-23503 => x"C0C0BFA4B092C0B0",
-23502 => x"C0C0BFA4B092C0A4",
-23501 => x"C0C0BFA4B092C0F9",
-23500 => x"C0C0BFA4B092C0C0",
-23499 => x"C0C0BFA4B0999090",
-23498 => x"C0C0BFA4B0999080",
-23497 => x"C0C0BFA4B09990F8",
-23496 => x"C0C0BFA4B0999082",
-23495 => x"C0C0BFA4B0999092",
-23494 => x"C0C0BFA4B0999099",
-23493 => x"C0C0BFA4B09990B0",
-23492 => x"C0C0BFA4B09990A4",
-23491 => x"C0C0BFA4B09990F9",
-23490 => x"C0C0BFA4B09990C0",
-23489 => x"C0C0BFA4B0998090",
-23488 => x"C0C0BFA4B0998080",
-23487 => x"C0C0BFA4B09980F8",
-23486 => x"C0C0BFA4B0998082",
-23485 => x"C0C0BFA4B0998092",
-23484 => x"C0C0BFA4B0998099",
-23483 => x"C0C0BFA4B09980B0",
-23482 => x"C0C0BFA4B09980A4",
-23481 => x"C0C0BFA4B09980F9",
-23480 => x"C0C0BFA4B09980C0",
-23479 => x"C0C0BFA4B099F890",
-23478 => x"C0C0BFA4B099F880",
-23477 => x"C0C0BFA4B099F8F8",
-23476 => x"C0C0BFA4B099F882",
-23475 => x"C0C0BFA4B099F892",
-23474 => x"C0C0BFA4B099F899",
-23473 => x"C0C0BFA4B099F8B0",
-23472 => x"C0C0BFA4B099F8A4",
-23471 => x"C0C0BFA4B099F8F9",
-23470 => x"C0C0BFA4B099F8C0",
-23469 => x"C0C0BFA4B0998290",
-23468 => x"C0C0BFA4B0998280",
-23467 => x"C0C0BFA4B09982F8",
-23466 => x"C0C0BFA4B0998282",
-23465 => x"C0C0BFA4B0998292",
-23464 => x"C0C0BFA4B0998299",
-23463 => x"C0C0BFA4B09982B0",
-23462 => x"C0C0BFA4B09982A4",
-23461 => x"C0C0BFA4B09982F9",
-23460 => x"C0C0BFA4B09982C0",
-23459 => x"C0C0BFA4B0999290",
-23458 => x"C0C0BFA4B0999280",
-23457 => x"C0C0BFA4B09992F8",
-23456 => x"C0C0BFA4B0999282",
-23455 => x"C0C0BFA4B0999292",
-23454 => x"C0C0BFA4B0999299",
-23453 => x"C0C0BFA4B09992B0",
-23452 => x"C0C0BFA4B09992A4",
-23451 => x"C0C0BFA4B09992F9",
-23450 => x"C0C0BFA4B09992C0",
-23449 => x"C0C0BFA4B0999990",
-23448 => x"C0C0BFA4B0999980",
-23447 => x"C0C0BFA4B09999F8",
-23446 => x"C0C0BFA4B0999982",
-23445 => x"C0C0BFA4B0999992",
-23444 => x"C0C0BFA4B0999999",
-23443 => x"C0C0BFA4B09999B0",
-23442 => x"C0C0BFA4B09999A4",
-23441 => x"C0C0BFA4B09999F9",
-23440 => x"C0C0BFA4B09999C0",
-23439 => x"C0C0BFA4B099B090",
-23438 => x"C0C0BFA4B099B080",
-23437 => x"C0C0BFA4B099B0F8",
-23436 => x"C0C0BFA4B099B082",
-23435 => x"C0C0BFA4B099B092",
-23434 => x"C0C0BFA4B099B099",
-23433 => x"C0C0BFA4B099B0B0",
-23432 => x"C0C0BFA4B099B0A4",
-23431 => x"C0C0BFA4B099B0F9",
-23430 => x"C0C0BFA4B099B0C0",
-23429 => x"C0C0BFA4B099A490",
-23428 => x"C0C0BFA4B099A480",
-23427 => x"C0C0BFA4B099A4F8",
-23426 => x"C0C0BFA4B099A482",
-23425 => x"C0C0BFA4B099A492",
-23424 => x"C0C0BFA4B099A499",
-23423 => x"C0C0BFA4B099A4B0",
-23422 => x"C0C0BFA4B099A4A4",
-23421 => x"C0C0BFA4B099A4F9",
-23420 => x"C0C0BFA4B099A4C0",
-23419 => x"C0C0BFA4B099F990",
-23418 => x"C0C0BFA4B099F980",
-23417 => x"C0C0BFA4B099F9F8",
-23416 => x"C0C0BFA4B099F982",
-23415 => x"C0C0BFA4B099F992",
-23414 => x"C0C0BFA4B099F999",
-23413 => x"C0C0BFA4B099F9B0",
-23412 => x"C0C0BFA4B099F9A4",
-23411 => x"C0C0BFA4B099F9F9",
-23410 => x"C0C0BFA4B099F9C0",
-23409 => x"C0C0BFA4B099C090",
-23408 => x"C0C0BFA4B099C080",
-23407 => x"C0C0BFA4B099C0F8",
-23406 => x"C0C0BFA4B099C082",
-23405 => x"C0C0BFA4B099C092",
-23404 => x"C0C0BFA4B099C099",
-23403 => x"C0C0BFA4B099C0B0",
-23402 => x"C0C0BFA4B099C0A4",
-23401 => x"C0C0BFA4B099C0F9",
-23400 => x"C0C0BFA4B099C0C0",
-23399 => x"C0C0BFA4B0B09090",
-23398 => x"C0C0BFA4B0B09080",
-23397 => x"C0C0BFA4B0B090F8",
-23396 => x"C0C0BFA4B0B09082",
-23395 => x"C0C0BFA4B0B09092",
-23394 => x"C0C0BFA4B0B09099",
-23393 => x"C0C0BFA4B0B090B0",
-23392 => x"C0C0BFA4B0B090A4",
-23391 => x"C0C0BFA4B0B090F9",
-23390 => x"C0C0BFA4B0B090C0",
-23389 => x"C0C0BFA4B0B08090",
-23388 => x"C0C0BFA4B0B08080",
-23387 => x"C0C0BFA4B0B080F8",
-23386 => x"C0C0BFA4B0B08082",
-23385 => x"C0C0BFA4B0B08092",
-23384 => x"C0C0BFA4B0B08099",
-23383 => x"C0C0BFA4B0B080B0",
-23382 => x"C0C0BFA4B0B080A4",
-23381 => x"C0C0BFA4B0B080F9",
-23380 => x"C0C0BFA4B0B080C0",
-23379 => x"C0C0BFA4B0B0F890",
-23378 => x"C0C0BFA4B0B0F880",
-23377 => x"C0C0BFA4B0B0F8F8",
-23376 => x"C0C0BFA4B0B0F882",
-23375 => x"C0C0BFA4B0B0F892",
-23374 => x"C0C0BFA4B0B0F899",
-23373 => x"C0C0BFA4B0B0F8B0",
-23372 => x"C0C0BFA4B0B0F8A4",
-23371 => x"C0C0BFA4B0B0F8F9",
-23370 => x"C0C0BFA4B0B0F8C0",
-23369 => x"C0C0BFA4B0B08290",
-23368 => x"C0C0BFA4B0B08280",
-23367 => x"C0C0BFA4B0B082F8",
-23366 => x"C0C0BFA4B0B08282",
-23365 => x"C0C0BFA4B0B08292",
-23364 => x"C0C0BFA4B0B08299",
-23363 => x"C0C0BFA4B0B082B0",
-23362 => x"C0C0BFA4B0B082A4",
-23361 => x"C0C0BFA4B0B082F9",
-23360 => x"C0C0BFA4B0B082C0",
-23359 => x"C0C0BFA4B0B09290",
-23358 => x"C0C0BFA4B0B09280",
-23357 => x"C0C0BFA4B0B092F8",
-23356 => x"C0C0BFA4B0B09282",
-23355 => x"C0C0BFA4B0B09292",
-23354 => x"C0C0BFA4B0B09299",
-23353 => x"C0C0BFA4B0B092B0",
-23352 => x"C0C0BFA4B0B092A4",
-23351 => x"C0C0BFA4B0B092F9",
-23350 => x"C0C0BFA4B0B092C0",
-23349 => x"C0C0BFA4B0B09990",
-23348 => x"C0C0BFA4B0B09980",
-23347 => x"C0C0BFA4B0B099F8",
-23346 => x"C0C0BFA4B0B09982",
-23345 => x"C0C0BFA4B0B09992",
-23344 => x"C0C0BFA4B0B09999",
-23343 => x"C0C0BFA4B0B099B0",
-23342 => x"C0C0BFA4B0B099A4",
-23341 => x"C0C0BFA4B0B099F9",
-23340 => x"C0C0BFA4B0B099C0",
-23339 => x"C0C0BFA4B0B0B090",
-23338 => x"C0C0BFA4B0B0B080",
-23337 => x"C0C0BFA4B0B0B0F8",
-23336 => x"C0C0BFA4B0B0B082",
-23335 => x"C0C0BFA4B0B0B092",
-23334 => x"C0C0BFA4B0B0B099",
-23333 => x"C0C0BFA4B0B0B0B0",
-23332 => x"C0C0BFA4B0B0B0A4",
-23331 => x"C0C0BFA4B0B0B0F9",
-23330 => x"C0C0BFA4B0B0B0C0",
-23329 => x"C0C0BFA4B0B0A490",
-23328 => x"C0C0BFA4B0B0A480",
-23327 => x"C0C0BFA4B0B0A4F8",
-23326 => x"C0C0BFA4B0B0A482",
-23325 => x"C0C0BFA4B0B0A492",
-23324 => x"C0C0BFA4B0B0A499",
-23323 => x"C0C0BFA4B0B0A4B0",
-23322 => x"C0C0BFA4B0B0A4A4",
-23321 => x"C0C0BFA4B0B0A4F9",
-23320 => x"C0C0BFA4B0B0A4C0",
-23319 => x"C0C0BFA4B0B0F990",
-23318 => x"C0C0BFA4B0B0F980",
-23317 => x"C0C0BFA4B0B0F9F8",
-23316 => x"C0C0BFA4B0B0F982",
-23315 => x"C0C0BFA4B0B0F992",
-23314 => x"C0C0BFA4B0B0F999",
-23313 => x"C0C0BFA4B0B0F9B0",
-23312 => x"C0C0BFA4B0B0F9A4",
-23311 => x"C0C0BFA4B0B0F9F9",
-23310 => x"C0C0BFA4B0B0F9C0",
-23309 => x"C0C0BFA4B0B0C090",
-23308 => x"C0C0BFA4B0B0C080",
-23307 => x"C0C0BFA4B0B0C0F8",
-23306 => x"C0C0BFA4B0B0C082",
-23305 => x"C0C0BFA4B0B0C092",
-23304 => x"C0C0BFA4B0B0C099",
-23303 => x"C0C0BFA4B0B0C0B0",
-23302 => x"C0C0BFA4B0B0C0A4",
-23301 => x"C0C0BFA4B0B0C0F9",
-23300 => x"C0C0BFA4B0B0C0C0",
-23299 => x"C0C0BFA4B0A49090",
-23298 => x"C0C0BFA4B0A49080",
-23297 => x"C0C0BFA4B0A490F8",
-23296 => x"C0C0BFA4B0A49082",
-23295 => x"C0C0BFA4B0A49092",
-23294 => x"C0C0BFA4B0A49099",
-23293 => x"C0C0BFA4B0A490B0",
-23292 => x"C0C0BFA4B0A490A4",
-23291 => x"C0C0BFA4B0A490F9",
-23290 => x"C0C0BFA4B0A490C0",
-23289 => x"C0C0BFA4B0A48090",
-23288 => x"C0C0BFA4B0A48080",
-23287 => x"C0C0BFA4B0A480F8",
-23286 => x"C0C0BFA4B0A48082",
-23285 => x"C0C0BFA4B0A48092",
-23284 => x"C0C0BFA4B0A48099",
-23283 => x"C0C0BFA4B0A480B0",
-23282 => x"C0C0BFA4B0A480A4",
-23281 => x"C0C0BFA4B0A480F9",
-23280 => x"C0C0BFA4B0A480C0",
-23279 => x"C0C0BFA4B0A4F890",
-23278 => x"C0C0BFA4B0A4F880",
-23277 => x"C0C0BFA4B0A4F8F8",
-23276 => x"C0C0BFA4B0A4F882",
-23275 => x"C0C0BFA4B0A4F892",
-23274 => x"C0C0BFA4B0A4F899",
-23273 => x"C0C0BFA4B0A4F8B0",
-23272 => x"C0C0BFA4B0A4F8A4",
-23271 => x"C0C0BFA4B0A4F8F9",
-23270 => x"C0C0BFA4B0A4F8C0",
-23269 => x"C0C0BFA4B0A48290",
-23268 => x"C0C0BFA4B0A48280",
-23267 => x"C0C0BFA4B0A482F8",
-23266 => x"C0C0BFA4B0A48282",
-23265 => x"C0C0BFA4B0A48292",
-23264 => x"C0C0BFA4B0A48299",
-23263 => x"C0C0BFA4B0A482B0",
-23262 => x"C0C0BFA4B0A482A4",
-23261 => x"C0C0BFA4B0A482F9",
-23260 => x"C0C0BFA4B0A482C0",
-23259 => x"C0C0BFA4B0A49290",
-23258 => x"C0C0BFA4B0A49280",
-23257 => x"C0C0BFA4B0A492F8",
-23256 => x"C0C0BFA4B0A49282",
-23255 => x"C0C0BFA4B0A49292",
-23254 => x"C0C0BFA4B0A49299",
-23253 => x"C0C0BFA4B0A492B0",
-23252 => x"C0C0BFA4B0A492A4",
-23251 => x"C0C0BFA4B0A492F9",
-23250 => x"C0C0BFA4B0A492C0",
-23249 => x"C0C0BFA4B0A49990",
-23248 => x"C0C0BFA4B0A49980",
-23247 => x"C0C0BFA4B0A499F8",
-23246 => x"C0C0BFA4B0A49982",
-23245 => x"C0C0BFA4B0A49992",
-23244 => x"C0C0BFA4B0A49999",
-23243 => x"C0C0BFA4B0A499B0",
-23242 => x"C0C0BFA4B0A499A4",
-23241 => x"C0C0BFA4B0A499F9",
-23240 => x"C0C0BFA4B0A499C0",
-23239 => x"C0C0BFA4B0A4B090",
-23238 => x"C0C0BFA4B0A4B080",
-23237 => x"C0C0BFA4B0A4B0F8",
-23236 => x"C0C0BFA4B0A4B082",
-23235 => x"C0C0BFA4B0A4B092",
-23234 => x"C0C0BFA4B0A4B099",
-23233 => x"C0C0BFA4B0A4B0B0",
-23232 => x"C0C0BFA4B0A4B0A4",
-23231 => x"C0C0BFA4B0A4B0F9",
-23230 => x"C0C0BFA4B0A4B0C0",
-23229 => x"C0C0BFA4B0A4A490",
-23228 => x"C0C0BFA4B0A4A480",
-23227 => x"C0C0BFA4B0A4A4F8",
-23226 => x"C0C0BFA4B0A4A482",
-23225 => x"C0C0BFA4B0A4A492",
-23224 => x"C0C0BFA4B0A4A499",
-23223 => x"C0C0BFA4B0A4A4B0",
-23222 => x"C0C0BFA4B0A4A4A4",
-23221 => x"C0C0BFA4B0A4A4F9",
-23220 => x"C0C0BFA4B0A4A4C0",
-23219 => x"C0C0BFA4B0A4F990",
-23218 => x"C0C0BFA4B0A4F980",
-23217 => x"C0C0BFA4B0A4F9F8",
-23216 => x"C0C0BFA4B0A4F982",
-23215 => x"C0C0BFA4B0A4F992",
-23214 => x"C0C0BFA4B0A4F999",
-23213 => x"C0C0BFA4B0A4F9B0",
-23212 => x"C0C0BFA4B0A4F9A4",
-23211 => x"C0C0BFA4B0A4F9F9",
-23210 => x"C0C0BFA4B0A4F9C0",
-23209 => x"C0C0BFA4B0A4C090",
-23208 => x"C0C0BFA4B0A4C080",
-23207 => x"C0C0BFA4B0A4C0F8",
-23206 => x"C0C0BFA4B0A4C082",
-23205 => x"C0C0BFA4B0A4C092",
-23204 => x"C0C0BFA4B0A4C099",
-23203 => x"C0C0BFA4B0A4C0B0",
-23202 => x"C0C0BFA4B0A4C0A4",
-23201 => x"C0C0BFA4B0A4C0F9",
-23200 => x"C0C0BFA4B0A4C0C0",
-23199 => x"C0C0BFA4B0F99090",
-23198 => x"C0C0BFA4B0F99080",
-23197 => x"C0C0BFA4B0F990F8",
-23196 => x"C0C0BFA4B0F99082",
-23195 => x"C0C0BFA4B0F99092",
-23194 => x"C0C0BFA4B0F99099",
-23193 => x"C0C0BFA4B0F990B0",
-23192 => x"C0C0BFA4B0F990A4",
-23191 => x"C0C0BFA4B0F990F9",
-23190 => x"C0C0BFA4B0F990C0",
-23189 => x"C0C0BFA4B0F98090",
-23188 => x"C0C0BFA4B0F98080",
-23187 => x"C0C0BFA4B0F980F8",
-23186 => x"C0C0BFA4B0F98082",
-23185 => x"C0C0BFA4B0F98092",
-23184 => x"C0C0BFA4B0F98099",
-23183 => x"C0C0BFA4B0F980B0",
-23182 => x"C0C0BFA4B0F980A4",
-23181 => x"C0C0BFA4B0F980F9",
-23180 => x"C0C0BFA4B0F980C0",
-23179 => x"C0C0BFA4B0F9F890",
-23178 => x"C0C0BFA4B0F9F880",
-23177 => x"C0C0BFA4B0F9F8F8",
-23176 => x"C0C0BFA4B0F9F882",
-23175 => x"C0C0BFA4B0F9F892",
-23174 => x"C0C0BFA4B0F9F899",
-23173 => x"C0C0BFA4B0F9F8B0",
-23172 => x"C0C0BFA4B0F9F8A4",
-23171 => x"C0C0BFA4B0F9F8F9",
-23170 => x"C0C0BFA4B0F9F8C0",
-23169 => x"C0C0BFA4B0F98290",
-23168 => x"C0C0BFA4B0F98280",
-23167 => x"C0C0BFA4B0F982F8",
-23166 => x"C0C0BFA4B0F98282",
-23165 => x"C0C0BFA4B0F98292",
-23164 => x"C0C0BFA4B0F98299",
-23163 => x"C0C0BFA4B0F982B0",
-23162 => x"C0C0BFA4B0F982A4",
-23161 => x"C0C0BFA4B0F982F9",
-23160 => x"C0C0BFA4B0F982C0",
-23159 => x"C0C0BFA4B0F99290",
-23158 => x"C0C0BFA4B0F99280",
-23157 => x"C0C0BFA4B0F992F8",
-23156 => x"C0C0BFA4B0F99282",
-23155 => x"C0C0BFA4B0F99292",
-23154 => x"C0C0BFA4B0F99299",
-23153 => x"C0C0BFA4B0F992B0",
-23152 => x"C0C0BFA4B0F992A4",
-23151 => x"C0C0BFA4B0F992F9",
-23150 => x"C0C0BFA4B0F992C0",
-23149 => x"C0C0BFA4B0F99990",
-23148 => x"C0C0BFA4B0F99980",
-23147 => x"C0C0BFA4B0F999F8",
-23146 => x"C0C0BFA4B0F99982",
-23145 => x"C0C0BFA4B0F99992",
-23144 => x"C0C0BFA4B0F99999",
-23143 => x"C0C0BFA4B0F999B0",
-23142 => x"C0C0BFA4B0F999A4",
-23141 => x"C0C0BFA4B0F999F9",
-23140 => x"C0C0BFA4B0F999C0",
-23139 => x"C0C0BFA4B0F9B090",
-23138 => x"C0C0BFA4B0F9B080",
-23137 => x"C0C0BFA4B0F9B0F8",
-23136 => x"C0C0BFA4B0F9B082",
-23135 => x"C0C0BFA4B0F9B092",
-23134 => x"C0C0BFA4B0F9B099",
-23133 => x"C0C0BFA4B0F9B0B0",
-23132 => x"C0C0BFA4B0F9B0A4",
-23131 => x"C0C0BFA4B0F9B0F9",
-23130 => x"C0C0BFA4B0F9B0C0",
-23129 => x"C0C0BFA4B0F9A490",
-23128 => x"C0C0BFA4B0F9A480",
-23127 => x"C0C0BFA4B0F9A4F8",
-23126 => x"C0C0BFA4B0F9A482",
-23125 => x"C0C0BFA4B0F9A492",
-23124 => x"C0C0BFA4B0F9A499",
-23123 => x"C0C0BFA4B0F9A4B0",
-23122 => x"C0C0BFA4B0F9A4A4",
-23121 => x"C0C0BFA4B0F9A4F9",
-23120 => x"C0C0BFA4B0F9A4C0",
-23119 => x"C0C0BFA4B0F9F990",
-23118 => x"C0C0BFA4B0F9F980",
-23117 => x"C0C0BFA4B0F9F9F8",
-23116 => x"C0C0BFA4B0F9F982",
-23115 => x"C0C0BFA4B0F9F992",
-23114 => x"C0C0BFA4B0F9F999",
-23113 => x"C0C0BFA4B0F9F9B0",
-23112 => x"C0C0BFA4B0F9F9A4",
-23111 => x"C0C0BFA4B0F9F9F9",
-23110 => x"C0C0BFA4B0F9F9C0",
-23109 => x"C0C0BFA4B0F9C090",
-23108 => x"C0C0BFA4B0F9C080",
-23107 => x"C0C0BFA4B0F9C0F8",
-23106 => x"C0C0BFA4B0F9C082",
-23105 => x"C0C0BFA4B0F9C092",
-23104 => x"C0C0BFA4B0F9C099",
-23103 => x"C0C0BFA4B0F9C0B0",
-23102 => x"C0C0BFA4B0F9C0A4",
-23101 => x"C0C0BFA4B0F9C0F9",
-23100 => x"C0C0BFA4B0F9C0C0",
-23099 => x"C0C0BFA4B0C09090",
-23098 => x"C0C0BFA4B0C09080",
-23097 => x"C0C0BFA4B0C090F8",
-23096 => x"C0C0BFA4B0C09082",
-23095 => x"C0C0BFA4B0C09092",
-23094 => x"C0C0BFA4B0C09099",
-23093 => x"C0C0BFA4B0C090B0",
-23092 => x"C0C0BFA4B0C090A4",
-23091 => x"C0C0BFA4B0C090F9",
-23090 => x"C0C0BFA4B0C090C0",
-23089 => x"C0C0BFA4B0C08090",
-23088 => x"C0C0BFA4B0C08080",
-23087 => x"C0C0BFA4B0C080F8",
-23086 => x"C0C0BFA4B0C08082",
-23085 => x"C0C0BFA4B0C08092",
-23084 => x"C0C0BFA4B0C08099",
-23083 => x"C0C0BFA4B0C080B0",
-23082 => x"C0C0BFA4B0C080A4",
-23081 => x"C0C0BFA4B0C080F9",
-23080 => x"C0C0BFA4B0C080C0",
-23079 => x"C0C0BFA4B0C0F890",
-23078 => x"C0C0BFA4B0C0F880",
-23077 => x"C0C0BFA4B0C0F8F8",
-23076 => x"C0C0BFA4B0C0F882",
-23075 => x"C0C0BFA4B0C0F892",
-23074 => x"C0C0BFA4B0C0F899",
-23073 => x"C0C0BFA4B0C0F8B0",
-23072 => x"C0C0BFA4B0C0F8A4",
-23071 => x"C0C0BFA4B0C0F8F9",
-23070 => x"C0C0BFA4B0C0F8C0",
-23069 => x"C0C0BFA4B0C08290",
-23068 => x"C0C0BFA4B0C08280",
-23067 => x"C0C0BFA4B0C082F8",
-23066 => x"C0C0BFA4B0C08282",
-23065 => x"C0C0BFA4B0C08292",
-23064 => x"C0C0BFA4B0C08299",
-23063 => x"C0C0BFA4B0C082B0",
-23062 => x"C0C0BFA4B0C082A4",
-23061 => x"C0C0BFA4B0C082F9",
-23060 => x"C0C0BFA4B0C082C0",
-23059 => x"C0C0BFA4B0C09290",
-23058 => x"C0C0BFA4B0C09280",
-23057 => x"C0C0BFA4B0C092F8",
-23056 => x"C0C0BFA4B0C09282",
-23055 => x"C0C0BFA4B0C09292",
-23054 => x"C0C0BFA4B0C09299",
-23053 => x"C0C0BFA4B0C092B0",
-23052 => x"C0C0BFA4B0C092A4",
-23051 => x"C0C0BFA4B0C092F9",
-23050 => x"C0C0BFA4B0C092C0",
-23049 => x"C0C0BFA4B0C09990",
-23048 => x"C0C0BFA4B0C09980",
-23047 => x"C0C0BFA4B0C099F8",
-23046 => x"C0C0BFA4B0C09982",
-23045 => x"C0C0BFA4B0C09992",
-23044 => x"C0C0BFA4B0C09999",
-23043 => x"C0C0BFA4B0C099B0",
-23042 => x"C0C0BFA4B0C099A4",
-23041 => x"C0C0BFA4B0C099F9",
-23040 => x"C0C0BFA4B0C099C0",
-23039 => x"C0C0BFA4B0C0B090",
-23038 => x"C0C0BFA4B0C0B080",
-23037 => x"C0C0BFA4B0C0B0F8",
-23036 => x"C0C0BFA4B0C0B082",
-23035 => x"C0C0BFA4B0C0B092",
-23034 => x"C0C0BFA4B0C0B099",
-23033 => x"C0C0BFA4B0C0B0B0",
-23032 => x"C0C0BFA4B0C0B0A4",
-23031 => x"C0C0BFA4B0C0B0F9",
-23030 => x"C0C0BFA4B0C0B0C0",
-23029 => x"C0C0BFA4B0C0A490",
-23028 => x"C0C0BFA4B0C0A480",
-23027 => x"C0C0BFA4B0C0A4F8",
-23026 => x"C0C0BFA4B0C0A482",
-23025 => x"C0C0BFA4B0C0A492",
-23024 => x"C0C0BFA4B0C0A499",
-23023 => x"C0C0BFA4B0C0A4B0",
-23022 => x"C0C0BFA4B0C0A4A4",
-23021 => x"C0C0BFA4B0C0A4F9",
-23020 => x"C0C0BFA4B0C0A4C0",
-23019 => x"C0C0BFA4B0C0F990",
-23018 => x"C0C0BFA4B0C0F980",
-23017 => x"C0C0BFA4B0C0F9F8",
-23016 => x"C0C0BFA4B0C0F982",
-23015 => x"C0C0BFA4B0C0F992",
-23014 => x"C0C0BFA4B0C0F999",
-23013 => x"C0C0BFA4B0C0F9B0",
-23012 => x"C0C0BFA4B0C0F9A4",
-23011 => x"C0C0BFA4B0C0F9F9",
-23010 => x"C0C0BFA4B0C0F9C0",
-23009 => x"C0C0BFA4B0C0C090",
-23008 => x"C0C0BFA4B0C0C080",
-23007 => x"C0C0BFA4B0C0C0F8",
-23006 => x"C0C0BFA4B0C0C082",
-23005 => x"C0C0BFA4B0C0C092",
-23004 => x"C0C0BFA4B0C0C099",
-23003 => x"C0C0BFA4B0C0C0B0",
-23002 => x"C0C0BFA4B0C0C0A4",
-23001 => x"C0C0BFA4B0C0C0F9",
-23000 => x"C0C0BFA4B0C0C0C0",
-22999 => x"C0C0BFA4A4909090",
-22998 => x"C0C0BFA4A4909080",
-22997 => x"C0C0BFA4A49090F8",
-22996 => x"C0C0BFA4A4909082",
-22995 => x"C0C0BFA4A4909092",
-22994 => x"C0C0BFA4A4909099",
-22993 => x"C0C0BFA4A49090B0",
-22992 => x"C0C0BFA4A49090A4",
-22991 => x"C0C0BFA4A49090F9",
-22990 => x"C0C0BFA4A49090C0",
-22989 => x"C0C0BFA4A4908090",
-22988 => x"C0C0BFA4A4908080",
-22987 => x"C0C0BFA4A49080F8",
-22986 => x"C0C0BFA4A4908082",
-22985 => x"C0C0BFA4A4908092",
-22984 => x"C0C0BFA4A4908099",
-22983 => x"C0C0BFA4A49080B0",
-22982 => x"C0C0BFA4A49080A4",
-22981 => x"C0C0BFA4A49080F9",
-22980 => x"C0C0BFA4A49080C0",
-22979 => x"C0C0BFA4A490F890",
-22978 => x"C0C0BFA4A490F880",
-22977 => x"C0C0BFA4A490F8F8",
-22976 => x"C0C0BFA4A490F882",
-22975 => x"C0C0BFA4A490F892",
-22974 => x"C0C0BFA4A490F899",
-22973 => x"C0C0BFA4A490F8B0",
-22972 => x"C0C0BFA4A490F8A4",
-22971 => x"C0C0BFA4A490F8F9",
-22970 => x"C0C0BFA4A490F8C0",
-22969 => x"C0C0BFA4A4908290",
-22968 => x"C0C0BFA4A4908280",
-22967 => x"C0C0BFA4A49082F8",
-22966 => x"C0C0BFA4A4908282",
-22965 => x"C0C0BFA4A4908292",
-22964 => x"C0C0BFA4A4908299",
-22963 => x"C0C0BFA4A49082B0",
-22962 => x"C0C0BFA4A49082A4",
-22961 => x"C0C0BFA4A49082F9",
-22960 => x"C0C0BFA4A49082C0",
-22959 => x"C0C0BFA4A4909290",
-22958 => x"C0C0BFA4A4909280",
-22957 => x"C0C0BFA4A49092F8",
-22956 => x"C0C0BFA4A4909282",
-22955 => x"C0C0BFA4A4909292",
-22954 => x"C0C0BFA4A4909299",
-22953 => x"C0C0BFA4A49092B0",
-22952 => x"C0C0BFA4A49092A4",
-22951 => x"C0C0BFA4A49092F9",
-22950 => x"C0C0BFA4A49092C0",
-22949 => x"C0C0BFA4A4909990",
-22948 => x"C0C0BFA4A4909980",
-22947 => x"C0C0BFA4A49099F8",
-22946 => x"C0C0BFA4A4909982",
-22945 => x"C0C0BFA4A4909992",
-22944 => x"C0C0BFA4A4909999",
-22943 => x"C0C0BFA4A49099B0",
-22942 => x"C0C0BFA4A49099A4",
-22941 => x"C0C0BFA4A49099F9",
-22940 => x"C0C0BFA4A49099C0",
-22939 => x"C0C0BFA4A490B090",
-22938 => x"C0C0BFA4A490B080",
-22937 => x"C0C0BFA4A490B0F8",
-22936 => x"C0C0BFA4A490B082",
-22935 => x"C0C0BFA4A490B092",
-22934 => x"C0C0BFA4A490B099",
-22933 => x"C0C0BFA4A490B0B0",
-22932 => x"C0C0BFA4A490B0A4",
-22931 => x"C0C0BFA4A490B0F9",
-22930 => x"C0C0BFA4A490B0C0",
-22929 => x"C0C0BFA4A490A490",
-22928 => x"C0C0BFA4A490A480",
-22927 => x"C0C0BFA4A490A4F8",
-22926 => x"C0C0BFA4A490A482",
-22925 => x"C0C0BFA4A490A492",
-22924 => x"C0C0BFA4A490A499",
-22923 => x"C0C0BFA4A490A4B0",
-22922 => x"C0C0BFA4A490A4A4",
-22921 => x"C0C0BFA4A490A4F9",
-22920 => x"C0C0BFA4A490A4C0",
-22919 => x"C0C0BFA4A490F990",
-22918 => x"C0C0BFA4A490F980",
-22917 => x"C0C0BFA4A490F9F8",
-22916 => x"C0C0BFA4A490F982",
-22915 => x"C0C0BFA4A490F992",
-22914 => x"C0C0BFA4A490F999",
-22913 => x"C0C0BFA4A490F9B0",
-22912 => x"C0C0BFA4A490F9A4",
-22911 => x"C0C0BFA4A490F9F9",
-22910 => x"C0C0BFA4A490F9C0",
-22909 => x"C0C0BFA4A490C090",
-22908 => x"C0C0BFA4A490C080",
-22907 => x"C0C0BFA4A490C0F8",
-22906 => x"C0C0BFA4A490C082",
-22905 => x"C0C0BFA4A490C092",
-22904 => x"C0C0BFA4A490C099",
-22903 => x"C0C0BFA4A490C0B0",
-22902 => x"C0C0BFA4A490C0A4",
-22901 => x"C0C0BFA4A490C0F9",
-22900 => x"C0C0BFA4A490C0C0",
-22899 => x"C0C0BFA4A4809090",
-22898 => x"C0C0BFA4A4809080",
-22897 => x"C0C0BFA4A48090F8",
-22896 => x"C0C0BFA4A4809082",
-22895 => x"C0C0BFA4A4809092",
-22894 => x"C0C0BFA4A4809099",
-22893 => x"C0C0BFA4A48090B0",
-22892 => x"C0C0BFA4A48090A4",
-22891 => x"C0C0BFA4A48090F9",
-22890 => x"C0C0BFA4A48090C0",
-22889 => x"C0C0BFA4A4808090",
-22888 => x"C0C0BFA4A4808080",
-22887 => x"C0C0BFA4A48080F8",
-22886 => x"C0C0BFA4A4808082",
-22885 => x"C0C0BFA4A4808092",
-22884 => x"C0C0BFA4A4808099",
-22883 => x"C0C0BFA4A48080B0",
-22882 => x"C0C0BFA4A48080A4",
-22881 => x"C0C0BFA4A48080F9",
-22880 => x"C0C0BFA4A48080C0",
-22879 => x"C0C0BFA4A480F890",
-22878 => x"C0C0BFA4A480F880",
-22877 => x"C0C0BFA4A480F8F8",
-22876 => x"C0C0BFA4A480F882",
-22875 => x"C0C0BFA4A480F892",
-22874 => x"C0C0BFA4A480F899",
-22873 => x"C0C0BFA4A480F8B0",
-22872 => x"C0C0BFA4A480F8A4",
-22871 => x"C0C0BFA4A480F8F9",
-22870 => x"C0C0BFA4A480F8C0",
-22869 => x"C0C0BFA4A4808290",
-22868 => x"C0C0BFA4A4808280",
-22867 => x"C0C0BFA4A48082F8",
-22866 => x"C0C0BFA4A4808282",
-22865 => x"C0C0BFA4A4808292",
-22864 => x"C0C0BFA4A4808299",
-22863 => x"C0C0BFA4A48082B0",
-22862 => x"C0C0BFA4A48082A4",
-22861 => x"C0C0BFA4A48082F9",
-22860 => x"C0C0BFA4A48082C0",
-22859 => x"C0C0BFA4A4809290",
-22858 => x"C0C0BFA4A4809280",
-22857 => x"C0C0BFA4A48092F8",
-22856 => x"C0C0BFA4A4809282",
-22855 => x"C0C0BFA4A4809292",
-22854 => x"C0C0BFA4A4809299",
-22853 => x"C0C0BFA4A48092B0",
-22852 => x"C0C0BFA4A48092A4",
-22851 => x"C0C0BFA4A48092F9",
-22850 => x"C0C0BFA4A48092C0",
-22849 => x"C0C0BFA4A4809990",
-22848 => x"C0C0BFA4A4809980",
-22847 => x"C0C0BFA4A48099F8",
-22846 => x"C0C0BFA4A4809982",
-22845 => x"C0C0BFA4A4809992",
-22844 => x"C0C0BFA4A4809999",
-22843 => x"C0C0BFA4A48099B0",
-22842 => x"C0C0BFA4A48099A4",
-22841 => x"C0C0BFA4A48099F9",
-22840 => x"C0C0BFA4A48099C0",
-22839 => x"C0C0BFA4A480B090",
-22838 => x"C0C0BFA4A480B080",
-22837 => x"C0C0BFA4A480B0F8",
-22836 => x"C0C0BFA4A480B082",
-22835 => x"C0C0BFA4A480B092",
-22834 => x"C0C0BFA4A480B099",
-22833 => x"C0C0BFA4A480B0B0",
-22832 => x"C0C0BFA4A480B0A4",
-22831 => x"C0C0BFA4A480B0F9",
-22830 => x"C0C0BFA4A480B0C0",
-22829 => x"C0C0BFA4A480A490",
-22828 => x"C0C0BFA4A480A480",
-22827 => x"C0C0BFA4A480A4F8",
-22826 => x"C0C0BFA4A480A482",
-22825 => x"C0C0BFA4A480A492",
-22824 => x"C0C0BFA4A480A499",
-22823 => x"C0C0BFA4A480A4B0",
-22822 => x"C0C0BFA4A480A4A4",
-22821 => x"C0C0BFA4A480A4F9",
-22820 => x"C0C0BFA4A480A4C0",
-22819 => x"C0C0BFA4A480F990",
-22818 => x"C0C0BFA4A480F980",
-22817 => x"C0C0BFA4A480F9F8",
-22816 => x"C0C0BFA4A480F982",
-22815 => x"C0C0BFA4A480F992",
-22814 => x"C0C0BFA4A480F999",
-22813 => x"C0C0BFA4A480F9B0",
-22812 => x"C0C0BFA4A480F9A4",
-22811 => x"C0C0BFA4A480F9F9",
-22810 => x"C0C0BFA4A480F9C0",
-22809 => x"C0C0BFA4A480C090",
-22808 => x"C0C0BFA4A480C080",
-22807 => x"C0C0BFA4A480C0F8",
-22806 => x"C0C0BFA4A480C082",
-22805 => x"C0C0BFA4A480C092",
-22804 => x"C0C0BFA4A480C099",
-22803 => x"C0C0BFA4A480C0B0",
-22802 => x"C0C0BFA4A480C0A4",
-22801 => x"C0C0BFA4A480C0F9",
-22800 => x"C0C0BFA4A480C0C0",
-22799 => x"C0C0BFA4A4F89090",
-22798 => x"C0C0BFA4A4F89080",
-22797 => x"C0C0BFA4A4F890F8",
-22796 => x"C0C0BFA4A4F89082",
-22795 => x"C0C0BFA4A4F89092",
-22794 => x"C0C0BFA4A4F89099",
-22793 => x"C0C0BFA4A4F890B0",
-22792 => x"C0C0BFA4A4F890A4",
-22791 => x"C0C0BFA4A4F890F9",
-22790 => x"C0C0BFA4A4F890C0",
-22789 => x"C0C0BFA4A4F88090",
-22788 => x"C0C0BFA4A4F88080",
-22787 => x"C0C0BFA4A4F880F8",
-22786 => x"C0C0BFA4A4F88082",
-22785 => x"C0C0BFA4A4F88092",
-22784 => x"C0C0BFA4A4F88099",
-22783 => x"C0C0BFA4A4F880B0",
-22782 => x"C0C0BFA4A4F880A4",
-22781 => x"C0C0BFA4A4F880F9",
-22780 => x"C0C0BFA4A4F880C0",
-22779 => x"C0C0BFA4A4F8F890",
-22778 => x"C0C0BFA4A4F8F880",
-22777 => x"C0C0BFA4A4F8F8F8",
-22776 => x"C0C0BFA4A4F8F882",
-22775 => x"C0C0BFA4A4F8F892",
-22774 => x"C0C0BFA4A4F8F899",
-22773 => x"C0C0BFA4A4F8F8B0",
-22772 => x"C0C0BFA4A4F8F8A4",
-22771 => x"C0C0BFA4A4F8F8F9",
-22770 => x"C0C0BFA4A4F8F8C0",
-22769 => x"C0C0BFA4A4F88290",
-22768 => x"C0C0BFA4A4F88280",
-22767 => x"C0C0BFA4A4F882F8",
-22766 => x"C0C0BFA4A4F88282",
-22765 => x"C0C0BFA4A4F88292",
-22764 => x"C0C0BFA4A4F88299",
-22763 => x"C0C0BFA4A4F882B0",
-22762 => x"C0C0BFA4A4F882A4",
-22761 => x"C0C0BFA4A4F882F9",
-22760 => x"C0C0BFA4A4F882C0",
-22759 => x"C0C0BFA4A4F89290",
-22758 => x"C0C0BFA4A4F89280",
-22757 => x"C0C0BFA4A4F892F8",
-22756 => x"C0C0BFA4A4F89282",
-22755 => x"C0C0BFA4A4F89292",
-22754 => x"C0C0BFA4A4F89299",
-22753 => x"C0C0BFA4A4F892B0",
-22752 => x"C0C0BFA4A4F892A4",
-22751 => x"C0C0BFA4A4F892F9",
-22750 => x"C0C0BFA4A4F892C0",
-22749 => x"C0C0BFA4A4F89990",
-22748 => x"C0C0BFA4A4F89980",
-22747 => x"C0C0BFA4A4F899F8",
-22746 => x"C0C0BFA4A4F89982",
-22745 => x"C0C0BFA4A4F89992",
-22744 => x"C0C0BFA4A4F89999",
-22743 => x"C0C0BFA4A4F899B0",
-22742 => x"C0C0BFA4A4F899A4",
-22741 => x"C0C0BFA4A4F899F9",
-22740 => x"C0C0BFA4A4F899C0",
-22739 => x"C0C0BFA4A4F8B090",
-22738 => x"C0C0BFA4A4F8B080",
-22737 => x"C0C0BFA4A4F8B0F8",
-22736 => x"C0C0BFA4A4F8B082",
-22735 => x"C0C0BFA4A4F8B092",
-22734 => x"C0C0BFA4A4F8B099",
-22733 => x"C0C0BFA4A4F8B0B0",
-22732 => x"C0C0BFA4A4F8B0A4",
-22731 => x"C0C0BFA4A4F8B0F9",
-22730 => x"C0C0BFA4A4F8B0C0",
-22729 => x"C0C0BFA4A4F8A490",
-22728 => x"C0C0BFA4A4F8A480",
-22727 => x"C0C0BFA4A4F8A4F8",
-22726 => x"C0C0BFA4A4F8A482",
-22725 => x"C0C0BFA4A4F8A492",
-22724 => x"C0C0BFA4A4F8A499",
-22723 => x"C0C0BFA4A4F8A4B0",
-22722 => x"C0C0BFA4A4F8A4A4",
-22721 => x"C0C0BFA4A4F8A4F9",
-22720 => x"C0C0BFA4A4F8A4C0",
-22719 => x"C0C0BFA4A4F8F990",
-22718 => x"C0C0BFA4A4F8F980",
-22717 => x"C0C0BFA4A4F8F9F8",
-22716 => x"C0C0BFA4A4F8F982",
-22715 => x"C0C0BFA4A4F8F992",
-22714 => x"C0C0BFA4A4F8F999",
-22713 => x"C0C0BFA4A4F8F9B0",
-22712 => x"C0C0BFA4A4F8F9A4",
-22711 => x"C0C0BFA4A4F8F9F9",
-22710 => x"C0C0BFA4A4F8F9C0",
-22709 => x"C0C0BFA4A4F8C090",
-22708 => x"C0C0BFA4A4F8C080",
-22707 => x"C0C0BFA4A4F8C0F8",
-22706 => x"C0C0BFA4A4F8C082",
-22705 => x"C0C0BFA4A4F8C092",
-22704 => x"C0C0BFA4A4F8C099",
-22703 => x"C0C0BFA4A4F8C0B0",
-22702 => x"C0C0BFA4A4F8C0A4",
-22701 => x"C0C0BFA4A4F8C0F9",
-22700 => x"C0C0BFA4A4F8C0C0",
-22699 => x"C0C0BFA4A4829090",
-22698 => x"C0C0BFA4A4829080",
-22697 => x"C0C0BFA4A48290F8",
-22696 => x"C0C0BFA4A4829082",
-22695 => x"C0C0BFA4A4829092",
-22694 => x"C0C0BFA4A4829099",
-22693 => x"C0C0BFA4A48290B0",
-22692 => x"C0C0BFA4A48290A4",
-22691 => x"C0C0BFA4A48290F9",
-22690 => x"C0C0BFA4A48290C0",
-22689 => x"C0C0BFA4A4828090",
-22688 => x"C0C0BFA4A4828080",
-22687 => x"C0C0BFA4A48280F8",
-22686 => x"C0C0BFA4A4828082",
-22685 => x"C0C0BFA4A4828092",
-22684 => x"C0C0BFA4A4828099",
-22683 => x"C0C0BFA4A48280B0",
-22682 => x"C0C0BFA4A48280A4",
-22681 => x"C0C0BFA4A48280F9",
-22680 => x"C0C0BFA4A48280C0",
-22679 => x"C0C0BFA4A482F890",
-22678 => x"C0C0BFA4A482F880",
-22677 => x"C0C0BFA4A482F8F8",
-22676 => x"C0C0BFA4A482F882",
-22675 => x"C0C0BFA4A482F892",
-22674 => x"C0C0BFA4A482F899",
-22673 => x"C0C0BFA4A482F8B0",
-22672 => x"C0C0BFA4A482F8A4",
-22671 => x"C0C0BFA4A482F8F9",
-22670 => x"C0C0BFA4A482F8C0",
-22669 => x"C0C0BFA4A4828290",
-22668 => x"C0C0BFA4A4828280",
-22667 => x"C0C0BFA4A48282F8",
-22666 => x"C0C0BFA4A4828282",
-22665 => x"C0C0BFA4A4828292",
-22664 => x"C0C0BFA4A4828299",
-22663 => x"C0C0BFA4A48282B0",
-22662 => x"C0C0BFA4A48282A4",
-22661 => x"C0C0BFA4A48282F9",
-22660 => x"C0C0BFA4A48282C0",
-22659 => x"C0C0BFA4A4829290",
-22658 => x"C0C0BFA4A4829280",
-22657 => x"C0C0BFA4A48292F8",
-22656 => x"C0C0BFA4A4829282",
-22655 => x"C0C0BFA4A4829292",
-22654 => x"C0C0BFA4A4829299",
-22653 => x"C0C0BFA4A48292B0",
-22652 => x"C0C0BFA4A48292A4",
-22651 => x"C0C0BFA4A48292F9",
-22650 => x"C0C0BFA4A48292C0",
-22649 => x"C0C0BFA4A4829990",
-22648 => x"C0C0BFA4A4829980",
-22647 => x"C0C0BFA4A48299F8",
-22646 => x"C0C0BFA4A4829982",
-22645 => x"C0C0BFA4A4829992",
-22644 => x"C0C0BFA4A4829999",
-22643 => x"C0C0BFA4A48299B0",
-22642 => x"C0C0BFA4A48299A4",
-22641 => x"C0C0BFA4A48299F9",
-22640 => x"C0C0BFA4A48299C0",
-22639 => x"C0C0BFA4A482B090",
-22638 => x"C0C0BFA4A482B080",
-22637 => x"C0C0BFA4A482B0F8",
-22636 => x"C0C0BFA4A482B082",
-22635 => x"C0C0BFA4A482B092",
-22634 => x"C0C0BFA4A482B099",
-22633 => x"C0C0BFA4A482B0B0",
-22632 => x"C0C0BFA4A482B0A4",
-22631 => x"C0C0BFA4A482B0F9",
-22630 => x"C0C0BFA4A482B0C0",
-22629 => x"C0C0BFA4A482A490",
-22628 => x"C0C0BFA4A482A480",
-22627 => x"C0C0BFA4A482A4F8",
-22626 => x"C0C0BFA4A482A482",
-22625 => x"C0C0BFA4A482A492",
-22624 => x"C0C0BFA4A482A499",
-22623 => x"C0C0BFA4A482A4B0",
-22622 => x"C0C0BFA4A482A4A4",
-22621 => x"C0C0BFA4A482A4F9",
-22620 => x"C0C0BFA4A482A4C0",
-22619 => x"C0C0BFA4A482F990",
-22618 => x"C0C0BFA4A482F980",
-22617 => x"C0C0BFA4A482F9F8",
-22616 => x"C0C0BFA4A482F982",
-22615 => x"C0C0BFA4A482F992",
-22614 => x"C0C0BFA4A482F999",
-22613 => x"C0C0BFA4A482F9B0",
-22612 => x"C0C0BFA4A482F9A4",
-22611 => x"C0C0BFA4A482F9F9",
-22610 => x"C0C0BFA4A482F9C0",
-22609 => x"C0C0BFA4A482C090",
-22608 => x"C0C0BFA4A482C080",
-22607 => x"C0C0BFA4A482C0F8",
-22606 => x"C0C0BFA4A482C082",
-22605 => x"C0C0BFA4A482C092",
-22604 => x"C0C0BFA4A482C099",
-22603 => x"C0C0BFA4A482C0B0",
-22602 => x"C0C0BFA4A482C0A4",
-22601 => x"C0C0BFA4A482C0F9",
-22600 => x"C0C0BFA4A482C0C0",
-22599 => x"C0C0BFA4A4929090",
-22598 => x"C0C0BFA4A4929080",
-22597 => x"C0C0BFA4A49290F8",
-22596 => x"C0C0BFA4A4929082",
-22595 => x"C0C0BFA4A4929092",
-22594 => x"C0C0BFA4A4929099",
-22593 => x"C0C0BFA4A49290B0",
-22592 => x"C0C0BFA4A49290A4",
-22591 => x"C0C0BFA4A49290F9",
-22590 => x"C0C0BFA4A49290C0",
-22589 => x"C0C0BFA4A4928090",
-22588 => x"C0C0BFA4A4928080",
-22587 => x"C0C0BFA4A49280F8",
-22586 => x"C0C0BFA4A4928082",
-22585 => x"C0C0BFA4A4928092",
-22584 => x"C0C0BFA4A4928099",
-22583 => x"C0C0BFA4A49280B0",
-22582 => x"C0C0BFA4A49280A4",
-22581 => x"C0C0BFA4A49280F9",
-22580 => x"C0C0BFA4A49280C0",
-22579 => x"C0C0BFA4A492F890",
-22578 => x"C0C0BFA4A492F880",
-22577 => x"C0C0BFA4A492F8F8",
-22576 => x"C0C0BFA4A492F882",
-22575 => x"C0C0BFA4A492F892",
-22574 => x"C0C0BFA4A492F899",
-22573 => x"C0C0BFA4A492F8B0",
-22572 => x"C0C0BFA4A492F8A4",
-22571 => x"C0C0BFA4A492F8F9",
-22570 => x"C0C0BFA4A492F8C0",
-22569 => x"C0C0BFA4A4928290",
-22568 => x"C0C0BFA4A4928280",
-22567 => x"C0C0BFA4A49282F8",
-22566 => x"C0C0BFA4A4928282",
-22565 => x"C0C0BFA4A4928292",
-22564 => x"C0C0BFA4A4928299",
-22563 => x"C0C0BFA4A49282B0",
-22562 => x"C0C0BFA4A49282A4",
-22561 => x"C0C0BFA4A49282F9",
-22560 => x"C0C0BFA4A49282C0",
-22559 => x"C0C0BFA4A4929290",
-22558 => x"C0C0BFA4A4929280",
-22557 => x"C0C0BFA4A49292F8",
-22556 => x"C0C0BFA4A4929282",
-22555 => x"C0C0BFA4A4929292",
-22554 => x"C0C0BFA4A4929299",
-22553 => x"C0C0BFA4A49292B0",
-22552 => x"C0C0BFA4A49292A4",
-22551 => x"C0C0BFA4A49292F9",
-22550 => x"C0C0BFA4A49292C0",
-22549 => x"C0C0BFA4A4929990",
-22548 => x"C0C0BFA4A4929980",
-22547 => x"C0C0BFA4A49299F8",
-22546 => x"C0C0BFA4A4929982",
-22545 => x"C0C0BFA4A4929992",
-22544 => x"C0C0BFA4A4929999",
-22543 => x"C0C0BFA4A49299B0",
-22542 => x"C0C0BFA4A49299A4",
-22541 => x"C0C0BFA4A49299F9",
-22540 => x"C0C0BFA4A49299C0",
-22539 => x"C0C0BFA4A492B090",
-22538 => x"C0C0BFA4A492B080",
-22537 => x"C0C0BFA4A492B0F8",
-22536 => x"C0C0BFA4A492B082",
-22535 => x"C0C0BFA4A492B092",
-22534 => x"C0C0BFA4A492B099",
-22533 => x"C0C0BFA4A492B0B0",
-22532 => x"C0C0BFA4A492B0A4",
-22531 => x"C0C0BFA4A492B0F9",
-22530 => x"C0C0BFA4A492B0C0",
-22529 => x"C0C0BFA4A492A490",
-22528 => x"C0C0BFA4A492A480",
-22527 => x"C0C0BFA4A492A4F8",
-22526 => x"C0C0BFA4A492A482",
-22525 => x"C0C0BFA4A492A492",
-22524 => x"C0C0BFA4A492A499",
-22523 => x"C0C0BFA4A492A4B0",
-22522 => x"C0C0BFA4A492A4A4",
-22521 => x"C0C0BFA4A492A4F9",
-22520 => x"C0C0BFA4A492A4C0",
-22519 => x"C0C0BFA4A492F990",
-22518 => x"C0C0BFA4A492F980",
-22517 => x"C0C0BFA4A492F9F8",
-22516 => x"C0C0BFA4A492F982",
-22515 => x"C0C0BFA4A492F992",
-22514 => x"C0C0BFA4A492F999",
-22513 => x"C0C0BFA4A492F9B0",
-22512 => x"C0C0BFA4A492F9A4",
-22511 => x"C0C0BFA4A492F9F9",
-22510 => x"C0C0BFA4A492F9C0",
-22509 => x"C0C0BFA4A492C090",
-22508 => x"C0C0BFA4A492C080",
-22507 => x"C0C0BFA4A492C0F8",
-22506 => x"C0C0BFA4A492C082",
-22505 => x"C0C0BFA4A492C092",
-22504 => x"C0C0BFA4A492C099",
-22503 => x"C0C0BFA4A492C0B0",
-22502 => x"C0C0BFA4A492C0A4",
-22501 => x"C0C0BFA4A492C0F9",
-22500 => x"C0C0BFA4A492C0C0",
-22499 => x"C0C0BFA4A4999090",
-22498 => x"C0C0BFA4A4999080",
-22497 => x"C0C0BFA4A49990F8",
-22496 => x"C0C0BFA4A4999082",
-22495 => x"C0C0BFA4A4999092",
-22494 => x"C0C0BFA4A4999099",
-22493 => x"C0C0BFA4A49990B0",
-22492 => x"C0C0BFA4A49990A4",
-22491 => x"C0C0BFA4A49990F9",
-22490 => x"C0C0BFA4A49990C0",
-22489 => x"C0C0BFA4A4998090",
-22488 => x"C0C0BFA4A4998080",
-22487 => x"C0C0BFA4A49980F8",
-22486 => x"C0C0BFA4A4998082",
-22485 => x"C0C0BFA4A4998092",
-22484 => x"C0C0BFA4A4998099",
-22483 => x"C0C0BFA4A49980B0",
-22482 => x"C0C0BFA4A49980A4",
-22481 => x"C0C0BFA4A49980F9",
-22480 => x"C0C0BFA4A49980C0",
-22479 => x"C0C0BFA4A499F890",
-22478 => x"C0C0BFA4A499F880",
-22477 => x"C0C0BFA4A499F8F8",
-22476 => x"C0C0BFA4A499F882",
-22475 => x"C0C0BFA4A499F892",
-22474 => x"C0C0BFA4A499F899",
-22473 => x"C0C0BFA4A499F8B0",
-22472 => x"C0C0BFA4A499F8A4",
-22471 => x"C0C0BFA4A499F8F9",
-22470 => x"C0C0BFA4A499F8C0",
-22469 => x"C0C0BFA4A4998290",
-22468 => x"C0C0BFA4A4998280",
-22467 => x"C0C0BFA4A49982F8",
-22466 => x"C0C0BFA4A4998282",
-22465 => x"C0C0BFA4A4998292",
-22464 => x"C0C0BFA4A4998299",
-22463 => x"C0C0BFA4A49982B0",
-22462 => x"C0C0BFA4A49982A4",
-22461 => x"C0C0BFA4A49982F9",
-22460 => x"C0C0BFA4A49982C0",
-22459 => x"C0C0BFA4A4999290",
-22458 => x"C0C0BFA4A4999280",
-22457 => x"C0C0BFA4A49992F8",
-22456 => x"C0C0BFA4A4999282",
-22455 => x"C0C0BFA4A4999292",
-22454 => x"C0C0BFA4A4999299",
-22453 => x"C0C0BFA4A49992B0",
-22452 => x"C0C0BFA4A49992A4",
-22451 => x"C0C0BFA4A49992F9",
-22450 => x"C0C0BFA4A49992C0",
-22449 => x"C0C0BFA4A4999990",
-22448 => x"C0C0BFA4A4999980",
-22447 => x"C0C0BFA4A49999F8",
-22446 => x"C0C0BFA4A4999982",
-22445 => x"C0C0BFA4A4999992",
-22444 => x"C0C0BFA4A4999999",
-22443 => x"C0C0BFA4A49999B0",
-22442 => x"C0C0BFA4A49999A4",
-22441 => x"C0C0BFA4A49999F9",
-22440 => x"C0C0BFA4A49999C0",
-22439 => x"C0C0BFA4A499B090",
-22438 => x"C0C0BFA4A499B080",
-22437 => x"C0C0BFA4A499B0F8",
-22436 => x"C0C0BFA4A499B082",
-22435 => x"C0C0BFA4A499B092",
-22434 => x"C0C0BFA4A499B099",
-22433 => x"C0C0BFA4A499B0B0",
-22432 => x"C0C0BFA4A499B0A4",
-22431 => x"C0C0BFA4A499B0F9",
-22430 => x"C0C0BFA4A499B0C0",
-22429 => x"C0C0BFA4A499A490",
-22428 => x"C0C0BFA4A499A480",
-22427 => x"C0C0BFA4A499A4F8",
-22426 => x"C0C0BFA4A499A482",
-22425 => x"C0C0BFA4A499A492",
-22424 => x"C0C0BFA4A499A499",
-22423 => x"C0C0BFA4A499A4B0",
-22422 => x"C0C0BFA4A499A4A4",
-22421 => x"C0C0BFA4A499A4F9",
-22420 => x"C0C0BFA4A499A4C0",
-22419 => x"C0C0BFA4A499F990",
-22418 => x"C0C0BFA4A499F980",
-22417 => x"C0C0BFA4A499F9F8",
-22416 => x"C0C0BFA4A499F982",
-22415 => x"C0C0BFA4A499F992",
-22414 => x"C0C0BFA4A499F999",
-22413 => x"C0C0BFA4A499F9B0",
-22412 => x"C0C0BFA4A499F9A4",
-22411 => x"C0C0BFA4A499F9F9",
-22410 => x"C0C0BFA4A499F9C0",
-22409 => x"C0C0BFA4A499C090",
-22408 => x"C0C0BFA4A499C080",
-22407 => x"C0C0BFA4A499C0F8",
-22406 => x"C0C0BFA4A499C082",
-22405 => x"C0C0BFA4A499C092",
-22404 => x"C0C0BFA4A499C099",
-22403 => x"C0C0BFA4A499C0B0",
-22402 => x"C0C0BFA4A499C0A4",
-22401 => x"C0C0BFA4A499C0F9",
-22400 => x"C0C0BFA4A499C0C0",
-22399 => x"C0C0BFA4A4B09090",
-22398 => x"C0C0BFA4A4B09080",
-22397 => x"C0C0BFA4A4B090F8",
-22396 => x"C0C0BFA4A4B09082",
-22395 => x"C0C0BFA4A4B09092",
-22394 => x"C0C0BFA4A4B09099",
-22393 => x"C0C0BFA4A4B090B0",
-22392 => x"C0C0BFA4A4B090A4",
-22391 => x"C0C0BFA4A4B090F9",
-22390 => x"C0C0BFA4A4B090C0",
-22389 => x"C0C0BFA4A4B08090",
-22388 => x"C0C0BFA4A4B08080",
-22387 => x"C0C0BFA4A4B080F8",
-22386 => x"C0C0BFA4A4B08082",
-22385 => x"C0C0BFA4A4B08092",
-22384 => x"C0C0BFA4A4B08099",
-22383 => x"C0C0BFA4A4B080B0",
-22382 => x"C0C0BFA4A4B080A4",
-22381 => x"C0C0BFA4A4B080F9",
-22380 => x"C0C0BFA4A4B080C0",
-22379 => x"C0C0BFA4A4B0F890",
-22378 => x"C0C0BFA4A4B0F880",
-22377 => x"C0C0BFA4A4B0F8F8",
-22376 => x"C0C0BFA4A4B0F882",
-22375 => x"C0C0BFA4A4B0F892",
-22374 => x"C0C0BFA4A4B0F899",
-22373 => x"C0C0BFA4A4B0F8B0",
-22372 => x"C0C0BFA4A4B0F8A4",
-22371 => x"C0C0BFA4A4B0F8F9",
-22370 => x"C0C0BFA4A4B0F8C0",
-22369 => x"C0C0BFA4A4B08290",
-22368 => x"C0C0BFA4A4B08280",
-22367 => x"C0C0BFA4A4B082F8",
-22366 => x"C0C0BFA4A4B08282",
-22365 => x"C0C0BFA4A4B08292",
-22364 => x"C0C0BFA4A4B08299",
-22363 => x"C0C0BFA4A4B082B0",
-22362 => x"C0C0BFA4A4B082A4",
-22361 => x"C0C0BFA4A4B082F9",
-22360 => x"C0C0BFA4A4B082C0",
-22359 => x"C0C0BFA4A4B09290",
-22358 => x"C0C0BFA4A4B09280",
-22357 => x"C0C0BFA4A4B092F8",
-22356 => x"C0C0BFA4A4B09282",
-22355 => x"C0C0BFA4A4B09292",
-22354 => x"C0C0BFA4A4B09299",
-22353 => x"C0C0BFA4A4B092B0",
-22352 => x"C0C0BFA4A4B092A4",
-22351 => x"C0C0BFA4A4B092F9",
-22350 => x"C0C0BFA4A4B092C0",
-22349 => x"C0C0BFA4A4B09990",
-22348 => x"C0C0BFA4A4B09980",
-22347 => x"C0C0BFA4A4B099F8",
-22346 => x"C0C0BFA4A4B09982",
-22345 => x"C0C0BFA4A4B09992",
-22344 => x"C0C0BFA4A4B09999",
-22343 => x"C0C0BFA4A4B099B0",
-22342 => x"C0C0BFA4A4B099A4",
-22341 => x"C0C0BFA4A4B099F9",
-22340 => x"C0C0BFA4A4B099C0",
-22339 => x"C0C0BFA4A4B0B090",
-22338 => x"C0C0BFA4A4B0B080",
-22337 => x"C0C0BFA4A4B0B0F8",
-22336 => x"C0C0BFA4A4B0B082",
-22335 => x"C0C0BFA4A4B0B092",
-22334 => x"C0C0BFA4A4B0B099",
-22333 => x"C0C0BFA4A4B0B0B0",
-22332 => x"C0C0BFA4A4B0B0A4",
-22331 => x"C0C0BFA4A4B0B0F9",
-22330 => x"C0C0BFA4A4B0B0C0",
-22329 => x"C0C0BFA4A4B0A490",
-22328 => x"C0C0BFA4A4B0A480",
-22327 => x"C0C0BFA4A4B0A4F8",
-22326 => x"C0C0BFA4A4B0A482",
-22325 => x"C0C0BFA4A4B0A492",
-22324 => x"C0C0BFA4A4B0A499",
-22323 => x"C0C0BFA4A4B0A4B0",
-22322 => x"C0C0BFA4A4B0A4A4",
-22321 => x"C0C0BFA4A4B0A4F9",
-22320 => x"C0C0BFA4A4B0A4C0",
-22319 => x"C0C0BFA4A4B0F990",
-22318 => x"C0C0BFA4A4B0F980",
-22317 => x"C0C0BFA4A4B0F9F8",
-22316 => x"C0C0BFA4A4B0F982",
-22315 => x"C0C0BFA4A4B0F992",
-22314 => x"C0C0BFA4A4B0F999",
-22313 => x"C0C0BFA4A4B0F9B0",
-22312 => x"C0C0BFA4A4B0F9A4",
-22311 => x"C0C0BFA4A4B0F9F9",
-22310 => x"C0C0BFA4A4B0F9C0",
-22309 => x"C0C0BFA4A4B0C090",
-22308 => x"C0C0BFA4A4B0C080",
-22307 => x"C0C0BFA4A4B0C0F8",
-22306 => x"C0C0BFA4A4B0C082",
-22305 => x"C0C0BFA4A4B0C092",
-22304 => x"C0C0BFA4A4B0C099",
-22303 => x"C0C0BFA4A4B0C0B0",
-22302 => x"C0C0BFA4A4B0C0A4",
-22301 => x"C0C0BFA4A4B0C0F9",
-22300 => x"C0C0BFA4A4B0C0C0",
-22299 => x"C0C0BFA4A4A49090",
-22298 => x"C0C0BFA4A4A49080",
-22297 => x"C0C0BFA4A4A490F8",
-22296 => x"C0C0BFA4A4A49082",
-22295 => x"C0C0BFA4A4A49092",
-22294 => x"C0C0BFA4A4A49099",
-22293 => x"C0C0BFA4A4A490B0",
-22292 => x"C0C0BFA4A4A490A4",
-22291 => x"C0C0BFA4A4A490F9",
-22290 => x"C0C0BFA4A4A490C0",
-22289 => x"C0C0BFA4A4A48090",
-22288 => x"C0C0BFA4A4A48080",
-22287 => x"C0C0BFA4A4A480F8",
-22286 => x"C0C0BFA4A4A48082",
-22285 => x"C0C0BFA4A4A48092",
-22284 => x"C0C0BFA4A4A48099",
-22283 => x"C0C0BFA4A4A480B0",
-22282 => x"C0C0BFA4A4A480A4",
-22281 => x"C0C0BFA4A4A480F9",
-22280 => x"C0C0BFA4A4A480C0",
-22279 => x"C0C0BFA4A4A4F890",
-22278 => x"C0C0BFA4A4A4F880",
-22277 => x"C0C0BFA4A4A4F8F8",
-22276 => x"C0C0BFA4A4A4F882",
-22275 => x"C0C0BFA4A4A4F892",
-22274 => x"C0C0BFA4A4A4F899",
-22273 => x"C0C0BFA4A4A4F8B0",
-22272 => x"C0C0BFA4A4A4F8A4",
-22271 => x"C0C0BFA4A4A4F8F9",
-22270 => x"C0C0BFA4A4A4F8C0",
-22269 => x"C0C0BFA4A4A48290",
-22268 => x"C0C0BFA4A4A48280",
-22267 => x"C0C0BFA4A4A482F8",
-22266 => x"C0C0BFA4A4A48282",
-22265 => x"C0C0BFA4A4A48292",
-22264 => x"C0C0BFA4A4A48299",
-22263 => x"C0C0BFA4A4A482B0",
-22262 => x"C0C0BFA4A4A482A4",
-22261 => x"C0C0BFA4A4A482F9",
-22260 => x"C0C0BFA4A4A482C0",
-22259 => x"C0C0BFA4A4A49290",
-22258 => x"C0C0BFA4A4A49280",
-22257 => x"C0C0BFA4A4A492F8",
-22256 => x"C0C0BFA4A4A49282",
-22255 => x"C0C0BFA4A4A49292",
-22254 => x"C0C0BFA4A4A49299",
-22253 => x"C0C0BFA4A4A492B0",
-22252 => x"C0C0BFA4A4A492A4",
-22251 => x"C0C0BFA4A4A492F9",
-22250 => x"C0C0BFA4A4A492C0",
-22249 => x"C0C0BFA4A4A49990",
-22248 => x"C0C0BFA4A4A49980",
-22247 => x"C0C0BFA4A4A499F8",
-22246 => x"C0C0BFA4A4A49982",
-22245 => x"C0C0BFA4A4A49992",
-22244 => x"C0C0BFA4A4A49999",
-22243 => x"C0C0BFA4A4A499B0",
-22242 => x"C0C0BFA4A4A499A4",
-22241 => x"C0C0BFA4A4A499F9",
-22240 => x"C0C0BFA4A4A499C0",
-22239 => x"C0C0BFA4A4A4B090",
-22238 => x"C0C0BFA4A4A4B080",
-22237 => x"C0C0BFA4A4A4B0F8",
-22236 => x"C0C0BFA4A4A4B082",
-22235 => x"C0C0BFA4A4A4B092",
-22234 => x"C0C0BFA4A4A4B099",
-22233 => x"C0C0BFA4A4A4B0B0",
-22232 => x"C0C0BFA4A4A4B0A4",
-22231 => x"C0C0BFA4A4A4B0F9",
-22230 => x"C0C0BFA4A4A4B0C0",
-22229 => x"C0C0BFA4A4A4A490",
-22228 => x"C0C0BFA4A4A4A480",
-22227 => x"C0C0BFA4A4A4A4F8",
-22226 => x"C0C0BFA4A4A4A482",
-22225 => x"C0C0BFA4A4A4A492",
-22224 => x"C0C0BFA4A4A4A499",
-22223 => x"C0C0BFA4A4A4A4B0",
-22222 => x"C0C0BFA4A4A4A4A4",
-22221 => x"C0C0BFA4A4A4A4F9",
-22220 => x"C0C0BFA4A4A4A4C0",
-22219 => x"C0C0BFA4A4A4F990",
-22218 => x"C0C0BFA4A4A4F980",
-22217 => x"C0C0BFA4A4A4F9F8",
-22216 => x"C0C0BFA4A4A4F982",
-22215 => x"C0C0BFA4A4A4F992",
-22214 => x"C0C0BFA4A4A4F999",
-22213 => x"C0C0BFA4A4A4F9B0",
-22212 => x"C0C0BFA4A4A4F9A4",
-22211 => x"C0C0BFA4A4A4F9F9",
-22210 => x"C0C0BFA4A4A4F9C0",
-22209 => x"C0C0BFA4A4A4C090",
-22208 => x"C0C0BFA4A4A4C080",
-22207 => x"C0C0BFA4A4A4C0F8",
-22206 => x"C0C0BFA4A4A4C082",
-22205 => x"C0C0BFA4A4A4C092",
-22204 => x"C0C0BFA4A4A4C099",
-22203 => x"C0C0BFA4A4A4C0B0",
-22202 => x"C0C0BFA4A4A4C0A4",
-22201 => x"C0C0BFA4A4A4C0F9",
-22200 => x"C0C0BFA4A4A4C0C0",
-22199 => x"C0C0BFA4A4F99090",
-22198 => x"C0C0BFA4A4F99080",
-22197 => x"C0C0BFA4A4F990F8",
-22196 => x"C0C0BFA4A4F99082",
-22195 => x"C0C0BFA4A4F99092",
-22194 => x"C0C0BFA4A4F99099",
-22193 => x"C0C0BFA4A4F990B0",
-22192 => x"C0C0BFA4A4F990A4",
-22191 => x"C0C0BFA4A4F990F9",
-22190 => x"C0C0BFA4A4F990C0",
-22189 => x"C0C0BFA4A4F98090",
-22188 => x"C0C0BFA4A4F98080",
-22187 => x"C0C0BFA4A4F980F8",
-22186 => x"C0C0BFA4A4F98082",
-22185 => x"C0C0BFA4A4F98092",
-22184 => x"C0C0BFA4A4F98099",
-22183 => x"C0C0BFA4A4F980B0",
-22182 => x"C0C0BFA4A4F980A4",
-22181 => x"C0C0BFA4A4F980F9",
-22180 => x"C0C0BFA4A4F980C0",
-22179 => x"C0C0BFA4A4F9F890",
-22178 => x"C0C0BFA4A4F9F880",
-22177 => x"C0C0BFA4A4F9F8F8",
-22176 => x"C0C0BFA4A4F9F882",
-22175 => x"C0C0BFA4A4F9F892",
-22174 => x"C0C0BFA4A4F9F899",
-22173 => x"C0C0BFA4A4F9F8B0",
-22172 => x"C0C0BFA4A4F9F8A4",
-22171 => x"C0C0BFA4A4F9F8F9",
-22170 => x"C0C0BFA4A4F9F8C0",
-22169 => x"C0C0BFA4A4F98290",
-22168 => x"C0C0BFA4A4F98280",
-22167 => x"C0C0BFA4A4F982F8",
-22166 => x"C0C0BFA4A4F98282",
-22165 => x"C0C0BFA4A4F98292",
-22164 => x"C0C0BFA4A4F98299",
-22163 => x"C0C0BFA4A4F982B0",
-22162 => x"C0C0BFA4A4F982A4",
-22161 => x"C0C0BFA4A4F982F9",
-22160 => x"C0C0BFA4A4F982C0",
-22159 => x"C0C0BFA4A4F99290",
-22158 => x"C0C0BFA4A4F99280",
-22157 => x"C0C0BFA4A4F992F8",
-22156 => x"C0C0BFA4A4F99282",
-22155 => x"C0C0BFA4A4F99292",
-22154 => x"C0C0BFA4A4F99299",
-22153 => x"C0C0BFA4A4F992B0",
-22152 => x"C0C0BFA4A4F992A4",
-22151 => x"C0C0BFA4A4F992F9",
-22150 => x"C0C0BFA4A4F992C0",
-22149 => x"C0C0BFA4A4F99990",
-22148 => x"C0C0BFA4A4F99980",
-22147 => x"C0C0BFA4A4F999F8",
-22146 => x"C0C0BFA4A4F99982",
-22145 => x"C0C0BFA4A4F99992",
-22144 => x"C0C0BFA4A4F99999",
-22143 => x"C0C0BFA4A4F999B0",
-22142 => x"C0C0BFA4A4F999A4",
-22141 => x"C0C0BFA4A4F999F9",
-22140 => x"C0C0BFA4A4F999C0",
-22139 => x"C0C0BFA4A4F9B090",
-22138 => x"C0C0BFA4A4F9B080",
-22137 => x"C0C0BFA4A4F9B0F8",
-22136 => x"C0C0BFA4A4F9B082",
-22135 => x"C0C0BFA4A4F9B092",
-22134 => x"C0C0BFA4A4F9B099",
-22133 => x"C0C0BFA4A4F9B0B0",
-22132 => x"C0C0BFA4A4F9B0A4",
-22131 => x"C0C0BFA4A4F9B0F9",
-22130 => x"C0C0BFA4A4F9B0C0",
-22129 => x"C0C0BFA4A4F9A490",
-22128 => x"C0C0BFA4A4F9A480",
-22127 => x"C0C0BFA4A4F9A4F8",
-22126 => x"C0C0BFA4A4F9A482",
-22125 => x"C0C0BFA4A4F9A492",
-22124 => x"C0C0BFA4A4F9A499",
-22123 => x"C0C0BFA4A4F9A4B0",
-22122 => x"C0C0BFA4A4F9A4A4",
-22121 => x"C0C0BFA4A4F9A4F9",
-22120 => x"C0C0BFA4A4F9A4C0",
-22119 => x"C0C0BFA4A4F9F990",
-22118 => x"C0C0BFA4A4F9F980",
-22117 => x"C0C0BFA4A4F9F9F8",
-22116 => x"C0C0BFA4A4F9F982",
-22115 => x"C0C0BFA4A4F9F992",
-22114 => x"C0C0BFA4A4F9F999",
-22113 => x"C0C0BFA4A4F9F9B0",
-22112 => x"C0C0BFA4A4F9F9A4",
-22111 => x"C0C0BFA4A4F9F9F9",
-22110 => x"C0C0BFA4A4F9F9C0",
-22109 => x"C0C0BFA4A4F9C090",
-22108 => x"C0C0BFA4A4F9C080",
-22107 => x"C0C0BFA4A4F9C0F8",
-22106 => x"C0C0BFA4A4F9C082",
-22105 => x"C0C0BFA4A4F9C092",
-22104 => x"C0C0BFA4A4F9C099",
-22103 => x"C0C0BFA4A4F9C0B0",
-22102 => x"C0C0BFA4A4F9C0A4",
-22101 => x"C0C0BFA4A4F9C0F9",
-22100 => x"C0C0BFA4A4F9C0C0",
-22099 => x"C0C0BFA4A4C09090",
-22098 => x"C0C0BFA4A4C09080",
-22097 => x"C0C0BFA4A4C090F8",
-22096 => x"C0C0BFA4A4C09082",
-22095 => x"C0C0BFA4A4C09092",
-22094 => x"C0C0BFA4A4C09099",
-22093 => x"C0C0BFA4A4C090B0",
-22092 => x"C0C0BFA4A4C090A4",
-22091 => x"C0C0BFA4A4C090F9",
-22090 => x"C0C0BFA4A4C090C0",
-22089 => x"C0C0BFA4A4C08090",
-22088 => x"C0C0BFA4A4C08080",
-22087 => x"C0C0BFA4A4C080F8",
-22086 => x"C0C0BFA4A4C08082",
-22085 => x"C0C0BFA4A4C08092",
-22084 => x"C0C0BFA4A4C08099",
-22083 => x"C0C0BFA4A4C080B0",
-22082 => x"C0C0BFA4A4C080A4",
-22081 => x"C0C0BFA4A4C080F9",
-22080 => x"C0C0BFA4A4C080C0",
-22079 => x"C0C0BFA4A4C0F890",
-22078 => x"C0C0BFA4A4C0F880",
-22077 => x"C0C0BFA4A4C0F8F8",
-22076 => x"C0C0BFA4A4C0F882",
-22075 => x"C0C0BFA4A4C0F892",
-22074 => x"C0C0BFA4A4C0F899",
-22073 => x"C0C0BFA4A4C0F8B0",
-22072 => x"C0C0BFA4A4C0F8A4",
-22071 => x"C0C0BFA4A4C0F8F9",
-22070 => x"C0C0BFA4A4C0F8C0",
-22069 => x"C0C0BFA4A4C08290",
-22068 => x"C0C0BFA4A4C08280",
-22067 => x"C0C0BFA4A4C082F8",
-22066 => x"C0C0BFA4A4C08282",
-22065 => x"C0C0BFA4A4C08292",
-22064 => x"C0C0BFA4A4C08299",
-22063 => x"C0C0BFA4A4C082B0",
-22062 => x"C0C0BFA4A4C082A4",
-22061 => x"C0C0BFA4A4C082F9",
-22060 => x"C0C0BFA4A4C082C0",
-22059 => x"C0C0BFA4A4C09290",
-22058 => x"C0C0BFA4A4C09280",
-22057 => x"C0C0BFA4A4C092F8",
-22056 => x"C0C0BFA4A4C09282",
-22055 => x"C0C0BFA4A4C09292",
-22054 => x"C0C0BFA4A4C09299",
-22053 => x"C0C0BFA4A4C092B0",
-22052 => x"C0C0BFA4A4C092A4",
-22051 => x"C0C0BFA4A4C092F9",
-22050 => x"C0C0BFA4A4C092C0",
-22049 => x"C0C0BFA4A4C09990",
-22048 => x"C0C0BFA4A4C09980",
-22047 => x"C0C0BFA4A4C099F8",
-22046 => x"C0C0BFA4A4C09982",
-22045 => x"C0C0BFA4A4C09992",
-22044 => x"C0C0BFA4A4C09999",
-22043 => x"C0C0BFA4A4C099B0",
-22042 => x"C0C0BFA4A4C099A4",
-22041 => x"C0C0BFA4A4C099F9",
-22040 => x"C0C0BFA4A4C099C0",
-22039 => x"C0C0BFA4A4C0B090",
-22038 => x"C0C0BFA4A4C0B080",
-22037 => x"C0C0BFA4A4C0B0F8",
-22036 => x"C0C0BFA4A4C0B082",
-22035 => x"C0C0BFA4A4C0B092",
-22034 => x"C0C0BFA4A4C0B099",
-22033 => x"C0C0BFA4A4C0B0B0",
-22032 => x"C0C0BFA4A4C0B0A4",
-22031 => x"C0C0BFA4A4C0B0F9",
-22030 => x"C0C0BFA4A4C0B0C0",
-22029 => x"C0C0BFA4A4C0A490",
-22028 => x"C0C0BFA4A4C0A480",
-22027 => x"C0C0BFA4A4C0A4F8",
-22026 => x"C0C0BFA4A4C0A482",
-22025 => x"C0C0BFA4A4C0A492",
-22024 => x"C0C0BFA4A4C0A499",
-22023 => x"C0C0BFA4A4C0A4B0",
-22022 => x"C0C0BFA4A4C0A4A4",
-22021 => x"C0C0BFA4A4C0A4F9",
-22020 => x"C0C0BFA4A4C0A4C0",
-22019 => x"C0C0BFA4A4C0F990",
-22018 => x"C0C0BFA4A4C0F980",
-22017 => x"C0C0BFA4A4C0F9F8",
-22016 => x"C0C0BFA4A4C0F982",
-22015 => x"C0C0BFA4A4C0F992",
-22014 => x"C0C0BFA4A4C0F999",
-22013 => x"C0C0BFA4A4C0F9B0",
-22012 => x"C0C0BFA4A4C0F9A4",
-22011 => x"C0C0BFA4A4C0F9F9",
-22010 => x"C0C0BFA4A4C0F9C0",
-22009 => x"C0C0BFA4A4C0C090",
-22008 => x"C0C0BFA4A4C0C080",
-22007 => x"C0C0BFA4A4C0C0F8",
-22006 => x"C0C0BFA4A4C0C082",
-22005 => x"C0C0BFA4A4C0C092",
-22004 => x"C0C0BFA4A4C0C099",
-22003 => x"C0C0BFA4A4C0C0B0",
-22002 => x"C0C0BFA4A4C0C0A4",
-22001 => x"C0C0BFA4A4C0C0F9",
-22000 => x"C0C0BFA4A4C0C0C0",
-21999 => x"C0C0BFA4F9909090",
-21998 => x"C0C0BFA4F9909080",
-21997 => x"C0C0BFA4F99090F8",
-21996 => x"C0C0BFA4F9909082",
-21995 => x"C0C0BFA4F9909092",
-21994 => x"C0C0BFA4F9909099",
-21993 => x"C0C0BFA4F99090B0",
-21992 => x"C0C0BFA4F99090A4",
-21991 => x"C0C0BFA4F99090F9",
-21990 => x"C0C0BFA4F99090C0",
-21989 => x"C0C0BFA4F9908090",
-21988 => x"C0C0BFA4F9908080",
-21987 => x"C0C0BFA4F99080F8",
-21986 => x"C0C0BFA4F9908082",
-21985 => x"C0C0BFA4F9908092",
-21984 => x"C0C0BFA4F9908099",
-21983 => x"C0C0BFA4F99080B0",
-21982 => x"C0C0BFA4F99080A4",
-21981 => x"C0C0BFA4F99080F9",
-21980 => x"C0C0BFA4F99080C0",
-21979 => x"C0C0BFA4F990F890",
-21978 => x"C0C0BFA4F990F880",
-21977 => x"C0C0BFA4F990F8F8",
-21976 => x"C0C0BFA4F990F882",
-21975 => x"C0C0BFA4F990F892",
-21974 => x"C0C0BFA4F990F899",
-21973 => x"C0C0BFA4F990F8B0",
-21972 => x"C0C0BFA4F990F8A4",
-21971 => x"C0C0BFA4F990F8F9",
-21970 => x"C0C0BFA4F990F8C0",
-21969 => x"C0C0BFA4F9908290",
-21968 => x"C0C0BFA4F9908280",
-21967 => x"C0C0BFA4F99082F8",
-21966 => x"C0C0BFA4F9908282",
-21965 => x"C0C0BFA4F9908292",
-21964 => x"C0C0BFA4F9908299",
-21963 => x"C0C0BFA4F99082B0",
-21962 => x"C0C0BFA4F99082A4",
-21961 => x"C0C0BFA4F99082F9",
-21960 => x"C0C0BFA4F99082C0",
-21959 => x"C0C0BFA4F9909290",
-21958 => x"C0C0BFA4F9909280",
-21957 => x"C0C0BFA4F99092F8",
-21956 => x"C0C0BFA4F9909282",
-21955 => x"C0C0BFA4F9909292",
-21954 => x"C0C0BFA4F9909299",
-21953 => x"C0C0BFA4F99092B0",
-21952 => x"C0C0BFA4F99092A4",
-21951 => x"C0C0BFA4F99092F9",
-21950 => x"C0C0BFA4F99092C0",
-21949 => x"C0C0BFA4F9909990",
-21948 => x"C0C0BFA4F9909980",
-21947 => x"C0C0BFA4F99099F8",
-21946 => x"C0C0BFA4F9909982",
-21945 => x"C0C0BFA4F9909992",
-21944 => x"C0C0BFA4F9909999",
-21943 => x"C0C0BFA4F99099B0",
-21942 => x"C0C0BFA4F99099A4",
-21941 => x"C0C0BFA4F99099F9",
-21940 => x"C0C0BFA4F99099C0",
-21939 => x"C0C0BFA4F990B090",
-21938 => x"C0C0BFA4F990B080",
-21937 => x"C0C0BFA4F990B0F8",
-21936 => x"C0C0BFA4F990B082",
-21935 => x"C0C0BFA4F990B092",
-21934 => x"C0C0BFA4F990B099",
-21933 => x"C0C0BFA4F990B0B0",
-21932 => x"C0C0BFA4F990B0A4",
-21931 => x"C0C0BFA4F990B0F9",
-21930 => x"C0C0BFA4F990B0C0",
-21929 => x"C0C0BFA4F990A490",
-21928 => x"C0C0BFA4F990A480",
-21927 => x"C0C0BFA4F990A4F8",
-21926 => x"C0C0BFA4F990A482",
-21925 => x"C0C0BFA4F990A492",
-21924 => x"C0C0BFA4F990A499",
-21923 => x"C0C0BFA4F990A4B0",
-21922 => x"C0C0BFA4F990A4A4",
-21921 => x"C0C0BFA4F990A4F9",
-21920 => x"C0C0BFA4F990A4C0",
-21919 => x"C0C0BFA4F990F990",
-21918 => x"C0C0BFA4F990F980",
-21917 => x"C0C0BFA4F990F9F8",
-21916 => x"C0C0BFA4F990F982",
-21915 => x"C0C0BFA4F990F992",
-21914 => x"C0C0BFA4F990F999",
-21913 => x"C0C0BFA4F990F9B0",
-21912 => x"C0C0BFA4F990F9A4",
-21911 => x"C0C0BFA4F990F9F9",
-21910 => x"C0C0BFA4F990F9C0",
-21909 => x"C0C0BFA4F990C090",
-21908 => x"C0C0BFA4F990C080",
-21907 => x"C0C0BFA4F990C0F8",
-21906 => x"C0C0BFA4F990C082",
-21905 => x"C0C0BFA4F990C092",
-21904 => x"C0C0BFA4F990C099",
-21903 => x"C0C0BFA4F990C0B0",
-21902 => x"C0C0BFA4F990C0A4",
-21901 => x"C0C0BFA4F990C0F9",
-21900 => x"C0C0BFA4F990C0C0",
-21899 => x"C0C0BFA4F9809090",
-21898 => x"C0C0BFA4F9809080",
-21897 => x"C0C0BFA4F98090F8",
-21896 => x"C0C0BFA4F9809082",
-21895 => x"C0C0BFA4F9809092",
-21894 => x"C0C0BFA4F9809099",
-21893 => x"C0C0BFA4F98090B0",
-21892 => x"C0C0BFA4F98090A4",
-21891 => x"C0C0BFA4F98090F9",
-21890 => x"C0C0BFA4F98090C0",
-21889 => x"C0C0BFA4F9808090",
-21888 => x"C0C0BFA4F9808080",
-21887 => x"C0C0BFA4F98080F8",
-21886 => x"C0C0BFA4F9808082",
-21885 => x"C0C0BFA4F9808092",
-21884 => x"C0C0BFA4F9808099",
-21883 => x"C0C0BFA4F98080B0",
-21882 => x"C0C0BFA4F98080A4",
-21881 => x"C0C0BFA4F98080F9",
-21880 => x"C0C0BFA4F98080C0",
-21879 => x"C0C0BFA4F980F890",
-21878 => x"C0C0BFA4F980F880",
-21877 => x"C0C0BFA4F980F8F8",
-21876 => x"C0C0BFA4F980F882",
-21875 => x"C0C0BFA4F980F892",
-21874 => x"C0C0BFA4F980F899",
-21873 => x"C0C0BFA4F980F8B0",
-21872 => x"C0C0BFA4F980F8A4",
-21871 => x"C0C0BFA4F980F8F9",
-21870 => x"C0C0BFA4F980F8C0",
-21869 => x"C0C0BFA4F9808290",
-21868 => x"C0C0BFA4F9808280",
-21867 => x"C0C0BFA4F98082F8",
-21866 => x"C0C0BFA4F9808282",
-21865 => x"C0C0BFA4F9808292",
-21864 => x"C0C0BFA4F9808299",
-21863 => x"C0C0BFA4F98082B0",
-21862 => x"C0C0BFA4F98082A4",
-21861 => x"C0C0BFA4F98082F9",
-21860 => x"C0C0BFA4F98082C0",
-21859 => x"C0C0BFA4F9809290",
-21858 => x"C0C0BFA4F9809280",
-21857 => x"C0C0BFA4F98092F8",
-21856 => x"C0C0BFA4F9809282",
-21855 => x"C0C0BFA4F9809292",
-21854 => x"C0C0BFA4F9809299",
-21853 => x"C0C0BFA4F98092B0",
-21852 => x"C0C0BFA4F98092A4",
-21851 => x"C0C0BFA4F98092F9",
-21850 => x"C0C0BFA4F98092C0",
-21849 => x"C0C0BFA4F9809990",
-21848 => x"C0C0BFA4F9809980",
-21847 => x"C0C0BFA4F98099F8",
-21846 => x"C0C0BFA4F9809982",
-21845 => x"C0C0BFA4F9809992",
-21844 => x"C0C0BFA4F9809999",
-21843 => x"C0C0BFA4F98099B0",
-21842 => x"C0C0BFA4F98099A4",
-21841 => x"C0C0BFA4F98099F9",
-21840 => x"C0C0BFA4F98099C0",
-21839 => x"C0C0BFA4F980B090",
-21838 => x"C0C0BFA4F980B080",
-21837 => x"C0C0BFA4F980B0F8",
-21836 => x"C0C0BFA4F980B082",
-21835 => x"C0C0BFA4F980B092",
-21834 => x"C0C0BFA4F980B099",
-21833 => x"C0C0BFA4F980B0B0",
-21832 => x"C0C0BFA4F980B0A4",
-21831 => x"C0C0BFA4F980B0F9",
-21830 => x"C0C0BFA4F980B0C0",
-21829 => x"C0C0BFA4F980A490",
-21828 => x"C0C0BFA4F980A480",
-21827 => x"C0C0BFA4F980A4F8",
-21826 => x"C0C0BFA4F980A482",
-21825 => x"C0C0BFA4F980A492",
-21824 => x"C0C0BFA4F980A499",
-21823 => x"C0C0BFA4F980A4B0",
-21822 => x"C0C0BFA4F980A4A4",
-21821 => x"C0C0BFA4F980A4F9",
-21820 => x"C0C0BFA4F980A4C0",
-21819 => x"C0C0BFA4F980F990",
-21818 => x"C0C0BFA4F980F980",
-21817 => x"C0C0BFA4F980F9F8",
-21816 => x"C0C0BFA4F980F982",
-21815 => x"C0C0BFA4F980F992",
-21814 => x"C0C0BFA4F980F999",
-21813 => x"C0C0BFA4F980F9B0",
-21812 => x"C0C0BFA4F980F9A4",
-21811 => x"C0C0BFA4F980F9F9",
-21810 => x"C0C0BFA4F980F9C0",
-21809 => x"C0C0BFA4F980C090",
-21808 => x"C0C0BFA4F980C080",
-21807 => x"C0C0BFA4F980C0F8",
-21806 => x"C0C0BFA4F980C082",
-21805 => x"C0C0BFA4F980C092",
-21804 => x"C0C0BFA4F980C099",
-21803 => x"C0C0BFA4F980C0B0",
-21802 => x"C0C0BFA4F980C0A4",
-21801 => x"C0C0BFA4F980C0F9",
-21800 => x"C0C0BFA4F980C0C0",
-21799 => x"C0C0BFA4F9F89090",
-21798 => x"C0C0BFA4F9F89080",
-21797 => x"C0C0BFA4F9F890F8",
-21796 => x"C0C0BFA4F9F89082",
-21795 => x"C0C0BFA4F9F89092",
-21794 => x"C0C0BFA4F9F89099",
-21793 => x"C0C0BFA4F9F890B0",
-21792 => x"C0C0BFA4F9F890A4",
-21791 => x"C0C0BFA4F9F890F9",
-21790 => x"C0C0BFA4F9F890C0",
-21789 => x"C0C0BFA4F9F88090",
-21788 => x"C0C0BFA4F9F88080",
-21787 => x"C0C0BFA4F9F880F8",
-21786 => x"C0C0BFA4F9F88082",
-21785 => x"C0C0BFA4F9F88092",
-21784 => x"C0C0BFA4F9F88099",
-21783 => x"C0C0BFA4F9F880B0",
-21782 => x"C0C0BFA4F9F880A4",
-21781 => x"C0C0BFA4F9F880F9",
-21780 => x"C0C0BFA4F9F880C0",
-21779 => x"C0C0BFA4F9F8F890",
-21778 => x"C0C0BFA4F9F8F880",
-21777 => x"C0C0BFA4F9F8F8F8",
-21776 => x"C0C0BFA4F9F8F882",
-21775 => x"C0C0BFA4F9F8F892",
-21774 => x"C0C0BFA4F9F8F899",
-21773 => x"C0C0BFA4F9F8F8B0",
-21772 => x"C0C0BFA4F9F8F8A4",
-21771 => x"C0C0BFA4F9F8F8F9",
-21770 => x"C0C0BFA4F9F8F8C0",
-21769 => x"C0C0BFA4F9F88290",
-21768 => x"C0C0BFA4F9F88280",
-21767 => x"C0C0BFA4F9F882F8",
-21766 => x"C0C0BFA4F9F88282",
-21765 => x"C0C0BFA4F9F88292",
-21764 => x"C0C0BFA4F9F88299",
-21763 => x"C0C0BFA4F9F882B0",
-21762 => x"C0C0BFA4F9F882A4",
-21761 => x"C0C0BFA4F9F882F9",
-21760 => x"C0C0BFA4F9F882C0",
-21759 => x"C0C0BFA4F9F89290",
-21758 => x"C0C0BFA4F9F89280",
-21757 => x"C0C0BFA4F9F892F8",
-21756 => x"C0C0BFA4F9F89282",
-21755 => x"C0C0BFA4F9F89292",
-21754 => x"C0C0BFA4F9F89299",
-21753 => x"C0C0BFA4F9F892B0",
-21752 => x"C0C0BFA4F9F892A4",
-21751 => x"C0C0BFA4F9F892F9",
-21750 => x"C0C0BFA4F9F892C0",
-21749 => x"C0C0BFA4F9F89990",
-21748 => x"C0C0BFA4F9F89980",
-21747 => x"C0C0BFA4F9F899F8",
-21746 => x"C0C0BFA4F9F89982",
-21745 => x"C0C0BFA4F9F89992",
-21744 => x"C0C0BFA4F9F89999",
-21743 => x"C0C0BFA4F9F899B0",
-21742 => x"C0C0BFA4F9F899A4",
-21741 => x"C0C0BFA4F9F899F9",
-21740 => x"C0C0BFA4F9F899C0",
-21739 => x"C0C0BFA4F9F8B090",
-21738 => x"C0C0BFA4F9F8B080",
-21737 => x"C0C0BFA4F9F8B0F8",
-21736 => x"C0C0BFA4F9F8B082",
-21735 => x"C0C0BFA4F9F8B092",
-21734 => x"C0C0BFA4F9F8B099",
-21733 => x"C0C0BFA4F9F8B0B0",
-21732 => x"C0C0BFA4F9F8B0A4",
-21731 => x"C0C0BFA4F9F8B0F9",
-21730 => x"C0C0BFA4F9F8B0C0",
-21729 => x"C0C0BFA4F9F8A490",
-21728 => x"C0C0BFA4F9F8A480",
-21727 => x"C0C0BFA4F9F8A4F8",
-21726 => x"C0C0BFA4F9F8A482",
-21725 => x"C0C0BFA4F9F8A492",
-21724 => x"C0C0BFA4F9F8A499",
-21723 => x"C0C0BFA4F9F8A4B0",
-21722 => x"C0C0BFA4F9F8A4A4",
-21721 => x"C0C0BFA4F9F8A4F9",
-21720 => x"C0C0BFA4F9F8A4C0",
-21719 => x"C0C0BFA4F9F8F990",
-21718 => x"C0C0BFA4F9F8F980",
-21717 => x"C0C0BFA4F9F8F9F8",
-21716 => x"C0C0BFA4F9F8F982",
-21715 => x"C0C0BFA4F9F8F992",
-21714 => x"C0C0BFA4F9F8F999",
-21713 => x"C0C0BFA4F9F8F9B0",
-21712 => x"C0C0BFA4F9F8F9A4",
-21711 => x"C0C0BFA4F9F8F9F9",
-21710 => x"C0C0BFA4F9F8F9C0",
-21709 => x"C0C0BFA4F9F8C090",
-21708 => x"C0C0BFA4F9F8C080",
-21707 => x"C0C0BFA4F9F8C0F8",
-21706 => x"C0C0BFA4F9F8C082",
-21705 => x"C0C0BFA4F9F8C092",
-21704 => x"C0C0BFA4F9F8C099",
-21703 => x"C0C0BFA4F9F8C0B0",
-21702 => x"C0C0BFA4F9F8C0A4",
-21701 => x"C0C0BFA4F9F8C0F9",
-21700 => x"C0C0BFA4F9F8C0C0",
-21699 => x"C0C0BFA4F9829090",
-21698 => x"C0C0BFA4F9829080",
-21697 => x"C0C0BFA4F98290F8",
-21696 => x"C0C0BFA4F9829082",
-21695 => x"C0C0BFA4F9829092",
-21694 => x"C0C0BFA4F9829099",
-21693 => x"C0C0BFA4F98290B0",
-21692 => x"C0C0BFA4F98290A4",
-21691 => x"C0C0BFA4F98290F9",
-21690 => x"C0C0BFA4F98290C0",
-21689 => x"C0C0BFA4F9828090",
-21688 => x"C0C0BFA4F9828080",
-21687 => x"C0C0BFA4F98280F8",
-21686 => x"C0C0BFA4F9828082",
-21685 => x"C0C0BFA4F9828092",
-21684 => x"C0C0BFA4F9828099",
-21683 => x"C0C0BFA4F98280B0",
-21682 => x"C0C0BFA4F98280A4",
-21681 => x"C0C0BFA4F98280F9",
-21680 => x"C0C0BFA4F98280C0",
-21679 => x"C0C0BFA4F982F890",
-21678 => x"C0C0BFA4F982F880",
-21677 => x"C0C0BFA4F982F8F8",
-21676 => x"C0C0BFA4F982F882",
-21675 => x"C0C0BFA4F982F892",
-21674 => x"C0C0BFA4F982F899",
-21673 => x"C0C0BFA4F982F8B0",
-21672 => x"C0C0BFA4F982F8A4",
-21671 => x"C0C0BFA4F982F8F9",
-21670 => x"C0C0BFA4F982F8C0",
-21669 => x"C0C0BFA4F9828290",
-21668 => x"C0C0BFA4F9828280",
-21667 => x"C0C0BFA4F98282F8",
-21666 => x"C0C0BFA4F9828282",
-21665 => x"C0C0BFA4F9828292",
-21664 => x"C0C0BFA4F9828299",
-21663 => x"C0C0BFA4F98282B0",
-21662 => x"C0C0BFA4F98282A4",
-21661 => x"C0C0BFA4F98282F9",
-21660 => x"C0C0BFA4F98282C0",
-21659 => x"C0C0BFA4F9829290",
-21658 => x"C0C0BFA4F9829280",
-21657 => x"C0C0BFA4F98292F8",
-21656 => x"C0C0BFA4F9829282",
-21655 => x"C0C0BFA4F9829292",
-21654 => x"C0C0BFA4F9829299",
-21653 => x"C0C0BFA4F98292B0",
-21652 => x"C0C0BFA4F98292A4",
-21651 => x"C0C0BFA4F98292F9",
-21650 => x"C0C0BFA4F98292C0",
-21649 => x"C0C0BFA4F9829990",
-21648 => x"C0C0BFA4F9829980",
-21647 => x"C0C0BFA4F98299F8",
-21646 => x"C0C0BFA4F9829982",
-21645 => x"C0C0BFA4F9829992",
-21644 => x"C0C0BFA4F9829999",
-21643 => x"C0C0BFA4F98299B0",
-21642 => x"C0C0BFA4F98299A4",
-21641 => x"C0C0BFA4F98299F9",
-21640 => x"C0C0BFA4F98299C0",
-21639 => x"C0C0BFA4F982B090",
-21638 => x"C0C0BFA4F982B080",
-21637 => x"C0C0BFA4F982B0F8",
-21636 => x"C0C0BFA4F982B082",
-21635 => x"C0C0BFA4F982B092",
-21634 => x"C0C0BFA4F982B099",
-21633 => x"C0C0BFA4F982B0B0",
-21632 => x"C0C0BFA4F982B0A4",
-21631 => x"C0C0BFA4F982B0F9",
-21630 => x"C0C0BFA4F982B0C0",
-21629 => x"C0C0BFA4F982A490",
-21628 => x"C0C0BFA4F982A480",
-21627 => x"C0C0BFA4F982A4F8",
-21626 => x"C0C0BFA4F982A482",
-21625 => x"C0C0BFA4F982A492",
-21624 => x"C0C0BFA4F982A499",
-21623 => x"C0C0BFA4F982A4B0",
-21622 => x"C0C0BFA4F982A4A4",
-21621 => x"C0C0BFA4F982A4F9",
-21620 => x"C0C0BFA4F982A4C0",
-21619 => x"C0C0BFA4F982F990",
-21618 => x"C0C0BFA4F982F980",
-21617 => x"C0C0BFA4F982F9F8",
-21616 => x"C0C0BFA4F982F982",
-21615 => x"C0C0BFA4F982F992",
-21614 => x"C0C0BFA4F982F999",
-21613 => x"C0C0BFA4F982F9B0",
-21612 => x"C0C0BFA4F982F9A4",
-21611 => x"C0C0BFA4F982F9F9",
-21610 => x"C0C0BFA4F982F9C0",
-21609 => x"C0C0BFA4F982C090",
-21608 => x"C0C0BFA4F982C080",
-21607 => x"C0C0BFA4F982C0F8",
-21606 => x"C0C0BFA4F982C082",
-21605 => x"C0C0BFA4F982C092",
-21604 => x"C0C0BFA4F982C099",
-21603 => x"C0C0BFA4F982C0B0",
-21602 => x"C0C0BFA4F982C0A4",
-21601 => x"C0C0BFA4F982C0F9",
-21600 => x"C0C0BFA4F982C0C0",
-21599 => x"C0C0BFA4F9929090",
-21598 => x"C0C0BFA4F9929080",
-21597 => x"C0C0BFA4F99290F8",
-21596 => x"C0C0BFA4F9929082",
-21595 => x"C0C0BFA4F9929092",
-21594 => x"C0C0BFA4F9929099",
-21593 => x"C0C0BFA4F99290B0",
-21592 => x"C0C0BFA4F99290A4",
-21591 => x"C0C0BFA4F99290F9",
-21590 => x"C0C0BFA4F99290C0",
-21589 => x"C0C0BFA4F9928090",
-21588 => x"C0C0BFA4F9928080",
-21587 => x"C0C0BFA4F99280F8",
-21586 => x"C0C0BFA4F9928082",
-21585 => x"C0C0BFA4F9928092",
-21584 => x"C0C0BFA4F9928099",
-21583 => x"C0C0BFA4F99280B0",
-21582 => x"C0C0BFA4F99280A4",
-21581 => x"C0C0BFA4F99280F9",
-21580 => x"C0C0BFA4F99280C0",
-21579 => x"C0C0BFA4F992F890",
-21578 => x"C0C0BFA4F992F880",
-21577 => x"C0C0BFA4F992F8F8",
-21576 => x"C0C0BFA4F992F882",
-21575 => x"C0C0BFA4F992F892",
-21574 => x"C0C0BFA4F992F899",
-21573 => x"C0C0BFA4F992F8B0",
-21572 => x"C0C0BFA4F992F8A4",
-21571 => x"C0C0BFA4F992F8F9",
-21570 => x"C0C0BFA4F992F8C0",
-21569 => x"C0C0BFA4F9928290",
-21568 => x"C0C0BFA4F9928280",
-21567 => x"C0C0BFA4F99282F8",
-21566 => x"C0C0BFA4F9928282",
-21565 => x"C0C0BFA4F9928292",
-21564 => x"C0C0BFA4F9928299",
-21563 => x"C0C0BFA4F99282B0",
-21562 => x"C0C0BFA4F99282A4",
-21561 => x"C0C0BFA4F99282F9",
-21560 => x"C0C0BFA4F99282C0",
-21559 => x"C0C0BFA4F9929290",
-21558 => x"C0C0BFA4F9929280",
-21557 => x"C0C0BFA4F99292F8",
-21556 => x"C0C0BFA4F9929282",
-21555 => x"C0C0BFA4F9929292",
-21554 => x"C0C0BFA4F9929299",
-21553 => x"C0C0BFA4F99292B0",
-21552 => x"C0C0BFA4F99292A4",
-21551 => x"C0C0BFA4F99292F9",
-21550 => x"C0C0BFA4F99292C0",
-21549 => x"C0C0BFA4F9929990",
-21548 => x"C0C0BFA4F9929980",
-21547 => x"C0C0BFA4F99299F8",
-21546 => x"C0C0BFA4F9929982",
-21545 => x"C0C0BFA4F9929992",
-21544 => x"C0C0BFA4F9929999",
-21543 => x"C0C0BFA4F99299B0",
-21542 => x"C0C0BFA4F99299A4",
-21541 => x"C0C0BFA4F99299F9",
-21540 => x"C0C0BFA4F99299C0",
-21539 => x"C0C0BFA4F992B090",
-21538 => x"C0C0BFA4F992B080",
-21537 => x"C0C0BFA4F992B0F8",
-21536 => x"C0C0BFA4F992B082",
-21535 => x"C0C0BFA4F992B092",
-21534 => x"C0C0BFA4F992B099",
-21533 => x"C0C0BFA4F992B0B0",
-21532 => x"C0C0BFA4F992B0A4",
-21531 => x"C0C0BFA4F992B0F9",
-21530 => x"C0C0BFA4F992B0C0",
-21529 => x"C0C0BFA4F992A490",
-21528 => x"C0C0BFA4F992A480",
-21527 => x"C0C0BFA4F992A4F8",
-21526 => x"C0C0BFA4F992A482",
-21525 => x"C0C0BFA4F992A492",
-21524 => x"C0C0BFA4F992A499",
-21523 => x"C0C0BFA4F992A4B0",
-21522 => x"C0C0BFA4F992A4A4",
-21521 => x"C0C0BFA4F992A4F9",
-21520 => x"C0C0BFA4F992A4C0",
-21519 => x"C0C0BFA4F992F990",
-21518 => x"C0C0BFA4F992F980",
-21517 => x"C0C0BFA4F992F9F8",
-21516 => x"C0C0BFA4F992F982",
-21515 => x"C0C0BFA4F992F992",
-21514 => x"C0C0BFA4F992F999",
-21513 => x"C0C0BFA4F992F9B0",
-21512 => x"C0C0BFA4F992F9A4",
-21511 => x"C0C0BFA4F992F9F9",
-21510 => x"C0C0BFA4F992F9C0",
-21509 => x"C0C0BFA4F992C090",
-21508 => x"C0C0BFA4F992C080",
-21507 => x"C0C0BFA4F992C0F8",
-21506 => x"C0C0BFA4F992C082",
-21505 => x"C0C0BFA4F992C092",
-21504 => x"C0C0BFA4F992C099",
-21503 => x"C0C0BFA4F992C0B0",
-21502 => x"C0C0BFA4F992C0A4",
-21501 => x"C0C0BFA4F992C0F9",
-21500 => x"C0C0BFA4F992C0C0",
-21499 => x"C0C0BFA4F9999090",
-21498 => x"C0C0BFA4F9999080",
-21497 => x"C0C0BFA4F99990F8",
-21496 => x"C0C0BFA4F9999082",
-21495 => x"C0C0BFA4F9999092",
-21494 => x"C0C0BFA4F9999099",
-21493 => x"C0C0BFA4F99990B0",
-21492 => x"C0C0BFA4F99990A4",
-21491 => x"C0C0BFA4F99990F9",
-21490 => x"C0C0BFA4F99990C0",
-21489 => x"C0C0BFA4F9998090",
-21488 => x"C0C0BFA4F9998080",
-21487 => x"C0C0BFA4F99980F8",
-21486 => x"C0C0BFA4F9998082",
-21485 => x"C0C0BFA4F9998092",
-21484 => x"C0C0BFA4F9998099",
-21483 => x"C0C0BFA4F99980B0",
-21482 => x"C0C0BFA4F99980A4",
-21481 => x"C0C0BFA4F99980F9",
-21480 => x"C0C0BFA4F99980C0",
-21479 => x"C0C0BFA4F999F890",
-21478 => x"C0C0BFA4F999F880",
-21477 => x"C0C0BFA4F999F8F8",
-21476 => x"C0C0BFA4F999F882",
-21475 => x"C0C0BFA4F999F892",
-21474 => x"C0C0BFA4F999F899",
-21473 => x"C0C0BFA4F999F8B0",
-21472 => x"C0C0BFA4F999F8A4",
-21471 => x"C0C0BFA4F999F8F9",
-21470 => x"C0C0BFA4F999F8C0",
-21469 => x"C0C0BFA4F9998290",
-21468 => x"C0C0BFA4F9998280",
-21467 => x"C0C0BFA4F99982F8",
-21466 => x"C0C0BFA4F9998282",
-21465 => x"C0C0BFA4F9998292",
-21464 => x"C0C0BFA4F9998299",
-21463 => x"C0C0BFA4F99982B0",
-21462 => x"C0C0BFA4F99982A4",
-21461 => x"C0C0BFA4F99982F9",
-21460 => x"C0C0BFA4F99982C0",
-21459 => x"C0C0BFA4F9999290",
-21458 => x"C0C0BFA4F9999280",
-21457 => x"C0C0BFA4F99992F8",
-21456 => x"C0C0BFA4F9999282",
-21455 => x"C0C0BFA4F9999292",
-21454 => x"C0C0BFA4F9999299",
-21453 => x"C0C0BFA4F99992B0",
-21452 => x"C0C0BFA4F99992A4",
-21451 => x"C0C0BFA4F99992F9",
-21450 => x"C0C0BFA4F99992C0",
-21449 => x"C0C0BFA4F9999990",
-21448 => x"C0C0BFA4F9999980",
-21447 => x"C0C0BFA4F99999F8",
-21446 => x"C0C0BFA4F9999982",
-21445 => x"C0C0BFA4F9999992",
-21444 => x"C0C0BFA4F9999999",
-21443 => x"C0C0BFA4F99999B0",
-21442 => x"C0C0BFA4F99999A4",
-21441 => x"C0C0BFA4F99999F9",
-21440 => x"C0C0BFA4F99999C0",
-21439 => x"C0C0BFA4F999B090",
-21438 => x"C0C0BFA4F999B080",
-21437 => x"C0C0BFA4F999B0F8",
-21436 => x"C0C0BFA4F999B082",
-21435 => x"C0C0BFA4F999B092",
-21434 => x"C0C0BFA4F999B099",
-21433 => x"C0C0BFA4F999B0B0",
-21432 => x"C0C0BFA4F999B0A4",
-21431 => x"C0C0BFA4F999B0F9",
-21430 => x"C0C0BFA4F999B0C0",
-21429 => x"C0C0BFA4F999A490",
-21428 => x"C0C0BFA4F999A480",
-21427 => x"C0C0BFA4F999A4F8",
-21426 => x"C0C0BFA4F999A482",
-21425 => x"C0C0BFA4F999A492",
-21424 => x"C0C0BFA4F999A499",
-21423 => x"C0C0BFA4F999A4B0",
-21422 => x"C0C0BFA4F999A4A4",
-21421 => x"C0C0BFA4F999A4F9",
-21420 => x"C0C0BFA4F999A4C0",
-21419 => x"C0C0BFA4F999F990",
-21418 => x"C0C0BFA4F999F980",
-21417 => x"C0C0BFA4F999F9F8",
-21416 => x"C0C0BFA4F999F982",
-21415 => x"C0C0BFA4F999F992",
-21414 => x"C0C0BFA4F999F999",
-21413 => x"C0C0BFA4F999F9B0",
-21412 => x"C0C0BFA4F999F9A4",
-21411 => x"C0C0BFA4F999F9F9",
-21410 => x"C0C0BFA4F999F9C0",
-21409 => x"C0C0BFA4F999C090",
-21408 => x"C0C0BFA4F999C080",
-21407 => x"C0C0BFA4F999C0F8",
-21406 => x"C0C0BFA4F999C082",
-21405 => x"C0C0BFA4F999C092",
-21404 => x"C0C0BFA4F999C099",
-21403 => x"C0C0BFA4F999C0B0",
-21402 => x"C0C0BFA4F999C0A4",
-21401 => x"C0C0BFA4F999C0F9",
-21400 => x"C0C0BFA4F999C0C0",
-21399 => x"C0C0BFA4F9B09090",
-21398 => x"C0C0BFA4F9B09080",
-21397 => x"C0C0BFA4F9B090F8",
-21396 => x"C0C0BFA4F9B09082",
-21395 => x"C0C0BFA4F9B09092",
-21394 => x"C0C0BFA4F9B09099",
-21393 => x"C0C0BFA4F9B090B0",
-21392 => x"C0C0BFA4F9B090A4",
-21391 => x"C0C0BFA4F9B090F9",
-21390 => x"C0C0BFA4F9B090C0",
-21389 => x"C0C0BFA4F9B08090",
-21388 => x"C0C0BFA4F9B08080",
-21387 => x"C0C0BFA4F9B080F8",
-21386 => x"C0C0BFA4F9B08082",
-21385 => x"C0C0BFA4F9B08092",
-21384 => x"C0C0BFA4F9B08099",
-21383 => x"C0C0BFA4F9B080B0",
-21382 => x"C0C0BFA4F9B080A4",
-21381 => x"C0C0BFA4F9B080F9",
-21380 => x"C0C0BFA4F9B080C0",
-21379 => x"C0C0BFA4F9B0F890",
-21378 => x"C0C0BFA4F9B0F880",
-21377 => x"C0C0BFA4F9B0F8F8",
-21376 => x"C0C0BFA4F9B0F882",
-21375 => x"C0C0BFA4F9B0F892",
-21374 => x"C0C0BFA4F9B0F899",
-21373 => x"C0C0BFA4F9B0F8B0",
-21372 => x"C0C0BFA4F9B0F8A4",
-21371 => x"C0C0BFA4F9B0F8F9",
-21370 => x"C0C0BFA4F9B0F8C0",
-21369 => x"C0C0BFA4F9B08290",
-21368 => x"C0C0BFA4F9B08280",
-21367 => x"C0C0BFA4F9B082F8",
-21366 => x"C0C0BFA4F9B08282",
-21365 => x"C0C0BFA4F9B08292",
-21364 => x"C0C0BFA4F9B08299",
-21363 => x"C0C0BFA4F9B082B0",
-21362 => x"C0C0BFA4F9B082A4",
-21361 => x"C0C0BFA4F9B082F9",
-21360 => x"C0C0BFA4F9B082C0",
-21359 => x"C0C0BFA4F9B09290",
-21358 => x"C0C0BFA4F9B09280",
-21357 => x"C0C0BFA4F9B092F8",
-21356 => x"C0C0BFA4F9B09282",
-21355 => x"C0C0BFA4F9B09292",
-21354 => x"C0C0BFA4F9B09299",
-21353 => x"C0C0BFA4F9B092B0",
-21352 => x"C0C0BFA4F9B092A4",
-21351 => x"C0C0BFA4F9B092F9",
-21350 => x"C0C0BFA4F9B092C0",
-21349 => x"C0C0BFA4F9B09990",
-21348 => x"C0C0BFA4F9B09980",
-21347 => x"C0C0BFA4F9B099F8",
-21346 => x"C0C0BFA4F9B09982",
-21345 => x"C0C0BFA4F9B09992",
-21344 => x"C0C0BFA4F9B09999",
-21343 => x"C0C0BFA4F9B099B0",
-21342 => x"C0C0BFA4F9B099A4",
-21341 => x"C0C0BFA4F9B099F9",
-21340 => x"C0C0BFA4F9B099C0",
-21339 => x"C0C0BFA4F9B0B090",
-21338 => x"C0C0BFA4F9B0B080",
-21337 => x"C0C0BFA4F9B0B0F8",
-21336 => x"C0C0BFA4F9B0B082",
-21335 => x"C0C0BFA4F9B0B092",
-21334 => x"C0C0BFA4F9B0B099",
-21333 => x"C0C0BFA4F9B0B0B0",
-21332 => x"C0C0BFA4F9B0B0A4",
-21331 => x"C0C0BFA4F9B0B0F9",
-21330 => x"C0C0BFA4F9B0B0C0",
-21329 => x"C0C0BFA4F9B0A490",
-21328 => x"C0C0BFA4F9B0A480",
-21327 => x"C0C0BFA4F9B0A4F8",
-21326 => x"C0C0BFA4F9B0A482",
-21325 => x"C0C0BFA4F9B0A492",
-21324 => x"C0C0BFA4F9B0A499",
-21323 => x"C0C0BFA4F9B0A4B0",
-21322 => x"C0C0BFA4F9B0A4A4",
-21321 => x"C0C0BFA4F9B0A4F9",
-21320 => x"C0C0BFA4F9B0A4C0",
-21319 => x"C0C0BFA4F9B0F990",
-21318 => x"C0C0BFA4F9B0F980",
-21317 => x"C0C0BFA4F9B0F9F8",
-21316 => x"C0C0BFA4F9B0F982",
-21315 => x"C0C0BFA4F9B0F992",
-21314 => x"C0C0BFA4F9B0F999",
-21313 => x"C0C0BFA4F9B0F9B0",
-21312 => x"C0C0BFA4F9B0F9A4",
-21311 => x"C0C0BFA4F9B0F9F9",
-21310 => x"C0C0BFA4F9B0F9C0",
-21309 => x"C0C0BFA4F9B0C090",
-21308 => x"C0C0BFA4F9B0C080",
-21307 => x"C0C0BFA4F9B0C0F8",
-21306 => x"C0C0BFA4F9B0C082",
-21305 => x"C0C0BFA4F9B0C092",
-21304 => x"C0C0BFA4F9B0C099",
-21303 => x"C0C0BFA4F9B0C0B0",
-21302 => x"C0C0BFA4F9B0C0A4",
-21301 => x"C0C0BFA4F9B0C0F9",
-21300 => x"C0C0BFA4F9B0C0C0",
-21299 => x"C0C0BFA4F9A49090",
-21298 => x"C0C0BFA4F9A49080",
-21297 => x"C0C0BFA4F9A490F8",
-21296 => x"C0C0BFA4F9A49082",
-21295 => x"C0C0BFA4F9A49092",
-21294 => x"C0C0BFA4F9A49099",
-21293 => x"C0C0BFA4F9A490B0",
-21292 => x"C0C0BFA4F9A490A4",
-21291 => x"C0C0BFA4F9A490F9",
-21290 => x"C0C0BFA4F9A490C0",
-21289 => x"C0C0BFA4F9A48090",
-21288 => x"C0C0BFA4F9A48080",
-21287 => x"C0C0BFA4F9A480F8",
-21286 => x"C0C0BFA4F9A48082",
-21285 => x"C0C0BFA4F9A48092",
-21284 => x"C0C0BFA4F9A48099",
-21283 => x"C0C0BFA4F9A480B0",
-21282 => x"C0C0BFA4F9A480A4",
-21281 => x"C0C0BFA4F9A480F9",
-21280 => x"C0C0BFA4F9A480C0",
-21279 => x"C0C0BFA4F9A4F890",
-21278 => x"C0C0BFA4F9A4F880",
-21277 => x"C0C0BFA4F9A4F8F8",
-21276 => x"C0C0BFA4F9A4F882",
-21275 => x"C0C0BFA4F9A4F892",
-21274 => x"C0C0BFA4F9A4F899",
-21273 => x"C0C0BFA4F9A4F8B0",
-21272 => x"C0C0BFA4F9A4F8A4",
-21271 => x"C0C0BFA4F9A4F8F9",
-21270 => x"C0C0BFA4F9A4F8C0",
-21269 => x"C0C0BFA4F9A48290",
-21268 => x"C0C0BFA4F9A48280",
-21267 => x"C0C0BFA4F9A482F8",
-21266 => x"C0C0BFA4F9A48282",
-21265 => x"C0C0BFA4F9A48292",
-21264 => x"C0C0BFA4F9A48299",
-21263 => x"C0C0BFA4F9A482B0",
-21262 => x"C0C0BFA4F9A482A4",
-21261 => x"C0C0BFA4F9A482F9",
-21260 => x"C0C0BFA4F9A482C0",
-21259 => x"C0C0BFA4F9A49290",
-21258 => x"C0C0BFA4F9A49280",
-21257 => x"C0C0BFA4F9A492F8",
-21256 => x"C0C0BFA4F9A49282",
-21255 => x"C0C0BFA4F9A49292",
-21254 => x"C0C0BFA4F9A49299",
-21253 => x"C0C0BFA4F9A492B0",
-21252 => x"C0C0BFA4F9A492A4",
-21251 => x"C0C0BFA4F9A492F9",
-21250 => x"C0C0BFA4F9A492C0",
-21249 => x"C0C0BFA4F9A49990",
-21248 => x"C0C0BFA4F9A49980",
-21247 => x"C0C0BFA4F9A499F8",
-21246 => x"C0C0BFA4F9A49982",
-21245 => x"C0C0BFA4F9A49992",
-21244 => x"C0C0BFA4F9A49999",
-21243 => x"C0C0BFA4F9A499B0",
-21242 => x"C0C0BFA4F9A499A4",
-21241 => x"C0C0BFA4F9A499F9",
-21240 => x"C0C0BFA4F9A499C0",
-21239 => x"C0C0BFA4F9A4B090",
-21238 => x"C0C0BFA4F9A4B080",
-21237 => x"C0C0BFA4F9A4B0F8",
-21236 => x"C0C0BFA4F9A4B082",
-21235 => x"C0C0BFA4F9A4B092",
-21234 => x"C0C0BFA4F9A4B099",
-21233 => x"C0C0BFA4F9A4B0B0",
-21232 => x"C0C0BFA4F9A4B0A4",
-21231 => x"C0C0BFA4F9A4B0F9",
-21230 => x"C0C0BFA4F9A4B0C0",
-21229 => x"C0C0BFA4F9A4A490",
-21228 => x"C0C0BFA4F9A4A480",
-21227 => x"C0C0BFA4F9A4A4F8",
-21226 => x"C0C0BFA4F9A4A482",
-21225 => x"C0C0BFA4F9A4A492",
-21224 => x"C0C0BFA4F9A4A499",
-21223 => x"C0C0BFA4F9A4A4B0",
-21222 => x"C0C0BFA4F9A4A4A4",
-21221 => x"C0C0BFA4F9A4A4F9",
-21220 => x"C0C0BFA4F9A4A4C0",
-21219 => x"C0C0BFA4F9A4F990",
-21218 => x"C0C0BFA4F9A4F980",
-21217 => x"C0C0BFA4F9A4F9F8",
-21216 => x"C0C0BFA4F9A4F982",
-21215 => x"C0C0BFA4F9A4F992",
-21214 => x"C0C0BFA4F9A4F999",
-21213 => x"C0C0BFA4F9A4F9B0",
-21212 => x"C0C0BFA4F9A4F9A4",
-21211 => x"C0C0BFA4F9A4F9F9",
-21210 => x"C0C0BFA4F9A4F9C0",
-21209 => x"C0C0BFA4F9A4C090",
-21208 => x"C0C0BFA4F9A4C080",
-21207 => x"C0C0BFA4F9A4C0F8",
-21206 => x"C0C0BFA4F9A4C082",
-21205 => x"C0C0BFA4F9A4C092",
-21204 => x"C0C0BFA4F9A4C099",
-21203 => x"C0C0BFA4F9A4C0B0",
-21202 => x"C0C0BFA4F9A4C0A4",
-21201 => x"C0C0BFA4F9A4C0F9",
-21200 => x"C0C0BFA4F9A4C0C0",
-21199 => x"C0C0BFA4F9F99090",
-21198 => x"C0C0BFA4F9F99080",
-21197 => x"C0C0BFA4F9F990F8",
-21196 => x"C0C0BFA4F9F99082",
-21195 => x"C0C0BFA4F9F99092",
-21194 => x"C0C0BFA4F9F99099",
-21193 => x"C0C0BFA4F9F990B0",
-21192 => x"C0C0BFA4F9F990A4",
-21191 => x"C0C0BFA4F9F990F9",
-21190 => x"C0C0BFA4F9F990C0",
-21189 => x"C0C0BFA4F9F98090",
-21188 => x"C0C0BFA4F9F98080",
-21187 => x"C0C0BFA4F9F980F8",
-21186 => x"C0C0BFA4F9F98082",
-21185 => x"C0C0BFA4F9F98092",
-21184 => x"C0C0BFA4F9F98099",
-21183 => x"C0C0BFA4F9F980B0",
-21182 => x"C0C0BFA4F9F980A4",
-21181 => x"C0C0BFA4F9F980F9",
-21180 => x"C0C0BFA4F9F980C0",
-21179 => x"C0C0BFA4F9F9F890",
-21178 => x"C0C0BFA4F9F9F880",
-21177 => x"C0C0BFA4F9F9F8F8",
-21176 => x"C0C0BFA4F9F9F882",
-21175 => x"C0C0BFA4F9F9F892",
-21174 => x"C0C0BFA4F9F9F899",
-21173 => x"C0C0BFA4F9F9F8B0",
-21172 => x"C0C0BFA4F9F9F8A4",
-21171 => x"C0C0BFA4F9F9F8F9",
-21170 => x"C0C0BFA4F9F9F8C0",
-21169 => x"C0C0BFA4F9F98290",
-21168 => x"C0C0BFA4F9F98280",
-21167 => x"C0C0BFA4F9F982F8",
-21166 => x"C0C0BFA4F9F98282",
-21165 => x"C0C0BFA4F9F98292",
-21164 => x"C0C0BFA4F9F98299",
-21163 => x"C0C0BFA4F9F982B0",
-21162 => x"C0C0BFA4F9F982A4",
-21161 => x"C0C0BFA4F9F982F9",
-21160 => x"C0C0BFA4F9F982C0",
-21159 => x"C0C0BFA4F9F99290",
-21158 => x"C0C0BFA4F9F99280",
-21157 => x"C0C0BFA4F9F992F8",
-21156 => x"C0C0BFA4F9F99282",
-21155 => x"C0C0BFA4F9F99292",
-21154 => x"C0C0BFA4F9F99299",
-21153 => x"C0C0BFA4F9F992B0",
-21152 => x"C0C0BFA4F9F992A4",
-21151 => x"C0C0BFA4F9F992F9",
-21150 => x"C0C0BFA4F9F992C0",
-21149 => x"C0C0BFA4F9F99990",
-21148 => x"C0C0BFA4F9F99980",
-21147 => x"C0C0BFA4F9F999F8",
-21146 => x"C0C0BFA4F9F99982",
-21145 => x"C0C0BFA4F9F99992",
-21144 => x"C0C0BFA4F9F99999",
-21143 => x"C0C0BFA4F9F999B0",
-21142 => x"C0C0BFA4F9F999A4",
-21141 => x"C0C0BFA4F9F999F9",
-21140 => x"C0C0BFA4F9F999C0",
-21139 => x"C0C0BFA4F9F9B090",
-21138 => x"C0C0BFA4F9F9B080",
-21137 => x"C0C0BFA4F9F9B0F8",
-21136 => x"C0C0BFA4F9F9B082",
-21135 => x"C0C0BFA4F9F9B092",
-21134 => x"C0C0BFA4F9F9B099",
-21133 => x"C0C0BFA4F9F9B0B0",
-21132 => x"C0C0BFA4F9F9B0A4",
-21131 => x"C0C0BFA4F9F9B0F9",
-21130 => x"C0C0BFA4F9F9B0C0",
-21129 => x"C0C0BFA4F9F9A490",
-21128 => x"C0C0BFA4F9F9A480",
-21127 => x"C0C0BFA4F9F9A4F8",
-21126 => x"C0C0BFA4F9F9A482",
-21125 => x"C0C0BFA4F9F9A492",
-21124 => x"C0C0BFA4F9F9A499",
-21123 => x"C0C0BFA4F9F9A4B0",
-21122 => x"C0C0BFA4F9F9A4A4",
-21121 => x"C0C0BFA4F9F9A4F9",
-21120 => x"C0C0BFA4F9F9A4C0",
-21119 => x"C0C0BFA4F9F9F990",
-21118 => x"C0C0BFA4F9F9F980",
-21117 => x"C0C0BFA4F9F9F9F8",
-21116 => x"C0C0BFA4F9F9F982",
-21115 => x"C0C0BFA4F9F9F992",
-21114 => x"C0C0BFA4F9F9F999",
-21113 => x"C0C0BFA4F9F9F9B0",
-21112 => x"C0C0BFA4F9F9F9A4",
-21111 => x"C0C0BFA4F9F9F9F9",
-21110 => x"C0C0BFA4F9F9F9C0",
-21109 => x"C0C0BFA4F9F9C090",
-21108 => x"C0C0BFA4F9F9C080",
-21107 => x"C0C0BFA4F9F9C0F8",
-21106 => x"C0C0BFA4F9F9C082",
-21105 => x"C0C0BFA4F9F9C092",
-21104 => x"C0C0BFA4F9F9C099",
-21103 => x"C0C0BFA4F9F9C0B0",
-21102 => x"C0C0BFA4F9F9C0A4",
-21101 => x"C0C0BFA4F9F9C0F9",
-21100 => x"C0C0BFA4F9F9C0C0",
-21099 => x"C0C0BFA4F9C09090",
-21098 => x"C0C0BFA4F9C09080",
-21097 => x"C0C0BFA4F9C090F8",
-21096 => x"C0C0BFA4F9C09082",
-21095 => x"C0C0BFA4F9C09092",
-21094 => x"C0C0BFA4F9C09099",
-21093 => x"C0C0BFA4F9C090B0",
-21092 => x"C0C0BFA4F9C090A4",
-21091 => x"C0C0BFA4F9C090F9",
-21090 => x"C0C0BFA4F9C090C0",
-21089 => x"C0C0BFA4F9C08090",
-21088 => x"C0C0BFA4F9C08080",
-21087 => x"C0C0BFA4F9C080F8",
-21086 => x"C0C0BFA4F9C08082",
-21085 => x"C0C0BFA4F9C08092",
-21084 => x"C0C0BFA4F9C08099",
-21083 => x"C0C0BFA4F9C080B0",
-21082 => x"C0C0BFA4F9C080A4",
-21081 => x"C0C0BFA4F9C080F9",
-21080 => x"C0C0BFA4F9C080C0",
-21079 => x"C0C0BFA4F9C0F890",
-21078 => x"C0C0BFA4F9C0F880",
-21077 => x"C0C0BFA4F9C0F8F8",
-21076 => x"C0C0BFA4F9C0F882",
-21075 => x"C0C0BFA4F9C0F892",
-21074 => x"C0C0BFA4F9C0F899",
-21073 => x"C0C0BFA4F9C0F8B0",
-21072 => x"C0C0BFA4F9C0F8A4",
-21071 => x"C0C0BFA4F9C0F8F9",
-21070 => x"C0C0BFA4F9C0F8C0",
-21069 => x"C0C0BFA4F9C08290",
-21068 => x"C0C0BFA4F9C08280",
-21067 => x"C0C0BFA4F9C082F8",
-21066 => x"C0C0BFA4F9C08282",
-21065 => x"C0C0BFA4F9C08292",
-21064 => x"C0C0BFA4F9C08299",
-21063 => x"C0C0BFA4F9C082B0",
-21062 => x"C0C0BFA4F9C082A4",
-21061 => x"C0C0BFA4F9C082F9",
-21060 => x"C0C0BFA4F9C082C0",
-21059 => x"C0C0BFA4F9C09290",
-21058 => x"C0C0BFA4F9C09280",
-21057 => x"C0C0BFA4F9C092F8",
-21056 => x"C0C0BFA4F9C09282",
-21055 => x"C0C0BFA4F9C09292",
-21054 => x"C0C0BFA4F9C09299",
-21053 => x"C0C0BFA4F9C092B0",
-21052 => x"C0C0BFA4F9C092A4",
-21051 => x"C0C0BFA4F9C092F9",
-21050 => x"C0C0BFA4F9C092C0",
-21049 => x"C0C0BFA4F9C09990",
-21048 => x"C0C0BFA4F9C09980",
-21047 => x"C0C0BFA4F9C099F8",
-21046 => x"C0C0BFA4F9C09982",
-21045 => x"C0C0BFA4F9C09992",
-21044 => x"C0C0BFA4F9C09999",
-21043 => x"C0C0BFA4F9C099B0",
-21042 => x"C0C0BFA4F9C099A4",
-21041 => x"C0C0BFA4F9C099F9",
-21040 => x"C0C0BFA4F9C099C0",
-21039 => x"C0C0BFA4F9C0B090",
-21038 => x"C0C0BFA4F9C0B080",
-21037 => x"C0C0BFA4F9C0B0F8",
-21036 => x"C0C0BFA4F9C0B082",
-21035 => x"C0C0BFA4F9C0B092",
-21034 => x"C0C0BFA4F9C0B099",
-21033 => x"C0C0BFA4F9C0B0B0",
-21032 => x"C0C0BFA4F9C0B0A4",
-21031 => x"C0C0BFA4F9C0B0F9",
-21030 => x"C0C0BFA4F9C0B0C0",
-21029 => x"C0C0BFA4F9C0A490",
-21028 => x"C0C0BFA4F9C0A480",
-21027 => x"C0C0BFA4F9C0A4F8",
-21026 => x"C0C0BFA4F9C0A482",
-21025 => x"C0C0BFA4F9C0A492",
-21024 => x"C0C0BFA4F9C0A499",
-21023 => x"C0C0BFA4F9C0A4B0",
-21022 => x"C0C0BFA4F9C0A4A4",
-21021 => x"C0C0BFA4F9C0A4F9",
-21020 => x"C0C0BFA4F9C0A4C0",
-21019 => x"C0C0BFA4F9C0F990",
-21018 => x"C0C0BFA4F9C0F980",
-21017 => x"C0C0BFA4F9C0F9F8",
-21016 => x"C0C0BFA4F9C0F982",
-21015 => x"C0C0BFA4F9C0F992",
-21014 => x"C0C0BFA4F9C0F999",
-21013 => x"C0C0BFA4F9C0F9B0",
-21012 => x"C0C0BFA4F9C0F9A4",
-21011 => x"C0C0BFA4F9C0F9F9",
-21010 => x"C0C0BFA4F9C0F9C0",
-21009 => x"C0C0BFA4F9C0C090",
-21008 => x"C0C0BFA4F9C0C080",
-21007 => x"C0C0BFA4F9C0C0F8",
-21006 => x"C0C0BFA4F9C0C082",
-21005 => x"C0C0BFA4F9C0C092",
-21004 => x"C0C0BFA4F9C0C099",
-21003 => x"C0C0BFA4F9C0C0B0",
-21002 => x"C0C0BFA4F9C0C0A4",
-21001 => x"C0C0BFA4F9C0C0F9",
-21000 => x"C0C0BFA4F9C0C0C0",
-20999 => x"C0C0BFA4C0909090",
-20998 => x"C0C0BFA4C0909080",
-20997 => x"C0C0BFA4C09090F8",
-20996 => x"C0C0BFA4C0909082",
-20995 => x"C0C0BFA4C0909092",
-20994 => x"C0C0BFA4C0909099",
-20993 => x"C0C0BFA4C09090B0",
-20992 => x"C0C0BFA4C09090A4",
-20991 => x"C0C0BFA4C09090F9",
-20990 => x"C0C0BFA4C09090C0",
-20989 => x"C0C0BFA4C0908090",
-20988 => x"C0C0BFA4C0908080",
-20987 => x"C0C0BFA4C09080F8",
-20986 => x"C0C0BFA4C0908082",
-20985 => x"C0C0BFA4C0908092",
-20984 => x"C0C0BFA4C0908099",
-20983 => x"C0C0BFA4C09080B0",
-20982 => x"C0C0BFA4C09080A4",
-20981 => x"C0C0BFA4C09080F9",
-20980 => x"C0C0BFA4C09080C0",
-20979 => x"C0C0BFA4C090F890",
-20978 => x"C0C0BFA4C090F880",
-20977 => x"C0C0BFA4C090F8F8",
-20976 => x"C0C0BFA4C090F882",
-20975 => x"C0C0BFA4C090F892",
-20974 => x"C0C0BFA4C090F899",
-20973 => x"C0C0BFA4C090F8B0",
-20972 => x"C0C0BFA4C090F8A4",
-20971 => x"C0C0BFA4C090F8F9",
-20970 => x"C0C0BFA4C090F8C0",
-20969 => x"C0C0BFA4C0908290",
-20968 => x"C0C0BFA4C0908280",
-20967 => x"C0C0BFA4C09082F8",
-20966 => x"C0C0BFA4C0908282",
-20965 => x"C0C0BFA4C0908292",
-20964 => x"C0C0BFA4C0908299",
-20963 => x"C0C0BFA4C09082B0",
-20962 => x"C0C0BFA4C09082A4",
-20961 => x"C0C0BFA4C09082F9",
-20960 => x"C0C0BFA4C09082C0",
-20959 => x"C0C0BFA4C0909290",
-20958 => x"C0C0BFA4C0909280",
-20957 => x"C0C0BFA4C09092F8",
-20956 => x"C0C0BFA4C0909282",
-20955 => x"C0C0BFA4C0909292",
-20954 => x"C0C0BFA4C0909299",
-20953 => x"C0C0BFA4C09092B0",
-20952 => x"C0C0BFA4C09092A4",
-20951 => x"C0C0BFA4C09092F9",
-20950 => x"C0C0BFA4C09092C0",
-20949 => x"C0C0BFA4C0909990",
-20948 => x"C0C0BFA4C0909980",
-20947 => x"C0C0BFA4C09099F8",
-20946 => x"C0C0BFA4C0909982",
-20945 => x"C0C0BFA4C0909992",
-20944 => x"C0C0BFA4C0909999",
-20943 => x"C0C0BFA4C09099B0",
-20942 => x"C0C0BFA4C09099A4",
-20941 => x"C0C0BFA4C09099F9",
-20940 => x"C0C0BFA4C09099C0",
-20939 => x"C0C0BFA4C090B090",
-20938 => x"C0C0BFA4C090B080",
-20937 => x"C0C0BFA4C090B0F8",
-20936 => x"C0C0BFA4C090B082",
-20935 => x"C0C0BFA4C090B092",
-20934 => x"C0C0BFA4C090B099",
-20933 => x"C0C0BFA4C090B0B0",
-20932 => x"C0C0BFA4C090B0A4",
-20931 => x"C0C0BFA4C090B0F9",
-20930 => x"C0C0BFA4C090B0C0",
-20929 => x"C0C0BFA4C090A490",
-20928 => x"C0C0BFA4C090A480",
-20927 => x"C0C0BFA4C090A4F8",
-20926 => x"C0C0BFA4C090A482",
-20925 => x"C0C0BFA4C090A492",
-20924 => x"C0C0BFA4C090A499",
-20923 => x"C0C0BFA4C090A4B0",
-20922 => x"C0C0BFA4C090A4A4",
-20921 => x"C0C0BFA4C090A4F9",
-20920 => x"C0C0BFA4C090A4C0",
-20919 => x"C0C0BFA4C090F990",
-20918 => x"C0C0BFA4C090F980",
-20917 => x"C0C0BFA4C090F9F8",
-20916 => x"C0C0BFA4C090F982",
-20915 => x"C0C0BFA4C090F992",
-20914 => x"C0C0BFA4C090F999",
-20913 => x"C0C0BFA4C090F9B0",
-20912 => x"C0C0BFA4C090F9A4",
-20911 => x"C0C0BFA4C090F9F9",
-20910 => x"C0C0BFA4C090F9C0",
-20909 => x"C0C0BFA4C090C090",
-20908 => x"C0C0BFA4C090C080",
-20907 => x"C0C0BFA4C090C0F8",
-20906 => x"C0C0BFA4C090C082",
-20905 => x"C0C0BFA4C090C092",
-20904 => x"C0C0BFA4C090C099",
-20903 => x"C0C0BFA4C090C0B0",
-20902 => x"C0C0BFA4C090C0A4",
-20901 => x"C0C0BFA4C090C0F9",
-20900 => x"C0C0BFA4C090C0C0",
-20899 => x"C0C0BFA4C0809090",
-20898 => x"C0C0BFA4C0809080",
-20897 => x"C0C0BFA4C08090F8",
-20896 => x"C0C0BFA4C0809082",
-20895 => x"C0C0BFA4C0809092",
-20894 => x"C0C0BFA4C0809099",
-20893 => x"C0C0BFA4C08090B0",
-20892 => x"C0C0BFA4C08090A4",
-20891 => x"C0C0BFA4C08090F9",
-20890 => x"C0C0BFA4C08090C0",
-20889 => x"C0C0BFA4C0808090",
-20888 => x"C0C0BFA4C0808080",
-20887 => x"C0C0BFA4C08080F8",
-20886 => x"C0C0BFA4C0808082",
-20885 => x"C0C0BFA4C0808092",
-20884 => x"C0C0BFA4C0808099",
-20883 => x"C0C0BFA4C08080B0",
-20882 => x"C0C0BFA4C08080A4",
-20881 => x"C0C0BFA4C08080F9",
-20880 => x"C0C0BFA4C08080C0",
-20879 => x"C0C0BFA4C080F890",
-20878 => x"C0C0BFA4C080F880",
-20877 => x"C0C0BFA4C080F8F8",
-20876 => x"C0C0BFA4C080F882",
-20875 => x"C0C0BFA4C080F892",
-20874 => x"C0C0BFA4C080F899",
-20873 => x"C0C0BFA4C080F8B0",
-20872 => x"C0C0BFA4C080F8A4",
-20871 => x"C0C0BFA4C080F8F9",
-20870 => x"C0C0BFA4C080F8C0",
-20869 => x"C0C0BFA4C0808290",
-20868 => x"C0C0BFA4C0808280",
-20867 => x"C0C0BFA4C08082F8",
-20866 => x"C0C0BFA4C0808282",
-20865 => x"C0C0BFA4C0808292",
-20864 => x"C0C0BFA4C0808299",
-20863 => x"C0C0BFA4C08082B0",
-20862 => x"C0C0BFA4C08082A4",
-20861 => x"C0C0BFA4C08082F9",
-20860 => x"C0C0BFA4C08082C0",
-20859 => x"C0C0BFA4C0809290",
-20858 => x"C0C0BFA4C0809280",
-20857 => x"C0C0BFA4C08092F8",
-20856 => x"C0C0BFA4C0809282",
-20855 => x"C0C0BFA4C0809292",
-20854 => x"C0C0BFA4C0809299",
-20853 => x"C0C0BFA4C08092B0",
-20852 => x"C0C0BFA4C08092A4",
-20851 => x"C0C0BFA4C08092F9",
-20850 => x"C0C0BFA4C08092C0",
-20849 => x"C0C0BFA4C0809990",
-20848 => x"C0C0BFA4C0809980",
-20847 => x"C0C0BFA4C08099F8",
-20846 => x"C0C0BFA4C0809982",
-20845 => x"C0C0BFA4C0809992",
-20844 => x"C0C0BFA4C0809999",
-20843 => x"C0C0BFA4C08099B0",
-20842 => x"C0C0BFA4C08099A4",
-20841 => x"C0C0BFA4C08099F9",
-20840 => x"C0C0BFA4C08099C0",
-20839 => x"C0C0BFA4C080B090",
-20838 => x"C0C0BFA4C080B080",
-20837 => x"C0C0BFA4C080B0F8",
-20836 => x"C0C0BFA4C080B082",
-20835 => x"C0C0BFA4C080B092",
-20834 => x"C0C0BFA4C080B099",
-20833 => x"C0C0BFA4C080B0B0",
-20832 => x"C0C0BFA4C080B0A4",
-20831 => x"C0C0BFA4C080B0F9",
-20830 => x"C0C0BFA4C080B0C0",
-20829 => x"C0C0BFA4C080A490",
-20828 => x"C0C0BFA4C080A480",
-20827 => x"C0C0BFA4C080A4F8",
-20826 => x"C0C0BFA4C080A482",
-20825 => x"C0C0BFA4C080A492",
-20824 => x"C0C0BFA4C080A499",
-20823 => x"C0C0BFA4C080A4B0",
-20822 => x"C0C0BFA4C080A4A4",
-20821 => x"C0C0BFA4C080A4F9",
-20820 => x"C0C0BFA4C080A4C0",
-20819 => x"C0C0BFA4C080F990",
-20818 => x"C0C0BFA4C080F980",
-20817 => x"C0C0BFA4C080F9F8",
-20816 => x"C0C0BFA4C080F982",
-20815 => x"C0C0BFA4C080F992",
-20814 => x"C0C0BFA4C080F999",
-20813 => x"C0C0BFA4C080F9B0",
-20812 => x"C0C0BFA4C080F9A4",
-20811 => x"C0C0BFA4C080F9F9",
-20810 => x"C0C0BFA4C080F9C0",
-20809 => x"C0C0BFA4C080C090",
-20808 => x"C0C0BFA4C080C080",
-20807 => x"C0C0BFA4C080C0F8",
-20806 => x"C0C0BFA4C080C082",
-20805 => x"C0C0BFA4C080C092",
-20804 => x"C0C0BFA4C080C099",
-20803 => x"C0C0BFA4C080C0B0",
-20802 => x"C0C0BFA4C080C0A4",
-20801 => x"C0C0BFA4C080C0F9",
-20800 => x"C0C0BFA4C080C0C0",
-20799 => x"C0C0BFA4C0F89090",
-20798 => x"C0C0BFA4C0F89080",
-20797 => x"C0C0BFA4C0F890F8",
-20796 => x"C0C0BFA4C0F89082",
-20795 => x"C0C0BFA4C0F89092",
-20794 => x"C0C0BFA4C0F89099",
-20793 => x"C0C0BFA4C0F890B0",
-20792 => x"C0C0BFA4C0F890A4",
-20791 => x"C0C0BFA4C0F890F9",
-20790 => x"C0C0BFA4C0F890C0",
-20789 => x"C0C0BFA4C0F88090",
-20788 => x"C0C0BFA4C0F88080",
-20787 => x"C0C0BFA4C0F880F8",
-20786 => x"C0C0BFA4C0F88082",
-20785 => x"C0C0BFA4C0F88092",
-20784 => x"C0C0BFA4C0F88099",
-20783 => x"C0C0BFA4C0F880B0",
-20782 => x"C0C0BFA4C0F880A4",
-20781 => x"C0C0BFA4C0F880F9",
-20780 => x"C0C0BFA4C0F880C0",
-20779 => x"C0C0BFA4C0F8F890",
-20778 => x"C0C0BFA4C0F8F880",
-20777 => x"C0C0BFA4C0F8F8F8",
-20776 => x"C0C0BFA4C0F8F882",
-20775 => x"C0C0BFA4C0F8F892",
-20774 => x"C0C0BFA4C0F8F899",
-20773 => x"C0C0BFA4C0F8F8B0",
-20772 => x"C0C0BFA4C0F8F8A4",
-20771 => x"C0C0BFA4C0F8F8F9",
-20770 => x"C0C0BFA4C0F8F8C0",
-20769 => x"C0C0BFA4C0F88290",
-20768 => x"C0C0BFA4C0F88280",
-20767 => x"C0C0BFA4C0F882F8",
-20766 => x"C0C0BFA4C0F88282",
-20765 => x"C0C0BFA4C0F88292",
-20764 => x"C0C0BFA4C0F88299",
-20763 => x"C0C0BFA4C0F882B0",
-20762 => x"C0C0BFA4C0F882A4",
-20761 => x"C0C0BFA4C0F882F9",
-20760 => x"C0C0BFA4C0F882C0",
-20759 => x"C0C0BFA4C0F89290",
-20758 => x"C0C0BFA4C0F89280",
-20757 => x"C0C0BFA4C0F892F8",
-20756 => x"C0C0BFA4C0F89282",
-20755 => x"C0C0BFA4C0F89292",
-20754 => x"C0C0BFA4C0F89299",
-20753 => x"C0C0BFA4C0F892B0",
-20752 => x"C0C0BFA4C0F892A4",
-20751 => x"C0C0BFA4C0F892F9",
-20750 => x"C0C0BFA4C0F892C0",
-20749 => x"C0C0BFA4C0F89990",
-20748 => x"C0C0BFA4C0F89980",
-20747 => x"C0C0BFA4C0F899F8",
-20746 => x"C0C0BFA4C0F89982",
-20745 => x"C0C0BFA4C0F89992",
-20744 => x"C0C0BFA4C0F89999",
-20743 => x"C0C0BFA4C0F899B0",
-20742 => x"C0C0BFA4C0F899A4",
-20741 => x"C0C0BFA4C0F899F9",
-20740 => x"C0C0BFA4C0F899C0",
-20739 => x"C0C0BFA4C0F8B090",
-20738 => x"C0C0BFA4C0F8B080",
-20737 => x"C0C0BFA4C0F8B0F8",
-20736 => x"C0C0BFA4C0F8B082",
-20735 => x"C0C0BFA4C0F8B092",
-20734 => x"C0C0BFA4C0F8B099",
-20733 => x"C0C0BFA4C0F8B0B0",
-20732 => x"C0C0BFA4C0F8B0A4",
-20731 => x"C0C0BFA4C0F8B0F9",
-20730 => x"C0C0BFA4C0F8B0C0",
-20729 => x"C0C0BFA4C0F8A490",
-20728 => x"C0C0BFA4C0F8A480",
-20727 => x"C0C0BFA4C0F8A4F8",
-20726 => x"C0C0BFA4C0F8A482",
-20725 => x"C0C0BFA4C0F8A492",
-20724 => x"C0C0BFA4C0F8A499",
-20723 => x"C0C0BFA4C0F8A4B0",
-20722 => x"C0C0BFA4C0F8A4A4",
-20721 => x"C0C0BFA4C0F8A4F9",
-20720 => x"C0C0BFA4C0F8A4C0",
-20719 => x"C0C0BFA4C0F8F990",
-20718 => x"C0C0BFA4C0F8F980",
-20717 => x"C0C0BFA4C0F8F9F8",
-20716 => x"C0C0BFA4C0F8F982",
-20715 => x"C0C0BFA4C0F8F992",
-20714 => x"C0C0BFA4C0F8F999",
-20713 => x"C0C0BFA4C0F8F9B0",
-20712 => x"C0C0BFA4C0F8F9A4",
-20711 => x"C0C0BFA4C0F8F9F9",
-20710 => x"C0C0BFA4C0F8F9C0",
-20709 => x"C0C0BFA4C0F8C090",
-20708 => x"C0C0BFA4C0F8C080",
-20707 => x"C0C0BFA4C0F8C0F8",
-20706 => x"C0C0BFA4C0F8C082",
-20705 => x"C0C0BFA4C0F8C092",
-20704 => x"C0C0BFA4C0F8C099",
-20703 => x"C0C0BFA4C0F8C0B0",
-20702 => x"C0C0BFA4C0F8C0A4",
-20701 => x"C0C0BFA4C0F8C0F9",
-20700 => x"C0C0BFA4C0F8C0C0",
-20699 => x"C0C0BFA4C0829090",
-20698 => x"C0C0BFA4C0829080",
-20697 => x"C0C0BFA4C08290F8",
-20696 => x"C0C0BFA4C0829082",
-20695 => x"C0C0BFA4C0829092",
-20694 => x"C0C0BFA4C0829099",
-20693 => x"C0C0BFA4C08290B0",
-20692 => x"C0C0BFA4C08290A4",
-20691 => x"C0C0BFA4C08290F9",
-20690 => x"C0C0BFA4C08290C0",
-20689 => x"C0C0BFA4C0828090",
-20688 => x"C0C0BFA4C0828080",
-20687 => x"C0C0BFA4C08280F8",
-20686 => x"C0C0BFA4C0828082",
-20685 => x"C0C0BFA4C0828092",
-20684 => x"C0C0BFA4C0828099",
-20683 => x"C0C0BFA4C08280B0",
-20682 => x"C0C0BFA4C08280A4",
-20681 => x"C0C0BFA4C08280F9",
-20680 => x"C0C0BFA4C08280C0",
-20679 => x"C0C0BFA4C082F890",
-20678 => x"C0C0BFA4C082F880",
-20677 => x"C0C0BFA4C082F8F8",
-20676 => x"C0C0BFA4C082F882",
-20675 => x"C0C0BFA4C082F892",
-20674 => x"C0C0BFA4C082F899",
-20673 => x"C0C0BFA4C082F8B0",
-20672 => x"C0C0BFA4C082F8A4",
-20671 => x"C0C0BFA4C082F8F9",
-20670 => x"C0C0BFA4C082F8C0",
-20669 => x"C0C0BFA4C0828290",
-20668 => x"C0C0BFA4C0828280",
-20667 => x"C0C0BFA4C08282F8",
-20666 => x"C0C0BFA4C0828282",
-20665 => x"C0C0BFA4C0828292",
-20664 => x"C0C0BFA4C0828299",
-20663 => x"C0C0BFA4C08282B0",
-20662 => x"C0C0BFA4C08282A4",
-20661 => x"C0C0BFA4C08282F9",
-20660 => x"C0C0BFA4C08282C0",
-20659 => x"C0C0BFA4C0829290",
-20658 => x"C0C0BFA4C0829280",
-20657 => x"C0C0BFA4C08292F8",
-20656 => x"C0C0BFA4C0829282",
-20655 => x"C0C0BFA4C0829292",
-20654 => x"C0C0BFA4C0829299",
-20653 => x"C0C0BFA4C08292B0",
-20652 => x"C0C0BFA4C08292A4",
-20651 => x"C0C0BFA4C08292F9",
-20650 => x"C0C0BFA4C08292C0",
-20649 => x"C0C0BFA4C0829990",
-20648 => x"C0C0BFA4C0829980",
-20647 => x"C0C0BFA4C08299F8",
-20646 => x"C0C0BFA4C0829982",
-20645 => x"C0C0BFA4C0829992",
-20644 => x"C0C0BFA4C0829999",
-20643 => x"C0C0BFA4C08299B0",
-20642 => x"C0C0BFA4C08299A4",
-20641 => x"C0C0BFA4C08299F9",
-20640 => x"C0C0BFA4C08299C0",
-20639 => x"C0C0BFA4C082B090",
-20638 => x"C0C0BFA4C082B080",
-20637 => x"C0C0BFA4C082B0F8",
-20636 => x"C0C0BFA4C082B082",
-20635 => x"C0C0BFA4C082B092",
-20634 => x"C0C0BFA4C082B099",
-20633 => x"C0C0BFA4C082B0B0",
-20632 => x"C0C0BFA4C082B0A4",
-20631 => x"C0C0BFA4C082B0F9",
-20630 => x"C0C0BFA4C082B0C0",
-20629 => x"C0C0BFA4C082A490",
-20628 => x"C0C0BFA4C082A480",
-20627 => x"C0C0BFA4C082A4F8",
-20626 => x"C0C0BFA4C082A482",
-20625 => x"C0C0BFA4C082A492",
-20624 => x"C0C0BFA4C082A499",
-20623 => x"C0C0BFA4C082A4B0",
-20622 => x"C0C0BFA4C082A4A4",
-20621 => x"C0C0BFA4C082A4F9",
-20620 => x"C0C0BFA4C082A4C0",
-20619 => x"C0C0BFA4C082F990",
-20618 => x"C0C0BFA4C082F980",
-20617 => x"C0C0BFA4C082F9F8",
-20616 => x"C0C0BFA4C082F982",
-20615 => x"C0C0BFA4C082F992",
-20614 => x"C0C0BFA4C082F999",
-20613 => x"C0C0BFA4C082F9B0",
-20612 => x"C0C0BFA4C082F9A4",
-20611 => x"C0C0BFA4C082F9F9",
-20610 => x"C0C0BFA4C082F9C0",
-20609 => x"C0C0BFA4C082C090",
-20608 => x"C0C0BFA4C082C080",
-20607 => x"C0C0BFA4C082C0F8",
-20606 => x"C0C0BFA4C082C082",
-20605 => x"C0C0BFA4C082C092",
-20604 => x"C0C0BFA4C082C099",
-20603 => x"C0C0BFA4C082C0B0",
-20602 => x"C0C0BFA4C082C0A4",
-20601 => x"C0C0BFA4C082C0F9",
-20600 => x"C0C0BFA4C082C0C0",
-20599 => x"C0C0BFA4C0929090",
-20598 => x"C0C0BFA4C0929080",
-20597 => x"C0C0BFA4C09290F8",
-20596 => x"C0C0BFA4C0929082",
-20595 => x"C0C0BFA4C0929092",
-20594 => x"C0C0BFA4C0929099",
-20593 => x"C0C0BFA4C09290B0",
-20592 => x"C0C0BFA4C09290A4",
-20591 => x"C0C0BFA4C09290F9",
-20590 => x"C0C0BFA4C09290C0",
-20589 => x"C0C0BFA4C0928090",
-20588 => x"C0C0BFA4C0928080",
-20587 => x"C0C0BFA4C09280F8",
-20586 => x"C0C0BFA4C0928082",
-20585 => x"C0C0BFA4C0928092",
-20584 => x"C0C0BFA4C0928099",
-20583 => x"C0C0BFA4C09280B0",
-20582 => x"C0C0BFA4C09280A4",
-20581 => x"C0C0BFA4C09280F9",
-20580 => x"C0C0BFA4C09280C0",
-20579 => x"C0C0BFA4C092F890",
-20578 => x"C0C0BFA4C092F880",
-20577 => x"C0C0BFA4C092F8F8",
-20576 => x"C0C0BFA4C092F882",
-20575 => x"C0C0BFA4C092F892",
-20574 => x"C0C0BFA4C092F899",
-20573 => x"C0C0BFA4C092F8B0",
-20572 => x"C0C0BFA4C092F8A4",
-20571 => x"C0C0BFA4C092F8F9",
-20570 => x"C0C0BFA4C092F8C0",
-20569 => x"C0C0BFA4C0928290",
-20568 => x"C0C0BFA4C0928280",
-20567 => x"C0C0BFA4C09282F8",
-20566 => x"C0C0BFA4C0928282",
-20565 => x"C0C0BFA4C0928292",
-20564 => x"C0C0BFA4C0928299",
-20563 => x"C0C0BFA4C09282B0",
-20562 => x"C0C0BFA4C09282A4",
-20561 => x"C0C0BFA4C09282F9",
-20560 => x"C0C0BFA4C09282C0",
-20559 => x"C0C0BFA4C0929290",
-20558 => x"C0C0BFA4C0929280",
-20557 => x"C0C0BFA4C09292F8",
-20556 => x"C0C0BFA4C0929282",
-20555 => x"C0C0BFA4C0929292",
-20554 => x"C0C0BFA4C0929299",
-20553 => x"C0C0BFA4C09292B0",
-20552 => x"C0C0BFA4C09292A4",
-20551 => x"C0C0BFA4C09292F9",
-20550 => x"C0C0BFA4C09292C0",
-20549 => x"C0C0BFA4C0929990",
-20548 => x"C0C0BFA4C0929980",
-20547 => x"C0C0BFA4C09299F8",
-20546 => x"C0C0BFA4C0929982",
-20545 => x"C0C0BFA4C0929992",
-20544 => x"C0C0BFA4C0929999",
-20543 => x"C0C0BFA4C09299B0",
-20542 => x"C0C0BFA4C09299A4",
-20541 => x"C0C0BFA4C09299F9",
-20540 => x"C0C0BFA4C09299C0",
-20539 => x"C0C0BFA4C092B090",
-20538 => x"C0C0BFA4C092B080",
-20537 => x"C0C0BFA4C092B0F8",
-20536 => x"C0C0BFA4C092B082",
-20535 => x"C0C0BFA4C092B092",
-20534 => x"C0C0BFA4C092B099",
-20533 => x"C0C0BFA4C092B0B0",
-20532 => x"C0C0BFA4C092B0A4",
-20531 => x"C0C0BFA4C092B0F9",
-20530 => x"C0C0BFA4C092B0C0",
-20529 => x"C0C0BFA4C092A490",
-20528 => x"C0C0BFA4C092A480",
-20527 => x"C0C0BFA4C092A4F8",
-20526 => x"C0C0BFA4C092A482",
-20525 => x"C0C0BFA4C092A492",
-20524 => x"C0C0BFA4C092A499",
-20523 => x"C0C0BFA4C092A4B0",
-20522 => x"C0C0BFA4C092A4A4",
-20521 => x"C0C0BFA4C092A4F9",
-20520 => x"C0C0BFA4C092A4C0",
-20519 => x"C0C0BFA4C092F990",
-20518 => x"C0C0BFA4C092F980",
-20517 => x"C0C0BFA4C092F9F8",
-20516 => x"C0C0BFA4C092F982",
-20515 => x"C0C0BFA4C092F992",
-20514 => x"C0C0BFA4C092F999",
-20513 => x"C0C0BFA4C092F9B0",
-20512 => x"C0C0BFA4C092F9A4",
-20511 => x"C0C0BFA4C092F9F9",
-20510 => x"C0C0BFA4C092F9C0",
-20509 => x"C0C0BFA4C092C090",
-20508 => x"C0C0BFA4C092C080",
-20507 => x"C0C0BFA4C092C0F8",
-20506 => x"C0C0BFA4C092C082",
-20505 => x"C0C0BFA4C092C092",
-20504 => x"C0C0BFA4C092C099",
-20503 => x"C0C0BFA4C092C0B0",
-20502 => x"C0C0BFA4C092C0A4",
-20501 => x"C0C0BFA4C092C0F9",
-20500 => x"C0C0BFA4C092C0C0",
-20499 => x"C0C0BFA4C0999090",
-20498 => x"C0C0BFA4C0999080",
-20497 => x"C0C0BFA4C09990F8",
-20496 => x"C0C0BFA4C0999082",
-20495 => x"C0C0BFA4C0999092",
-20494 => x"C0C0BFA4C0999099",
-20493 => x"C0C0BFA4C09990B0",
-20492 => x"C0C0BFA4C09990A4",
-20491 => x"C0C0BFA4C09990F9",
-20490 => x"C0C0BFA4C09990C0",
-20489 => x"C0C0BFA4C0998090",
-20488 => x"C0C0BFA4C0998080",
-20487 => x"C0C0BFA4C09980F8",
-20486 => x"C0C0BFA4C0998082",
-20485 => x"C0C0BFA4C0998092",
-20484 => x"C0C0BFA4C0998099",
-20483 => x"C0C0BFA4C09980B0",
-20482 => x"C0C0BFA4C09980A4",
-20481 => x"C0C0BFA4C09980F9",
-20480 => x"C0C0BFA4C09980C0",
-20479 => x"C0C0BFA4C099F890",
-20478 => x"C0C0BFA4C099F880",
-20477 => x"C0C0BFA4C099F8F8",
-20476 => x"C0C0BFA4C099F882",
-20475 => x"C0C0BFA4C099F892",
-20474 => x"C0C0BFA4C099F899",
-20473 => x"C0C0BFA4C099F8B0",
-20472 => x"C0C0BFA4C099F8A4",
-20471 => x"C0C0BFA4C099F8F9",
-20470 => x"C0C0BFA4C099F8C0",
-20469 => x"C0C0BFA4C0998290",
-20468 => x"C0C0BFA4C0998280",
-20467 => x"C0C0BFA4C09982F8",
-20466 => x"C0C0BFA4C0998282",
-20465 => x"C0C0BFA4C0998292",
-20464 => x"C0C0BFA4C0998299",
-20463 => x"C0C0BFA4C09982B0",
-20462 => x"C0C0BFA4C09982A4",
-20461 => x"C0C0BFA4C09982F9",
-20460 => x"C0C0BFA4C09982C0",
-20459 => x"C0C0BFA4C0999290",
-20458 => x"C0C0BFA4C0999280",
-20457 => x"C0C0BFA4C09992F8",
-20456 => x"C0C0BFA4C0999282",
-20455 => x"C0C0BFA4C0999292",
-20454 => x"C0C0BFA4C0999299",
-20453 => x"C0C0BFA4C09992B0",
-20452 => x"C0C0BFA4C09992A4",
-20451 => x"C0C0BFA4C09992F9",
-20450 => x"C0C0BFA4C09992C0",
-20449 => x"C0C0BFA4C0999990",
-20448 => x"C0C0BFA4C0999980",
-20447 => x"C0C0BFA4C09999F8",
-20446 => x"C0C0BFA4C0999982",
-20445 => x"C0C0BFA4C0999992",
-20444 => x"C0C0BFA4C0999999",
-20443 => x"C0C0BFA4C09999B0",
-20442 => x"C0C0BFA4C09999A4",
-20441 => x"C0C0BFA4C09999F9",
-20440 => x"C0C0BFA4C09999C0",
-20439 => x"C0C0BFA4C099B090",
-20438 => x"C0C0BFA4C099B080",
-20437 => x"C0C0BFA4C099B0F8",
-20436 => x"C0C0BFA4C099B082",
-20435 => x"C0C0BFA4C099B092",
-20434 => x"C0C0BFA4C099B099",
-20433 => x"C0C0BFA4C099B0B0",
-20432 => x"C0C0BFA4C099B0A4",
-20431 => x"C0C0BFA4C099B0F9",
-20430 => x"C0C0BFA4C099B0C0",
-20429 => x"C0C0BFA4C099A490",
-20428 => x"C0C0BFA4C099A480",
-20427 => x"C0C0BFA4C099A4F8",
-20426 => x"C0C0BFA4C099A482",
-20425 => x"C0C0BFA4C099A492",
-20424 => x"C0C0BFA4C099A499",
-20423 => x"C0C0BFA4C099A4B0",
-20422 => x"C0C0BFA4C099A4A4",
-20421 => x"C0C0BFA4C099A4F9",
-20420 => x"C0C0BFA4C099A4C0",
-20419 => x"C0C0BFA4C099F990",
-20418 => x"C0C0BFA4C099F980",
-20417 => x"C0C0BFA4C099F9F8",
-20416 => x"C0C0BFA4C099F982",
-20415 => x"C0C0BFA4C099F992",
-20414 => x"C0C0BFA4C099F999",
-20413 => x"C0C0BFA4C099F9B0",
-20412 => x"C0C0BFA4C099F9A4",
-20411 => x"C0C0BFA4C099F9F9",
-20410 => x"C0C0BFA4C099F9C0",
-20409 => x"C0C0BFA4C099C090",
-20408 => x"C0C0BFA4C099C080",
-20407 => x"C0C0BFA4C099C0F8",
-20406 => x"C0C0BFA4C099C082",
-20405 => x"C0C0BFA4C099C092",
-20404 => x"C0C0BFA4C099C099",
-20403 => x"C0C0BFA4C099C0B0",
-20402 => x"C0C0BFA4C099C0A4",
-20401 => x"C0C0BFA4C099C0F9",
-20400 => x"C0C0BFA4C099C0C0",
-20399 => x"C0C0BFA4C0B09090",
-20398 => x"C0C0BFA4C0B09080",
-20397 => x"C0C0BFA4C0B090F8",
-20396 => x"C0C0BFA4C0B09082",
-20395 => x"C0C0BFA4C0B09092",
-20394 => x"C0C0BFA4C0B09099",
-20393 => x"C0C0BFA4C0B090B0",
-20392 => x"C0C0BFA4C0B090A4",
-20391 => x"C0C0BFA4C0B090F9",
-20390 => x"C0C0BFA4C0B090C0",
-20389 => x"C0C0BFA4C0B08090",
-20388 => x"C0C0BFA4C0B08080",
-20387 => x"C0C0BFA4C0B080F8",
-20386 => x"C0C0BFA4C0B08082",
-20385 => x"C0C0BFA4C0B08092",
-20384 => x"C0C0BFA4C0B08099",
-20383 => x"C0C0BFA4C0B080B0",
-20382 => x"C0C0BFA4C0B080A4",
-20381 => x"C0C0BFA4C0B080F9",
-20380 => x"C0C0BFA4C0B080C0",
-20379 => x"C0C0BFA4C0B0F890",
-20378 => x"C0C0BFA4C0B0F880",
-20377 => x"C0C0BFA4C0B0F8F8",
-20376 => x"C0C0BFA4C0B0F882",
-20375 => x"C0C0BFA4C0B0F892",
-20374 => x"C0C0BFA4C0B0F899",
-20373 => x"C0C0BFA4C0B0F8B0",
-20372 => x"C0C0BFA4C0B0F8A4",
-20371 => x"C0C0BFA4C0B0F8F9",
-20370 => x"C0C0BFA4C0B0F8C0",
-20369 => x"C0C0BFA4C0B08290",
-20368 => x"C0C0BFA4C0B08280",
-20367 => x"C0C0BFA4C0B082F8",
-20366 => x"C0C0BFA4C0B08282",
-20365 => x"C0C0BFA4C0B08292",
-20364 => x"C0C0BFA4C0B08299",
-20363 => x"C0C0BFA4C0B082B0",
-20362 => x"C0C0BFA4C0B082A4",
-20361 => x"C0C0BFA4C0B082F9",
-20360 => x"C0C0BFA4C0B082C0",
-20359 => x"C0C0BFA4C0B09290",
-20358 => x"C0C0BFA4C0B09280",
-20357 => x"C0C0BFA4C0B092F8",
-20356 => x"C0C0BFA4C0B09282",
-20355 => x"C0C0BFA4C0B09292",
-20354 => x"C0C0BFA4C0B09299",
-20353 => x"C0C0BFA4C0B092B0",
-20352 => x"C0C0BFA4C0B092A4",
-20351 => x"C0C0BFA4C0B092F9",
-20350 => x"C0C0BFA4C0B092C0",
-20349 => x"C0C0BFA4C0B09990",
-20348 => x"C0C0BFA4C0B09980",
-20347 => x"C0C0BFA4C0B099F8",
-20346 => x"C0C0BFA4C0B09982",
-20345 => x"C0C0BFA4C0B09992",
-20344 => x"C0C0BFA4C0B09999",
-20343 => x"C0C0BFA4C0B099B0",
-20342 => x"C0C0BFA4C0B099A4",
-20341 => x"C0C0BFA4C0B099F9",
-20340 => x"C0C0BFA4C0B099C0",
-20339 => x"C0C0BFA4C0B0B090",
-20338 => x"C0C0BFA4C0B0B080",
-20337 => x"C0C0BFA4C0B0B0F8",
-20336 => x"C0C0BFA4C0B0B082",
-20335 => x"C0C0BFA4C0B0B092",
-20334 => x"C0C0BFA4C0B0B099",
-20333 => x"C0C0BFA4C0B0B0B0",
-20332 => x"C0C0BFA4C0B0B0A4",
-20331 => x"C0C0BFA4C0B0B0F9",
-20330 => x"C0C0BFA4C0B0B0C0",
-20329 => x"C0C0BFA4C0B0A490",
-20328 => x"C0C0BFA4C0B0A480",
-20327 => x"C0C0BFA4C0B0A4F8",
-20326 => x"C0C0BFA4C0B0A482",
-20325 => x"C0C0BFA4C0B0A492",
-20324 => x"C0C0BFA4C0B0A499",
-20323 => x"C0C0BFA4C0B0A4B0",
-20322 => x"C0C0BFA4C0B0A4A4",
-20321 => x"C0C0BFA4C0B0A4F9",
-20320 => x"C0C0BFA4C0B0A4C0",
-20319 => x"C0C0BFA4C0B0F990",
-20318 => x"C0C0BFA4C0B0F980",
-20317 => x"C0C0BFA4C0B0F9F8",
-20316 => x"C0C0BFA4C0B0F982",
-20315 => x"C0C0BFA4C0B0F992",
-20314 => x"C0C0BFA4C0B0F999",
-20313 => x"C0C0BFA4C0B0F9B0",
-20312 => x"C0C0BFA4C0B0F9A4",
-20311 => x"C0C0BFA4C0B0F9F9",
-20310 => x"C0C0BFA4C0B0F9C0",
-20309 => x"C0C0BFA4C0B0C090",
-20308 => x"C0C0BFA4C0B0C080",
-20307 => x"C0C0BFA4C0B0C0F8",
-20306 => x"C0C0BFA4C0B0C082",
-20305 => x"C0C0BFA4C0B0C092",
-20304 => x"C0C0BFA4C0B0C099",
-20303 => x"C0C0BFA4C0B0C0B0",
-20302 => x"C0C0BFA4C0B0C0A4",
-20301 => x"C0C0BFA4C0B0C0F9",
-20300 => x"C0C0BFA4C0B0C0C0",
-20299 => x"C0C0BFA4C0A49090",
-20298 => x"C0C0BFA4C0A49080",
-20297 => x"C0C0BFA4C0A490F8",
-20296 => x"C0C0BFA4C0A49082",
-20295 => x"C0C0BFA4C0A49092",
-20294 => x"C0C0BFA4C0A49099",
-20293 => x"C0C0BFA4C0A490B0",
-20292 => x"C0C0BFA4C0A490A4",
-20291 => x"C0C0BFA4C0A490F9",
-20290 => x"C0C0BFA4C0A490C0",
-20289 => x"C0C0BFA4C0A48090",
-20288 => x"C0C0BFA4C0A48080",
-20287 => x"C0C0BFA4C0A480F8",
-20286 => x"C0C0BFA4C0A48082",
-20285 => x"C0C0BFA4C0A48092",
-20284 => x"C0C0BFA4C0A48099",
-20283 => x"C0C0BFA4C0A480B0",
-20282 => x"C0C0BFA4C0A480A4",
-20281 => x"C0C0BFA4C0A480F9",
-20280 => x"C0C0BFA4C0A480C0",
-20279 => x"C0C0BFA4C0A4F890",
-20278 => x"C0C0BFA4C0A4F880",
-20277 => x"C0C0BFA4C0A4F8F8",
-20276 => x"C0C0BFA4C0A4F882",
-20275 => x"C0C0BFA4C0A4F892",
-20274 => x"C0C0BFA4C0A4F899",
-20273 => x"C0C0BFA4C0A4F8B0",
-20272 => x"C0C0BFA4C0A4F8A4",
-20271 => x"C0C0BFA4C0A4F8F9",
-20270 => x"C0C0BFA4C0A4F8C0",
-20269 => x"C0C0BFA4C0A48290",
-20268 => x"C0C0BFA4C0A48280",
-20267 => x"C0C0BFA4C0A482F8",
-20266 => x"C0C0BFA4C0A48282",
-20265 => x"C0C0BFA4C0A48292",
-20264 => x"C0C0BFA4C0A48299",
-20263 => x"C0C0BFA4C0A482B0",
-20262 => x"C0C0BFA4C0A482A4",
-20261 => x"C0C0BFA4C0A482F9",
-20260 => x"C0C0BFA4C0A482C0",
-20259 => x"C0C0BFA4C0A49290",
-20258 => x"C0C0BFA4C0A49280",
-20257 => x"C0C0BFA4C0A492F8",
-20256 => x"C0C0BFA4C0A49282",
-20255 => x"C0C0BFA4C0A49292",
-20254 => x"C0C0BFA4C0A49299",
-20253 => x"C0C0BFA4C0A492B0",
-20252 => x"C0C0BFA4C0A492A4",
-20251 => x"C0C0BFA4C0A492F9",
-20250 => x"C0C0BFA4C0A492C0",
-20249 => x"C0C0BFA4C0A49990",
-20248 => x"C0C0BFA4C0A49980",
-20247 => x"C0C0BFA4C0A499F8",
-20246 => x"C0C0BFA4C0A49982",
-20245 => x"C0C0BFA4C0A49992",
-20244 => x"C0C0BFA4C0A49999",
-20243 => x"C0C0BFA4C0A499B0",
-20242 => x"C0C0BFA4C0A499A4",
-20241 => x"C0C0BFA4C0A499F9",
-20240 => x"C0C0BFA4C0A499C0",
-20239 => x"C0C0BFA4C0A4B090",
-20238 => x"C0C0BFA4C0A4B080",
-20237 => x"C0C0BFA4C0A4B0F8",
-20236 => x"C0C0BFA4C0A4B082",
-20235 => x"C0C0BFA4C0A4B092",
-20234 => x"C0C0BFA4C0A4B099",
-20233 => x"C0C0BFA4C0A4B0B0",
-20232 => x"C0C0BFA4C0A4B0A4",
-20231 => x"C0C0BFA4C0A4B0F9",
-20230 => x"C0C0BFA4C0A4B0C0",
-20229 => x"C0C0BFA4C0A4A490",
-20228 => x"C0C0BFA4C0A4A480",
-20227 => x"C0C0BFA4C0A4A4F8",
-20226 => x"C0C0BFA4C0A4A482",
-20225 => x"C0C0BFA4C0A4A492",
-20224 => x"C0C0BFA4C0A4A499",
-20223 => x"C0C0BFA4C0A4A4B0",
-20222 => x"C0C0BFA4C0A4A4A4",
-20221 => x"C0C0BFA4C0A4A4F9",
-20220 => x"C0C0BFA4C0A4A4C0",
-20219 => x"C0C0BFA4C0A4F990",
-20218 => x"C0C0BFA4C0A4F980",
-20217 => x"C0C0BFA4C0A4F9F8",
-20216 => x"C0C0BFA4C0A4F982",
-20215 => x"C0C0BFA4C0A4F992",
-20214 => x"C0C0BFA4C0A4F999",
-20213 => x"C0C0BFA4C0A4F9B0",
-20212 => x"C0C0BFA4C0A4F9A4",
-20211 => x"C0C0BFA4C0A4F9F9",
-20210 => x"C0C0BFA4C0A4F9C0",
-20209 => x"C0C0BFA4C0A4C090",
-20208 => x"C0C0BFA4C0A4C080",
-20207 => x"C0C0BFA4C0A4C0F8",
-20206 => x"C0C0BFA4C0A4C082",
-20205 => x"C0C0BFA4C0A4C092",
-20204 => x"C0C0BFA4C0A4C099",
-20203 => x"C0C0BFA4C0A4C0B0",
-20202 => x"C0C0BFA4C0A4C0A4",
-20201 => x"C0C0BFA4C0A4C0F9",
-20200 => x"C0C0BFA4C0A4C0C0",
-20199 => x"C0C0BFA4C0F99090",
-20198 => x"C0C0BFA4C0F99080",
-20197 => x"C0C0BFA4C0F990F8",
-20196 => x"C0C0BFA4C0F99082",
-20195 => x"C0C0BFA4C0F99092",
-20194 => x"C0C0BFA4C0F99099",
-20193 => x"C0C0BFA4C0F990B0",
-20192 => x"C0C0BFA4C0F990A4",
-20191 => x"C0C0BFA4C0F990F9",
-20190 => x"C0C0BFA4C0F990C0",
-20189 => x"C0C0BFA4C0F98090",
-20188 => x"C0C0BFA4C0F98080",
-20187 => x"C0C0BFA4C0F980F8",
-20186 => x"C0C0BFA4C0F98082",
-20185 => x"C0C0BFA4C0F98092",
-20184 => x"C0C0BFA4C0F98099",
-20183 => x"C0C0BFA4C0F980B0",
-20182 => x"C0C0BFA4C0F980A4",
-20181 => x"C0C0BFA4C0F980F9",
-20180 => x"C0C0BFA4C0F980C0",
-20179 => x"C0C0BFA4C0F9F890",
-20178 => x"C0C0BFA4C0F9F880",
-20177 => x"C0C0BFA4C0F9F8F8",
-20176 => x"C0C0BFA4C0F9F882",
-20175 => x"C0C0BFA4C0F9F892",
-20174 => x"C0C0BFA4C0F9F899",
-20173 => x"C0C0BFA4C0F9F8B0",
-20172 => x"C0C0BFA4C0F9F8A4",
-20171 => x"C0C0BFA4C0F9F8F9",
-20170 => x"C0C0BFA4C0F9F8C0",
-20169 => x"C0C0BFA4C0F98290",
-20168 => x"C0C0BFA4C0F98280",
-20167 => x"C0C0BFA4C0F982F8",
-20166 => x"C0C0BFA4C0F98282",
-20165 => x"C0C0BFA4C0F98292",
-20164 => x"C0C0BFA4C0F98299",
-20163 => x"C0C0BFA4C0F982B0",
-20162 => x"C0C0BFA4C0F982A4",
-20161 => x"C0C0BFA4C0F982F9",
-20160 => x"C0C0BFA4C0F982C0",
-20159 => x"C0C0BFA4C0F99290",
-20158 => x"C0C0BFA4C0F99280",
-20157 => x"C0C0BFA4C0F992F8",
-20156 => x"C0C0BFA4C0F99282",
-20155 => x"C0C0BFA4C0F99292",
-20154 => x"C0C0BFA4C0F99299",
-20153 => x"C0C0BFA4C0F992B0",
-20152 => x"C0C0BFA4C0F992A4",
-20151 => x"C0C0BFA4C0F992F9",
-20150 => x"C0C0BFA4C0F992C0",
-20149 => x"C0C0BFA4C0F99990",
-20148 => x"C0C0BFA4C0F99980",
-20147 => x"C0C0BFA4C0F999F8",
-20146 => x"C0C0BFA4C0F99982",
-20145 => x"C0C0BFA4C0F99992",
-20144 => x"C0C0BFA4C0F99999",
-20143 => x"C0C0BFA4C0F999B0",
-20142 => x"C0C0BFA4C0F999A4",
-20141 => x"C0C0BFA4C0F999F9",
-20140 => x"C0C0BFA4C0F999C0",
-20139 => x"C0C0BFA4C0F9B090",
-20138 => x"C0C0BFA4C0F9B080",
-20137 => x"C0C0BFA4C0F9B0F8",
-20136 => x"C0C0BFA4C0F9B082",
-20135 => x"C0C0BFA4C0F9B092",
-20134 => x"C0C0BFA4C0F9B099",
-20133 => x"C0C0BFA4C0F9B0B0",
-20132 => x"C0C0BFA4C0F9B0A4",
-20131 => x"C0C0BFA4C0F9B0F9",
-20130 => x"C0C0BFA4C0F9B0C0",
-20129 => x"C0C0BFA4C0F9A490",
-20128 => x"C0C0BFA4C0F9A480",
-20127 => x"C0C0BFA4C0F9A4F8",
-20126 => x"C0C0BFA4C0F9A482",
-20125 => x"C0C0BFA4C0F9A492",
-20124 => x"C0C0BFA4C0F9A499",
-20123 => x"C0C0BFA4C0F9A4B0",
-20122 => x"C0C0BFA4C0F9A4A4",
-20121 => x"C0C0BFA4C0F9A4F9",
-20120 => x"C0C0BFA4C0F9A4C0",
-20119 => x"C0C0BFA4C0F9F990",
-20118 => x"C0C0BFA4C0F9F980",
-20117 => x"C0C0BFA4C0F9F9F8",
-20116 => x"C0C0BFA4C0F9F982",
-20115 => x"C0C0BFA4C0F9F992",
-20114 => x"C0C0BFA4C0F9F999",
-20113 => x"C0C0BFA4C0F9F9B0",
-20112 => x"C0C0BFA4C0F9F9A4",
-20111 => x"C0C0BFA4C0F9F9F9",
-20110 => x"C0C0BFA4C0F9F9C0",
-20109 => x"C0C0BFA4C0F9C090",
-20108 => x"C0C0BFA4C0F9C080",
-20107 => x"C0C0BFA4C0F9C0F8",
-20106 => x"C0C0BFA4C0F9C082",
-20105 => x"C0C0BFA4C0F9C092",
-20104 => x"C0C0BFA4C0F9C099",
-20103 => x"C0C0BFA4C0F9C0B0",
-20102 => x"C0C0BFA4C0F9C0A4",
-20101 => x"C0C0BFA4C0F9C0F9",
-20100 => x"C0C0BFA4C0F9C0C0",
-20099 => x"C0C0BFA4C0C09090",
-20098 => x"C0C0BFA4C0C09080",
-20097 => x"C0C0BFA4C0C090F8",
-20096 => x"C0C0BFA4C0C09082",
-20095 => x"C0C0BFA4C0C09092",
-20094 => x"C0C0BFA4C0C09099",
-20093 => x"C0C0BFA4C0C090B0",
-20092 => x"C0C0BFA4C0C090A4",
-20091 => x"C0C0BFA4C0C090F9",
-20090 => x"C0C0BFA4C0C090C0",
-20089 => x"C0C0BFA4C0C08090",
-20088 => x"C0C0BFA4C0C08080",
-20087 => x"C0C0BFA4C0C080F8",
-20086 => x"C0C0BFA4C0C08082",
-20085 => x"C0C0BFA4C0C08092",
-20084 => x"C0C0BFA4C0C08099",
-20083 => x"C0C0BFA4C0C080B0",
-20082 => x"C0C0BFA4C0C080A4",
-20081 => x"C0C0BFA4C0C080F9",
-20080 => x"C0C0BFA4C0C080C0",
-20079 => x"C0C0BFA4C0C0F890",
-20078 => x"C0C0BFA4C0C0F880",
-20077 => x"C0C0BFA4C0C0F8F8",
-20076 => x"C0C0BFA4C0C0F882",
-20075 => x"C0C0BFA4C0C0F892",
-20074 => x"C0C0BFA4C0C0F899",
-20073 => x"C0C0BFA4C0C0F8B0",
-20072 => x"C0C0BFA4C0C0F8A4",
-20071 => x"C0C0BFA4C0C0F8F9",
-20070 => x"C0C0BFA4C0C0F8C0",
-20069 => x"C0C0BFA4C0C08290",
-20068 => x"C0C0BFA4C0C08280",
-20067 => x"C0C0BFA4C0C082F8",
-20066 => x"C0C0BFA4C0C08282",
-20065 => x"C0C0BFA4C0C08292",
-20064 => x"C0C0BFA4C0C08299",
-20063 => x"C0C0BFA4C0C082B0",
-20062 => x"C0C0BFA4C0C082A4",
-20061 => x"C0C0BFA4C0C082F9",
-20060 => x"C0C0BFA4C0C082C0",
-20059 => x"C0C0BFA4C0C09290",
-20058 => x"C0C0BFA4C0C09280",
-20057 => x"C0C0BFA4C0C092F8",
-20056 => x"C0C0BFA4C0C09282",
-20055 => x"C0C0BFA4C0C09292",
-20054 => x"C0C0BFA4C0C09299",
-20053 => x"C0C0BFA4C0C092B0",
-20052 => x"C0C0BFA4C0C092A4",
-20051 => x"C0C0BFA4C0C092F9",
-20050 => x"C0C0BFA4C0C092C0",
-20049 => x"C0C0BFA4C0C09990",
-20048 => x"C0C0BFA4C0C09980",
-20047 => x"C0C0BFA4C0C099F8",
-20046 => x"C0C0BFA4C0C09982",
-20045 => x"C0C0BFA4C0C09992",
-20044 => x"C0C0BFA4C0C09999",
-20043 => x"C0C0BFA4C0C099B0",
-20042 => x"C0C0BFA4C0C099A4",
-20041 => x"C0C0BFA4C0C099F9",
-20040 => x"C0C0BFA4C0C099C0",
-20039 => x"C0C0BFA4C0C0B090",
-20038 => x"C0C0BFA4C0C0B080",
-20037 => x"C0C0BFA4C0C0B0F8",
-20036 => x"C0C0BFA4C0C0B082",
-20035 => x"C0C0BFA4C0C0B092",
-20034 => x"C0C0BFA4C0C0B099",
-20033 => x"C0C0BFA4C0C0B0B0",
-20032 => x"C0C0BFA4C0C0B0A4",
-20031 => x"C0C0BFA4C0C0B0F9",
-20030 => x"C0C0BFA4C0C0B0C0",
-20029 => x"C0C0BFA4C0C0A490",
-20028 => x"C0C0BFA4C0C0A480",
-20027 => x"C0C0BFA4C0C0A4F8",
-20026 => x"C0C0BFA4C0C0A482",
-20025 => x"C0C0BFA4C0C0A492",
-20024 => x"C0C0BFA4C0C0A499",
-20023 => x"C0C0BFA4C0C0A4B0",
-20022 => x"C0C0BFA4C0C0A4A4",
-20021 => x"C0C0BFA4C0C0A4F9",
-20020 => x"C0C0BFA4C0C0A4C0",
-20019 => x"C0C0BFA4C0C0F990",
-20018 => x"C0C0BFA4C0C0F980",
-20017 => x"C0C0BFA4C0C0F9F8",
-20016 => x"C0C0BFA4C0C0F982",
-20015 => x"C0C0BFA4C0C0F992",
-20014 => x"C0C0BFA4C0C0F999",
-20013 => x"C0C0BFA4C0C0F9B0",
-20012 => x"C0C0BFA4C0C0F9A4",
-20011 => x"C0C0BFA4C0C0F9F9",
-20010 => x"C0C0BFA4C0C0F9C0",
-20009 => x"C0C0BFA4C0C0C090",
-20008 => x"C0C0BFA4C0C0C080",
-20007 => x"C0C0BFA4C0C0C0F8",
-20006 => x"C0C0BFA4C0C0C082",
-20005 => x"C0C0BFA4C0C0C092",
-20004 => x"C0C0BFA4C0C0C099",
-20003 => x"C0C0BFA4C0C0C0B0",
-20002 => x"C0C0BFA4C0C0C0A4",
-20001 => x"C0C0BFA4C0C0C0F9",
-20000 => x"C0C0BFA4C0C0C0C0",
-19999 => x"C0C0BFF990909090",
-19998 => x"C0C0BFF990909080",
-19997 => x"C0C0BFF9909090F8",
-19996 => x"C0C0BFF990909082",
-19995 => x"C0C0BFF990909092",
-19994 => x"C0C0BFF990909099",
-19993 => x"C0C0BFF9909090B0",
-19992 => x"C0C0BFF9909090A4",
-19991 => x"C0C0BFF9909090F9",
-19990 => x"C0C0BFF9909090C0",
-19989 => x"C0C0BFF990908090",
-19988 => x"C0C0BFF990908080",
-19987 => x"C0C0BFF9909080F8",
-19986 => x"C0C0BFF990908082",
-19985 => x"C0C0BFF990908092",
-19984 => x"C0C0BFF990908099",
-19983 => x"C0C0BFF9909080B0",
-19982 => x"C0C0BFF9909080A4",
-19981 => x"C0C0BFF9909080F9",
-19980 => x"C0C0BFF9909080C0",
-19979 => x"C0C0BFF99090F890",
-19978 => x"C0C0BFF99090F880",
-19977 => x"C0C0BFF99090F8F8",
-19976 => x"C0C0BFF99090F882",
-19975 => x"C0C0BFF99090F892",
-19974 => x"C0C0BFF99090F899",
-19973 => x"C0C0BFF99090F8B0",
-19972 => x"C0C0BFF99090F8A4",
-19971 => x"C0C0BFF99090F8F9",
-19970 => x"C0C0BFF99090F8C0",
-19969 => x"C0C0BFF990908290",
-19968 => x"C0C0BFF990908280",
-19967 => x"C0C0BFF9909082F8",
-19966 => x"C0C0BFF990908282",
-19965 => x"C0C0BFF990908292",
-19964 => x"C0C0BFF990908299",
-19963 => x"C0C0BFF9909082B0",
-19962 => x"C0C0BFF9909082A4",
-19961 => x"C0C0BFF9909082F9",
-19960 => x"C0C0BFF9909082C0",
-19959 => x"C0C0BFF990909290",
-19958 => x"C0C0BFF990909280",
-19957 => x"C0C0BFF9909092F8",
-19956 => x"C0C0BFF990909282",
-19955 => x"C0C0BFF990909292",
-19954 => x"C0C0BFF990909299",
-19953 => x"C0C0BFF9909092B0",
-19952 => x"C0C0BFF9909092A4",
-19951 => x"C0C0BFF9909092F9",
-19950 => x"C0C0BFF9909092C0",
-19949 => x"C0C0BFF990909990",
-19948 => x"C0C0BFF990909980",
-19947 => x"C0C0BFF9909099F8",
-19946 => x"C0C0BFF990909982",
-19945 => x"C0C0BFF990909992",
-19944 => x"C0C0BFF990909999",
-19943 => x"C0C0BFF9909099B0",
-19942 => x"C0C0BFF9909099A4",
-19941 => x"C0C0BFF9909099F9",
-19940 => x"C0C0BFF9909099C0",
-19939 => x"C0C0BFF99090B090",
-19938 => x"C0C0BFF99090B080",
-19937 => x"C0C0BFF99090B0F8",
-19936 => x"C0C0BFF99090B082",
-19935 => x"C0C0BFF99090B092",
-19934 => x"C0C0BFF99090B099",
-19933 => x"C0C0BFF99090B0B0",
-19932 => x"C0C0BFF99090B0A4",
-19931 => x"C0C0BFF99090B0F9",
-19930 => x"C0C0BFF99090B0C0",
-19929 => x"C0C0BFF99090A490",
-19928 => x"C0C0BFF99090A480",
-19927 => x"C0C0BFF99090A4F8",
-19926 => x"C0C0BFF99090A482",
-19925 => x"C0C0BFF99090A492",
-19924 => x"C0C0BFF99090A499",
-19923 => x"C0C0BFF99090A4B0",
-19922 => x"C0C0BFF99090A4A4",
-19921 => x"C0C0BFF99090A4F9",
-19920 => x"C0C0BFF99090A4C0",
-19919 => x"C0C0BFF99090F990",
-19918 => x"C0C0BFF99090F980",
-19917 => x"C0C0BFF99090F9F8",
-19916 => x"C0C0BFF99090F982",
-19915 => x"C0C0BFF99090F992",
-19914 => x"C0C0BFF99090F999",
-19913 => x"C0C0BFF99090F9B0",
-19912 => x"C0C0BFF99090F9A4",
-19911 => x"C0C0BFF99090F9F9",
-19910 => x"C0C0BFF99090F9C0",
-19909 => x"C0C0BFF99090C090",
-19908 => x"C0C0BFF99090C080",
-19907 => x"C0C0BFF99090C0F8",
-19906 => x"C0C0BFF99090C082",
-19905 => x"C0C0BFF99090C092",
-19904 => x"C0C0BFF99090C099",
-19903 => x"C0C0BFF99090C0B0",
-19902 => x"C0C0BFF99090C0A4",
-19901 => x"C0C0BFF99090C0F9",
-19900 => x"C0C0BFF99090C0C0",
-19899 => x"C0C0BFF990809090",
-19898 => x"C0C0BFF990809080",
-19897 => x"C0C0BFF9908090F8",
-19896 => x"C0C0BFF990809082",
-19895 => x"C0C0BFF990809092",
-19894 => x"C0C0BFF990809099",
-19893 => x"C0C0BFF9908090B0",
-19892 => x"C0C0BFF9908090A4",
-19891 => x"C0C0BFF9908090F9",
-19890 => x"C0C0BFF9908090C0",
-19889 => x"C0C0BFF990808090",
-19888 => x"C0C0BFF990808080",
-19887 => x"C0C0BFF9908080F8",
-19886 => x"C0C0BFF990808082",
-19885 => x"C0C0BFF990808092",
-19884 => x"C0C0BFF990808099",
-19883 => x"C0C0BFF9908080B0",
-19882 => x"C0C0BFF9908080A4",
-19881 => x"C0C0BFF9908080F9",
-19880 => x"C0C0BFF9908080C0",
-19879 => x"C0C0BFF99080F890",
-19878 => x"C0C0BFF99080F880",
-19877 => x"C0C0BFF99080F8F8",
-19876 => x"C0C0BFF99080F882",
-19875 => x"C0C0BFF99080F892",
-19874 => x"C0C0BFF99080F899",
-19873 => x"C0C0BFF99080F8B0",
-19872 => x"C0C0BFF99080F8A4",
-19871 => x"C0C0BFF99080F8F9",
-19870 => x"C0C0BFF99080F8C0",
-19869 => x"C0C0BFF990808290",
-19868 => x"C0C0BFF990808280",
-19867 => x"C0C0BFF9908082F8",
-19866 => x"C0C0BFF990808282",
-19865 => x"C0C0BFF990808292",
-19864 => x"C0C0BFF990808299",
-19863 => x"C0C0BFF9908082B0",
-19862 => x"C0C0BFF9908082A4",
-19861 => x"C0C0BFF9908082F9",
-19860 => x"C0C0BFF9908082C0",
-19859 => x"C0C0BFF990809290",
-19858 => x"C0C0BFF990809280",
-19857 => x"C0C0BFF9908092F8",
-19856 => x"C0C0BFF990809282",
-19855 => x"C0C0BFF990809292",
-19854 => x"C0C0BFF990809299",
-19853 => x"C0C0BFF9908092B0",
-19852 => x"C0C0BFF9908092A4",
-19851 => x"C0C0BFF9908092F9",
-19850 => x"C0C0BFF9908092C0",
-19849 => x"C0C0BFF990809990",
-19848 => x"C0C0BFF990809980",
-19847 => x"C0C0BFF9908099F8",
-19846 => x"C0C0BFF990809982",
-19845 => x"C0C0BFF990809992",
-19844 => x"C0C0BFF990809999",
-19843 => x"C0C0BFF9908099B0",
-19842 => x"C0C0BFF9908099A4",
-19841 => x"C0C0BFF9908099F9",
-19840 => x"C0C0BFF9908099C0",
-19839 => x"C0C0BFF99080B090",
-19838 => x"C0C0BFF99080B080",
-19837 => x"C0C0BFF99080B0F8",
-19836 => x"C0C0BFF99080B082",
-19835 => x"C0C0BFF99080B092",
-19834 => x"C0C0BFF99080B099",
-19833 => x"C0C0BFF99080B0B0",
-19832 => x"C0C0BFF99080B0A4",
-19831 => x"C0C0BFF99080B0F9",
-19830 => x"C0C0BFF99080B0C0",
-19829 => x"C0C0BFF99080A490",
-19828 => x"C0C0BFF99080A480",
-19827 => x"C0C0BFF99080A4F8",
-19826 => x"C0C0BFF99080A482",
-19825 => x"C0C0BFF99080A492",
-19824 => x"C0C0BFF99080A499",
-19823 => x"C0C0BFF99080A4B0",
-19822 => x"C0C0BFF99080A4A4",
-19821 => x"C0C0BFF99080A4F9",
-19820 => x"C0C0BFF99080A4C0",
-19819 => x"C0C0BFF99080F990",
-19818 => x"C0C0BFF99080F980",
-19817 => x"C0C0BFF99080F9F8",
-19816 => x"C0C0BFF99080F982",
-19815 => x"C0C0BFF99080F992",
-19814 => x"C0C0BFF99080F999",
-19813 => x"C0C0BFF99080F9B0",
-19812 => x"C0C0BFF99080F9A4",
-19811 => x"C0C0BFF99080F9F9",
-19810 => x"C0C0BFF99080F9C0",
-19809 => x"C0C0BFF99080C090",
-19808 => x"C0C0BFF99080C080",
-19807 => x"C0C0BFF99080C0F8",
-19806 => x"C0C0BFF99080C082",
-19805 => x"C0C0BFF99080C092",
-19804 => x"C0C0BFF99080C099",
-19803 => x"C0C0BFF99080C0B0",
-19802 => x"C0C0BFF99080C0A4",
-19801 => x"C0C0BFF99080C0F9",
-19800 => x"C0C0BFF99080C0C0",
-19799 => x"C0C0BFF990F89090",
-19798 => x"C0C0BFF990F89080",
-19797 => x"C0C0BFF990F890F8",
-19796 => x"C0C0BFF990F89082",
-19795 => x"C0C0BFF990F89092",
-19794 => x"C0C0BFF990F89099",
-19793 => x"C0C0BFF990F890B0",
-19792 => x"C0C0BFF990F890A4",
-19791 => x"C0C0BFF990F890F9",
-19790 => x"C0C0BFF990F890C0",
-19789 => x"C0C0BFF990F88090",
-19788 => x"C0C0BFF990F88080",
-19787 => x"C0C0BFF990F880F8",
-19786 => x"C0C0BFF990F88082",
-19785 => x"C0C0BFF990F88092",
-19784 => x"C0C0BFF990F88099",
-19783 => x"C0C0BFF990F880B0",
-19782 => x"C0C0BFF990F880A4",
-19781 => x"C0C0BFF990F880F9",
-19780 => x"C0C0BFF990F880C0",
-19779 => x"C0C0BFF990F8F890",
-19778 => x"C0C0BFF990F8F880",
-19777 => x"C0C0BFF990F8F8F8",
-19776 => x"C0C0BFF990F8F882",
-19775 => x"C0C0BFF990F8F892",
-19774 => x"C0C0BFF990F8F899",
-19773 => x"C0C0BFF990F8F8B0",
-19772 => x"C0C0BFF990F8F8A4",
-19771 => x"C0C0BFF990F8F8F9",
-19770 => x"C0C0BFF990F8F8C0",
-19769 => x"C0C0BFF990F88290",
-19768 => x"C0C0BFF990F88280",
-19767 => x"C0C0BFF990F882F8",
-19766 => x"C0C0BFF990F88282",
-19765 => x"C0C0BFF990F88292",
-19764 => x"C0C0BFF990F88299",
-19763 => x"C0C0BFF990F882B0",
-19762 => x"C0C0BFF990F882A4",
-19761 => x"C0C0BFF990F882F9",
-19760 => x"C0C0BFF990F882C0",
-19759 => x"C0C0BFF990F89290",
-19758 => x"C0C0BFF990F89280",
-19757 => x"C0C0BFF990F892F8",
-19756 => x"C0C0BFF990F89282",
-19755 => x"C0C0BFF990F89292",
-19754 => x"C0C0BFF990F89299",
-19753 => x"C0C0BFF990F892B0",
-19752 => x"C0C0BFF990F892A4",
-19751 => x"C0C0BFF990F892F9",
-19750 => x"C0C0BFF990F892C0",
-19749 => x"C0C0BFF990F89990",
-19748 => x"C0C0BFF990F89980",
-19747 => x"C0C0BFF990F899F8",
-19746 => x"C0C0BFF990F89982",
-19745 => x"C0C0BFF990F89992",
-19744 => x"C0C0BFF990F89999",
-19743 => x"C0C0BFF990F899B0",
-19742 => x"C0C0BFF990F899A4",
-19741 => x"C0C0BFF990F899F9",
-19740 => x"C0C0BFF990F899C0",
-19739 => x"C0C0BFF990F8B090",
-19738 => x"C0C0BFF990F8B080",
-19737 => x"C0C0BFF990F8B0F8",
-19736 => x"C0C0BFF990F8B082",
-19735 => x"C0C0BFF990F8B092",
-19734 => x"C0C0BFF990F8B099",
-19733 => x"C0C0BFF990F8B0B0",
-19732 => x"C0C0BFF990F8B0A4",
-19731 => x"C0C0BFF990F8B0F9",
-19730 => x"C0C0BFF990F8B0C0",
-19729 => x"C0C0BFF990F8A490",
-19728 => x"C0C0BFF990F8A480",
-19727 => x"C0C0BFF990F8A4F8",
-19726 => x"C0C0BFF990F8A482",
-19725 => x"C0C0BFF990F8A492",
-19724 => x"C0C0BFF990F8A499",
-19723 => x"C0C0BFF990F8A4B0",
-19722 => x"C0C0BFF990F8A4A4",
-19721 => x"C0C0BFF990F8A4F9",
-19720 => x"C0C0BFF990F8A4C0",
-19719 => x"C0C0BFF990F8F990",
-19718 => x"C0C0BFF990F8F980",
-19717 => x"C0C0BFF990F8F9F8",
-19716 => x"C0C0BFF990F8F982",
-19715 => x"C0C0BFF990F8F992",
-19714 => x"C0C0BFF990F8F999",
-19713 => x"C0C0BFF990F8F9B0",
-19712 => x"C0C0BFF990F8F9A4",
-19711 => x"C0C0BFF990F8F9F9",
-19710 => x"C0C0BFF990F8F9C0",
-19709 => x"C0C0BFF990F8C090",
-19708 => x"C0C0BFF990F8C080",
-19707 => x"C0C0BFF990F8C0F8",
-19706 => x"C0C0BFF990F8C082",
-19705 => x"C0C0BFF990F8C092",
-19704 => x"C0C0BFF990F8C099",
-19703 => x"C0C0BFF990F8C0B0",
-19702 => x"C0C0BFF990F8C0A4",
-19701 => x"C0C0BFF990F8C0F9",
-19700 => x"C0C0BFF990F8C0C0",
-19699 => x"C0C0BFF990829090",
-19698 => x"C0C0BFF990829080",
-19697 => x"C0C0BFF9908290F8",
-19696 => x"C0C0BFF990829082",
-19695 => x"C0C0BFF990829092",
-19694 => x"C0C0BFF990829099",
-19693 => x"C0C0BFF9908290B0",
-19692 => x"C0C0BFF9908290A4",
-19691 => x"C0C0BFF9908290F9",
-19690 => x"C0C0BFF9908290C0",
-19689 => x"C0C0BFF990828090",
-19688 => x"C0C0BFF990828080",
-19687 => x"C0C0BFF9908280F8",
-19686 => x"C0C0BFF990828082",
-19685 => x"C0C0BFF990828092",
-19684 => x"C0C0BFF990828099",
-19683 => x"C0C0BFF9908280B0",
-19682 => x"C0C0BFF9908280A4",
-19681 => x"C0C0BFF9908280F9",
-19680 => x"C0C0BFF9908280C0",
-19679 => x"C0C0BFF99082F890",
-19678 => x"C0C0BFF99082F880",
-19677 => x"C0C0BFF99082F8F8",
-19676 => x"C0C0BFF99082F882",
-19675 => x"C0C0BFF99082F892",
-19674 => x"C0C0BFF99082F899",
-19673 => x"C0C0BFF99082F8B0",
-19672 => x"C0C0BFF99082F8A4",
-19671 => x"C0C0BFF99082F8F9",
-19670 => x"C0C0BFF99082F8C0",
-19669 => x"C0C0BFF990828290",
-19668 => x"C0C0BFF990828280",
-19667 => x"C0C0BFF9908282F8",
-19666 => x"C0C0BFF990828282",
-19665 => x"C0C0BFF990828292",
-19664 => x"C0C0BFF990828299",
-19663 => x"C0C0BFF9908282B0",
-19662 => x"C0C0BFF9908282A4",
-19661 => x"C0C0BFF9908282F9",
-19660 => x"C0C0BFF9908282C0",
-19659 => x"C0C0BFF990829290",
-19658 => x"C0C0BFF990829280",
-19657 => x"C0C0BFF9908292F8",
-19656 => x"C0C0BFF990829282",
-19655 => x"C0C0BFF990829292",
-19654 => x"C0C0BFF990829299",
-19653 => x"C0C0BFF9908292B0",
-19652 => x"C0C0BFF9908292A4",
-19651 => x"C0C0BFF9908292F9",
-19650 => x"C0C0BFF9908292C0",
-19649 => x"C0C0BFF990829990",
-19648 => x"C0C0BFF990829980",
-19647 => x"C0C0BFF9908299F8",
-19646 => x"C0C0BFF990829982",
-19645 => x"C0C0BFF990829992",
-19644 => x"C0C0BFF990829999",
-19643 => x"C0C0BFF9908299B0",
-19642 => x"C0C0BFF9908299A4",
-19641 => x"C0C0BFF9908299F9",
-19640 => x"C0C0BFF9908299C0",
-19639 => x"C0C0BFF99082B090",
-19638 => x"C0C0BFF99082B080",
-19637 => x"C0C0BFF99082B0F8",
-19636 => x"C0C0BFF99082B082",
-19635 => x"C0C0BFF99082B092",
-19634 => x"C0C0BFF99082B099",
-19633 => x"C0C0BFF99082B0B0",
-19632 => x"C0C0BFF99082B0A4",
-19631 => x"C0C0BFF99082B0F9",
-19630 => x"C0C0BFF99082B0C0",
-19629 => x"C0C0BFF99082A490",
-19628 => x"C0C0BFF99082A480",
-19627 => x"C0C0BFF99082A4F8",
-19626 => x"C0C0BFF99082A482",
-19625 => x"C0C0BFF99082A492",
-19624 => x"C0C0BFF99082A499",
-19623 => x"C0C0BFF99082A4B0",
-19622 => x"C0C0BFF99082A4A4",
-19621 => x"C0C0BFF99082A4F9",
-19620 => x"C0C0BFF99082A4C0",
-19619 => x"C0C0BFF99082F990",
-19618 => x"C0C0BFF99082F980",
-19617 => x"C0C0BFF99082F9F8",
-19616 => x"C0C0BFF99082F982",
-19615 => x"C0C0BFF99082F992",
-19614 => x"C0C0BFF99082F999",
-19613 => x"C0C0BFF99082F9B0",
-19612 => x"C0C0BFF99082F9A4",
-19611 => x"C0C0BFF99082F9F9",
-19610 => x"C0C0BFF99082F9C0",
-19609 => x"C0C0BFF99082C090",
-19608 => x"C0C0BFF99082C080",
-19607 => x"C0C0BFF99082C0F8",
-19606 => x"C0C0BFF99082C082",
-19605 => x"C0C0BFF99082C092",
-19604 => x"C0C0BFF99082C099",
-19603 => x"C0C0BFF99082C0B0",
-19602 => x"C0C0BFF99082C0A4",
-19601 => x"C0C0BFF99082C0F9",
-19600 => x"C0C0BFF99082C0C0",
-19599 => x"C0C0BFF990929090",
-19598 => x"C0C0BFF990929080",
-19597 => x"C0C0BFF9909290F8",
-19596 => x"C0C0BFF990929082",
-19595 => x"C0C0BFF990929092",
-19594 => x"C0C0BFF990929099",
-19593 => x"C0C0BFF9909290B0",
-19592 => x"C0C0BFF9909290A4",
-19591 => x"C0C0BFF9909290F9",
-19590 => x"C0C0BFF9909290C0",
-19589 => x"C0C0BFF990928090",
-19588 => x"C0C0BFF990928080",
-19587 => x"C0C0BFF9909280F8",
-19586 => x"C0C0BFF990928082",
-19585 => x"C0C0BFF990928092",
-19584 => x"C0C0BFF990928099",
-19583 => x"C0C0BFF9909280B0",
-19582 => x"C0C0BFF9909280A4",
-19581 => x"C0C0BFF9909280F9",
-19580 => x"C0C0BFF9909280C0",
-19579 => x"C0C0BFF99092F890",
-19578 => x"C0C0BFF99092F880",
-19577 => x"C0C0BFF99092F8F8",
-19576 => x"C0C0BFF99092F882",
-19575 => x"C0C0BFF99092F892",
-19574 => x"C0C0BFF99092F899",
-19573 => x"C0C0BFF99092F8B0",
-19572 => x"C0C0BFF99092F8A4",
-19571 => x"C0C0BFF99092F8F9",
-19570 => x"C0C0BFF99092F8C0",
-19569 => x"C0C0BFF990928290",
-19568 => x"C0C0BFF990928280",
-19567 => x"C0C0BFF9909282F8",
-19566 => x"C0C0BFF990928282",
-19565 => x"C0C0BFF990928292",
-19564 => x"C0C0BFF990928299",
-19563 => x"C0C0BFF9909282B0",
-19562 => x"C0C0BFF9909282A4",
-19561 => x"C0C0BFF9909282F9",
-19560 => x"C0C0BFF9909282C0",
-19559 => x"C0C0BFF990929290",
-19558 => x"C0C0BFF990929280",
-19557 => x"C0C0BFF9909292F8",
-19556 => x"C0C0BFF990929282",
-19555 => x"C0C0BFF990929292",
-19554 => x"C0C0BFF990929299",
-19553 => x"C0C0BFF9909292B0",
-19552 => x"C0C0BFF9909292A4",
-19551 => x"C0C0BFF9909292F9",
-19550 => x"C0C0BFF9909292C0",
-19549 => x"C0C0BFF990929990",
-19548 => x"C0C0BFF990929980",
-19547 => x"C0C0BFF9909299F8",
-19546 => x"C0C0BFF990929982",
-19545 => x"C0C0BFF990929992",
-19544 => x"C0C0BFF990929999",
-19543 => x"C0C0BFF9909299B0",
-19542 => x"C0C0BFF9909299A4",
-19541 => x"C0C0BFF9909299F9",
-19540 => x"C0C0BFF9909299C0",
-19539 => x"C0C0BFF99092B090",
-19538 => x"C0C0BFF99092B080",
-19537 => x"C0C0BFF99092B0F8",
-19536 => x"C0C0BFF99092B082",
-19535 => x"C0C0BFF99092B092",
-19534 => x"C0C0BFF99092B099",
-19533 => x"C0C0BFF99092B0B0",
-19532 => x"C0C0BFF99092B0A4",
-19531 => x"C0C0BFF99092B0F9",
-19530 => x"C0C0BFF99092B0C0",
-19529 => x"C0C0BFF99092A490",
-19528 => x"C0C0BFF99092A480",
-19527 => x"C0C0BFF99092A4F8",
-19526 => x"C0C0BFF99092A482",
-19525 => x"C0C0BFF99092A492",
-19524 => x"C0C0BFF99092A499",
-19523 => x"C0C0BFF99092A4B0",
-19522 => x"C0C0BFF99092A4A4",
-19521 => x"C0C0BFF99092A4F9",
-19520 => x"C0C0BFF99092A4C0",
-19519 => x"C0C0BFF99092F990",
-19518 => x"C0C0BFF99092F980",
-19517 => x"C0C0BFF99092F9F8",
-19516 => x"C0C0BFF99092F982",
-19515 => x"C0C0BFF99092F992",
-19514 => x"C0C0BFF99092F999",
-19513 => x"C0C0BFF99092F9B0",
-19512 => x"C0C0BFF99092F9A4",
-19511 => x"C0C0BFF99092F9F9",
-19510 => x"C0C0BFF99092F9C0",
-19509 => x"C0C0BFF99092C090",
-19508 => x"C0C0BFF99092C080",
-19507 => x"C0C0BFF99092C0F8",
-19506 => x"C0C0BFF99092C082",
-19505 => x"C0C0BFF99092C092",
-19504 => x"C0C0BFF99092C099",
-19503 => x"C0C0BFF99092C0B0",
-19502 => x"C0C0BFF99092C0A4",
-19501 => x"C0C0BFF99092C0F9",
-19500 => x"C0C0BFF99092C0C0",
-19499 => x"C0C0BFF990999090",
-19498 => x"C0C0BFF990999080",
-19497 => x"C0C0BFF9909990F8",
-19496 => x"C0C0BFF990999082",
-19495 => x"C0C0BFF990999092",
-19494 => x"C0C0BFF990999099",
-19493 => x"C0C0BFF9909990B0",
-19492 => x"C0C0BFF9909990A4",
-19491 => x"C0C0BFF9909990F9",
-19490 => x"C0C0BFF9909990C0",
-19489 => x"C0C0BFF990998090",
-19488 => x"C0C0BFF990998080",
-19487 => x"C0C0BFF9909980F8",
-19486 => x"C0C0BFF990998082",
-19485 => x"C0C0BFF990998092",
-19484 => x"C0C0BFF990998099",
-19483 => x"C0C0BFF9909980B0",
-19482 => x"C0C0BFF9909980A4",
-19481 => x"C0C0BFF9909980F9",
-19480 => x"C0C0BFF9909980C0",
-19479 => x"C0C0BFF99099F890",
-19478 => x"C0C0BFF99099F880",
-19477 => x"C0C0BFF99099F8F8",
-19476 => x"C0C0BFF99099F882",
-19475 => x"C0C0BFF99099F892",
-19474 => x"C0C0BFF99099F899",
-19473 => x"C0C0BFF99099F8B0",
-19472 => x"C0C0BFF99099F8A4",
-19471 => x"C0C0BFF99099F8F9",
-19470 => x"C0C0BFF99099F8C0",
-19469 => x"C0C0BFF990998290",
-19468 => x"C0C0BFF990998280",
-19467 => x"C0C0BFF9909982F8",
-19466 => x"C0C0BFF990998282",
-19465 => x"C0C0BFF990998292",
-19464 => x"C0C0BFF990998299",
-19463 => x"C0C0BFF9909982B0",
-19462 => x"C0C0BFF9909982A4",
-19461 => x"C0C0BFF9909982F9",
-19460 => x"C0C0BFF9909982C0",
-19459 => x"C0C0BFF990999290",
-19458 => x"C0C0BFF990999280",
-19457 => x"C0C0BFF9909992F8",
-19456 => x"C0C0BFF990999282",
-19455 => x"C0C0BFF990999292",
-19454 => x"C0C0BFF990999299",
-19453 => x"C0C0BFF9909992B0",
-19452 => x"C0C0BFF9909992A4",
-19451 => x"C0C0BFF9909992F9",
-19450 => x"C0C0BFF9909992C0",
-19449 => x"C0C0BFF990999990",
-19448 => x"C0C0BFF990999980",
-19447 => x"C0C0BFF9909999F8",
-19446 => x"C0C0BFF990999982",
-19445 => x"C0C0BFF990999992",
-19444 => x"C0C0BFF990999999",
-19443 => x"C0C0BFF9909999B0",
-19442 => x"C0C0BFF9909999A4",
-19441 => x"C0C0BFF9909999F9",
-19440 => x"C0C0BFF9909999C0",
-19439 => x"C0C0BFF99099B090",
-19438 => x"C0C0BFF99099B080",
-19437 => x"C0C0BFF99099B0F8",
-19436 => x"C0C0BFF99099B082",
-19435 => x"C0C0BFF99099B092",
-19434 => x"C0C0BFF99099B099",
-19433 => x"C0C0BFF99099B0B0",
-19432 => x"C0C0BFF99099B0A4",
-19431 => x"C0C0BFF99099B0F9",
-19430 => x"C0C0BFF99099B0C0",
-19429 => x"C0C0BFF99099A490",
-19428 => x"C0C0BFF99099A480",
-19427 => x"C0C0BFF99099A4F8",
-19426 => x"C0C0BFF99099A482",
-19425 => x"C0C0BFF99099A492",
-19424 => x"C0C0BFF99099A499",
-19423 => x"C0C0BFF99099A4B0",
-19422 => x"C0C0BFF99099A4A4",
-19421 => x"C0C0BFF99099A4F9",
-19420 => x"C0C0BFF99099A4C0",
-19419 => x"C0C0BFF99099F990",
-19418 => x"C0C0BFF99099F980",
-19417 => x"C0C0BFF99099F9F8",
-19416 => x"C0C0BFF99099F982",
-19415 => x"C0C0BFF99099F992",
-19414 => x"C0C0BFF99099F999",
-19413 => x"C0C0BFF99099F9B0",
-19412 => x"C0C0BFF99099F9A4",
-19411 => x"C0C0BFF99099F9F9",
-19410 => x"C0C0BFF99099F9C0",
-19409 => x"C0C0BFF99099C090",
-19408 => x"C0C0BFF99099C080",
-19407 => x"C0C0BFF99099C0F8",
-19406 => x"C0C0BFF99099C082",
-19405 => x"C0C0BFF99099C092",
-19404 => x"C0C0BFF99099C099",
-19403 => x"C0C0BFF99099C0B0",
-19402 => x"C0C0BFF99099C0A4",
-19401 => x"C0C0BFF99099C0F9",
-19400 => x"C0C0BFF99099C0C0",
-19399 => x"C0C0BFF990B09090",
-19398 => x"C0C0BFF990B09080",
-19397 => x"C0C0BFF990B090F8",
-19396 => x"C0C0BFF990B09082",
-19395 => x"C0C0BFF990B09092",
-19394 => x"C0C0BFF990B09099",
-19393 => x"C0C0BFF990B090B0",
-19392 => x"C0C0BFF990B090A4",
-19391 => x"C0C0BFF990B090F9",
-19390 => x"C0C0BFF990B090C0",
-19389 => x"C0C0BFF990B08090",
-19388 => x"C0C0BFF990B08080",
-19387 => x"C0C0BFF990B080F8",
-19386 => x"C0C0BFF990B08082",
-19385 => x"C0C0BFF990B08092",
-19384 => x"C0C0BFF990B08099",
-19383 => x"C0C0BFF990B080B0",
-19382 => x"C0C0BFF990B080A4",
-19381 => x"C0C0BFF990B080F9",
-19380 => x"C0C0BFF990B080C0",
-19379 => x"C0C0BFF990B0F890",
-19378 => x"C0C0BFF990B0F880",
-19377 => x"C0C0BFF990B0F8F8",
-19376 => x"C0C0BFF990B0F882",
-19375 => x"C0C0BFF990B0F892",
-19374 => x"C0C0BFF990B0F899",
-19373 => x"C0C0BFF990B0F8B0",
-19372 => x"C0C0BFF990B0F8A4",
-19371 => x"C0C0BFF990B0F8F9",
-19370 => x"C0C0BFF990B0F8C0",
-19369 => x"C0C0BFF990B08290",
-19368 => x"C0C0BFF990B08280",
-19367 => x"C0C0BFF990B082F8",
-19366 => x"C0C0BFF990B08282",
-19365 => x"C0C0BFF990B08292",
-19364 => x"C0C0BFF990B08299",
-19363 => x"C0C0BFF990B082B0",
-19362 => x"C0C0BFF990B082A4",
-19361 => x"C0C0BFF990B082F9",
-19360 => x"C0C0BFF990B082C0",
-19359 => x"C0C0BFF990B09290",
-19358 => x"C0C0BFF990B09280",
-19357 => x"C0C0BFF990B092F8",
-19356 => x"C0C0BFF990B09282",
-19355 => x"C0C0BFF990B09292",
-19354 => x"C0C0BFF990B09299",
-19353 => x"C0C0BFF990B092B0",
-19352 => x"C0C0BFF990B092A4",
-19351 => x"C0C0BFF990B092F9",
-19350 => x"C0C0BFF990B092C0",
-19349 => x"C0C0BFF990B09990",
-19348 => x"C0C0BFF990B09980",
-19347 => x"C0C0BFF990B099F8",
-19346 => x"C0C0BFF990B09982",
-19345 => x"C0C0BFF990B09992",
-19344 => x"C0C0BFF990B09999",
-19343 => x"C0C0BFF990B099B0",
-19342 => x"C0C0BFF990B099A4",
-19341 => x"C0C0BFF990B099F9",
-19340 => x"C0C0BFF990B099C0",
-19339 => x"C0C0BFF990B0B090",
-19338 => x"C0C0BFF990B0B080",
-19337 => x"C0C0BFF990B0B0F8",
-19336 => x"C0C0BFF990B0B082",
-19335 => x"C0C0BFF990B0B092",
-19334 => x"C0C0BFF990B0B099",
-19333 => x"C0C0BFF990B0B0B0",
-19332 => x"C0C0BFF990B0B0A4",
-19331 => x"C0C0BFF990B0B0F9",
-19330 => x"C0C0BFF990B0B0C0",
-19329 => x"C0C0BFF990B0A490",
-19328 => x"C0C0BFF990B0A480",
-19327 => x"C0C0BFF990B0A4F8",
-19326 => x"C0C0BFF990B0A482",
-19325 => x"C0C0BFF990B0A492",
-19324 => x"C0C0BFF990B0A499",
-19323 => x"C0C0BFF990B0A4B0",
-19322 => x"C0C0BFF990B0A4A4",
-19321 => x"C0C0BFF990B0A4F9",
-19320 => x"C0C0BFF990B0A4C0",
-19319 => x"C0C0BFF990B0F990",
-19318 => x"C0C0BFF990B0F980",
-19317 => x"C0C0BFF990B0F9F8",
-19316 => x"C0C0BFF990B0F982",
-19315 => x"C0C0BFF990B0F992",
-19314 => x"C0C0BFF990B0F999",
-19313 => x"C0C0BFF990B0F9B0",
-19312 => x"C0C0BFF990B0F9A4",
-19311 => x"C0C0BFF990B0F9F9",
-19310 => x"C0C0BFF990B0F9C0",
-19309 => x"C0C0BFF990B0C090",
-19308 => x"C0C0BFF990B0C080",
-19307 => x"C0C0BFF990B0C0F8",
-19306 => x"C0C0BFF990B0C082",
-19305 => x"C0C0BFF990B0C092",
-19304 => x"C0C0BFF990B0C099",
-19303 => x"C0C0BFF990B0C0B0",
-19302 => x"C0C0BFF990B0C0A4",
-19301 => x"C0C0BFF990B0C0F9",
-19300 => x"C0C0BFF990B0C0C0",
-19299 => x"C0C0BFF990A49090",
-19298 => x"C0C0BFF990A49080",
-19297 => x"C0C0BFF990A490F8",
-19296 => x"C0C0BFF990A49082",
-19295 => x"C0C0BFF990A49092",
-19294 => x"C0C0BFF990A49099",
-19293 => x"C0C0BFF990A490B0",
-19292 => x"C0C0BFF990A490A4",
-19291 => x"C0C0BFF990A490F9",
-19290 => x"C0C0BFF990A490C0",
-19289 => x"C0C0BFF990A48090",
-19288 => x"C0C0BFF990A48080",
-19287 => x"C0C0BFF990A480F8",
-19286 => x"C0C0BFF990A48082",
-19285 => x"C0C0BFF990A48092",
-19284 => x"C0C0BFF990A48099",
-19283 => x"C0C0BFF990A480B0",
-19282 => x"C0C0BFF990A480A4",
-19281 => x"C0C0BFF990A480F9",
-19280 => x"C0C0BFF990A480C0",
-19279 => x"C0C0BFF990A4F890",
-19278 => x"C0C0BFF990A4F880",
-19277 => x"C0C0BFF990A4F8F8",
-19276 => x"C0C0BFF990A4F882",
-19275 => x"C0C0BFF990A4F892",
-19274 => x"C0C0BFF990A4F899",
-19273 => x"C0C0BFF990A4F8B0",
-19272 => x"C0C0BFF990A4F8A4",
-19271 => x"C0C0BFF990A4F8F9",
-19270 => x"C0C0BFF990A4F8C0",
-19269 => x"C0C0BFF990A48290",
-19268 => x"C0C0BFF990A48280",
-19267 => x"C0C0BFF990A482F8",
-19266 => x"C0C0BFF990A48282",
-19265 => x"C0C0BFF990A48292",
-19264 => x"C0C0BFF990A48299",
-19263 => x"C0C0BFF990A482B0",
-19262 => x"C0C0BFF990A482A4",
-19261 => x"C0C0BFF990A482F9",
-19260 => x"C0C0BFF990A482C0",
-19259 => x"C0C0BFF990A49290",
-19258 => x"C0C0BFF990A49280",
-19257 => x"C0C0BFF990A492F8",
-19256 => x"C0C0BFF990A49282",
-19255 => x"C0C0BFF990A49292",
-19254 => x"C0C0BFF990A49299",
-19253 => x"C0C0BFF990A492B0",
-19252 => x"C0C0BFF990A492A4",
-19251 => x"C0C0BFF990A492F9",
-19250 => x"C0C0BFF990A492C0",
-19249 => x"C0C0BFF990A49990",
-19248 => x"C0C0BFF990A49980",
-19247 => x"C0C0BFF990A499F8",
-19246 => x"C0C0BFF990A49982",
-19245 => x"C0C0BFF990A49992",
-19244 => x"C0C0BFF990A49999",
-19243 => x"C0C0BFF990A499B0",
-19242 => x"C0C0BFF990A499A4",
-19241 => x"C0C0BFF990A499F9",
-19240 => x"C0C0BFF990A499C0",
-19239 => x"C0C0BFF990A4B090",
-19238 => x"C0C0BFF990A4B080",
-19237 => x"C0C0BFF990A4B0F8",
-19236 => x"C0C0BFF990A4B082",
-19235 => x"C0C0BFF990A4B092",
-19234 => x"C0C0BFF990A4B099",
-19233 => x"C0C0BFF990A4B0B0",
-19232 => x"C0C0BFF990A4B0A4",
-19231 => x"C0C0BFF990A4B0F9",
-19230 => x"C0C0BFF990A4B0C0",
-19229 => x"C0C0BFF990A4A490",
-19228 => x"C0C0BFF990A4A480",
-19227 => x"C0C0BFF990A4A4F8",
-19226 => x"C0C0BFF990A4A482",
-19225 => x"C0C0BFF990A4A492",
-19224 => x"C0C0BFF990A4A499",
-19223 => x"C0C0BFF990A4A4B0",
-19222 => x"C0C0BFF990A4A4A4",
-19221 => x"C0C0BFF990A4A4F9",
-19220 => x"C0C0BFF990A4A4C0",
-19219 => x"C0C0BFF990A4F990",
-19218 => x"C0C0BFF990A4F980",
-19217 => x"C0C0BFF990A4F9F8",
-19216 => x"C0C0BFF990A4F982",
-19215 => x"C0C0BFF990A4F992",
-19214 => x"C0C0BFF990A4F999",
-19213 => x"C0C0BFF990A4F9B0",
-19212 => x"C0C0BFF990A4F9A4",
-19211 => x"C0C0BFF990A4F9F9",
-19210 => x"C0C0BFF990A4F9C0",
-19209 => x"C0C0BFF990A4C090",
-19208 => x"C0C0BFF990A4C080",
-19207 => x"C0C0BFF990A4C0F8",
-19206 => x"C0C0BFF990A4C082",
-19205 => x"C0C0BFF990A4C092",
-19204 => x"C0C0BFF990A4C099",
-19203 => x"C0C0BFF990A4C0B0",
-19202 => x"C0C0BFF990A4C0A4",
-19201 => x"C0C0BFF990A4C0F9",
-19200 => x"C0C0BFF990A4C0C0",
-19199 => x"C0C0BFF990F99090",
-19198 => x"C0C0BFF990F99080",
-19197 => x"C0C0BFF990F990F8",
-19196 => x"C0C0BFF990F99082",
-19195 => x"C0C0BFF990F99092",
-19194 => x"C0C0BFF990F99099",
-19193 => x"C0C0BFF990F990B0",
-19192 => x"C0C0BFF990F990A4",
-19191 => x"C0C0BFF990F990F9",
-19190 => x"C0C0BFF990F990C0",
-19189 => x"C0C0BFF990F98090",
-19188 => x"C0C0BFF990F98080",
-19187 => x"C0C0BFF990F980F8",
-19186 => x"C0C0BFF990F98082",
-19185 => x"C0C0BFF990F98092",
-19184 => x"C0C0BFF990F98099",
-19183 => x"C0C0BFF990F980B0",
-19182 => x"C0C0BFF990F980A4",
-19181 => x"C0C0BFF990F980F9",
-19180 => x"C0C0BFF990F980C0",
-19179 => x"C0C0BFF990F9F890",
-19178 => x"C0C0BFF990F9F880",
-19177 => x"C0C0BFF990F9F8F8",
-19176 => x"C0C0BFF990F9F882",
-19175 => x"C0C0BFF990F9F892",
-19174 => x"C0C0BFF990F9F899",
-19173 => x"C0C0BFF990F9F8B0",
-19172 => x"C0C0BFF990F9F8A4",
-19171 => x"C0C0BFF990F9F8F9",
-19170 => x"C0C0BFF990F9F8C0",
-19169 => x"C0C0BFF990F98290",
-19168 => x"C0C0BFF990F98280",
-19167 => x"C0C0BFF990F982F8",
-19166 => x"C0C0BFF990F98282",
-19165 => x"C0C0BFF990F98292",
-19164 => x"C0C0BFF990F98299",
-19163 => x"C0C0BFF990F982B0",
-19162 => x"C0C0BFF990F982A4",
-19161 => x"C0C0BFF990F982F9",
-19160 => x"C0C0BFF990F982C0",
-19159 => x"C0C0BFF990F99290",
-19158 => x"C0C0BFF990F99280",
-19157 => x"C0C0BFF990F992F8",
-19156 => x"C0C0BFF990F99282",
-19155 => x"C0C0BFF990F99292",
-19154 => x"C0C0BFF990F99299",
-19153 => x"C0C0BFF990F992B0",
-19152 => x"C0C0BFF990F992A4",
-19151 => x"C0C0BFF990F992F9",
-19150 => x"C0C0BFF990F992C0",
-19149 => x"C0C0BFF990F99990",
-19148 => x"C0C0BFF990F99980",
-19147 => x"C0C0BFF990F999F8",
-19146 => x"C0C0BFF990F99982",
-19145 => x"C0C0BFF990F99992",
-19144 => x"C0C0BFF990F99999",
-19143 => x"C0C0BFF990F999B0",
-19142 => x"C0C0BFF990F999A4",
-19141 => x"C0C0BFF990F999F9",
-19140 => x"C0C0BFF990F999C0",
-19139 => x"C0C0BFF990F9B090",
-19138 => x"C0C0BFF990F9B080",
-19137 => x"C0C0BFF990F9B0F8",
-19136 => x"C0C0BFF990F9B082",
-19135 => x"C0C0BFF990F9B092",
-19134 => x"C0C0BFF990F9B099",
-19133 => x"C0C0BFF990F9B0B0",
-19132 => x"C0C0BFF990F9B0A4",
-19131 => x"C0C0BFF990F9B0F9",
-19130 => x"C0C0BFF990F9B0C0",
-19129 => x"C0C0BFF990F9A490",
-19128 => x"C0C0BFF990F9A480",
-19127 => x"C0C0BFF990F9A4F8",
-19126 => x"C0C0BFF990F9A482",
-19125 => x"C0C0BFF990F9A492",
-19124 => x"C0C0BFF990F9A499",
-19123 => x"C0C0BFF990F9A4B0",
-19122 => x"C0C0BFF990F9A4A4",
-19121 => x"C0C0BFF990F9A4F9",
-19120 => x"C0C0BFF990F9A4C0",
-19119 => x"C0C0BFF990F9F990",
-19118 => x"C0C0BFF990F9F980",
-19117 => x"C0C0BFF990F9F9F8",
-19116 => x"C0C0BFF990F9F982",
-19115 => x"C0C0BFF990F9F992",
-19114 => x"C0C0BFF990F9F999",
-19113 => x"C0C0BFF990F9F9B0",
-19112 => x"C0C0BFF990F9F9A4",
-19111 => x"C0C0BFF990F9F9F9",
-19110 => x"C0C0BFF990F9F9C0",
-19109 => x"C0C0BFF990F9C090",
-19108 => x"C0C0BFF990F9C080",
-19107 => x"C0C0BFF990F9C0F8",
-19106 => x"C0C0BFF990F9C082",
-19105 => x"C0C0BFF990F9C092",
-19104 => x"C0C0BFF990F9C099",
-19103 => x"C0C0BFF990F9C0B0",
-19102 => x"C0C0BFF990F9C0A4",
-19101 => x"C0C0BFF990F9C0F9",
-19100 => x"C0C0BFF990F9C0C0",
-19099 => x"C0C0BFF990C09090",
-19098 => x"C0C0BFF990C09080",
-19097 => x"C0C0BFF990C090F8",
-19096 => x"C0C0BFF990C09082",
-19095 => x"C0C0BFF990C09092",
-19094 => x"C0C0BFF990C09099",
-19093 => x"C0C0BFF990C090B0",
-19092 => x"C0C0BFF990C090A4",
-19091 => x"C0C0BFF990C090F9",
-19090 => x"C0C0BFF990C090C0",
-19089 => x"C0C0BFF990C08090",
-19088 => x"C0C0BFF990C08080",
-19087 => x"C0C0BFF990C080F8",
-19086 => x"C0C0BFF990C08082",
-19085 => x"C0C0BFF990C08092",
-19084 => x"C0C0BFF990C08099",
-19083 => x"C0C0BFF990C080B0",
-19082 => x"C0C0BFF990C080A4",
-19081 => x"C0C0BFF990C080F9",
-19080 => x"C0C0BFF990C080C0",
-19079 => x"C0C0BFF990C0F890",
-19078 => x"C0C0BFF990C0F880",
-19077 => x"C0C0BFF990C0F8F8",
-19076 => x"C0C0BFF990C0F882",
-19075 => x"C0C0BFF990C0F892",
-19074 => x"C0C0BFF990C0F899",
-19073 => x"C0C0BFF990C0F8B0",
-19072 => x"C0C0BFF990C0F8A4",
-19071 => x"C0C0BFF990C0F8F9",
-19070 => x"C0C0BFF990C0F8C0",
-19069 => x"C0C0BFF990C08290",
-19068 => x"C0C0BFF990C08280",
-19067 => x"C0C0BFF990C082F8",
-19066 => x"C0C0BFF990C08282",
-19065 => x"C0C0BFF990C08292",
-19064 => x"C0C0BFF990C08299",
-19063 => x"C0C0BFF990C082B0",
-19062 => x"C0C0BFF990C082A4",
-19061 => x"C0C0BFF990C082F9",
-19060 => x"C0C0BFF990C082C0",
-19059 => x"C0C0BFF990C09290",
-19058 => x"C0C0BFF990C09280",
-19057 => x"C0C0BFF990C092F8",
-19056 => x"C0C0BFF990C09282",
-19055 => x"C0C0BFF990C09292",
-19054 => x"C0C0BFF990C09299",
-19053 => x"C0C0BFF990C092B0",
-19052 => x"C0C0BFF990C092A4",
-19051 => x"C0C0BFF990C092F9",
-19050 => x"C0C0BFF990C092C0",
-19049 => x"C0C0BFF990C09990",
-19048 => x"C0C0BFF990C09980",
-19047 => x"C0C0BFF990C099F8",
-19046 => x"C0C0BFF990C09982",
-19045 => x"C0C0BFF990C09992",
-19044 => x"C0C0BFF990C09999",
-19043 => x"C0C0BFF990C099B0",
-19042 => x"C0C0BFF990C099A4",
-19041 => x"C0C0BFF990C099F9",
-19040 => x"C0C0BFF990C099C0",
-19039 => x"C0C0BFF990C0B090",
-19038 => x"C0C0BFF990C0B080",
-19037 => x"C0C0BFF990C0B0F8",
-19036 => x"C0C0BFF990C0B082",
-19035 => x"C0C0BFF990C0B092",
-19034 => x"C0C0BFF990C0B099",
-19033 => x"C0C0BFF990C0B0B0",
-19032 => x"C0C0BFF990C0B0A4",
-19031 => x"C0C0BFF990C0B0F9",
-19030 => x"C0C0BFF990C0B0C0",
-19029 => x"C0C0BFF990C0A490",
-19028 => x"C0C0BFF990C0A480",
-19027 => x"C0C0BFF990C0A4F8",
-19026 => x"C0C0BFF990C0A482",
-19025 => x"C0C0BFF990C0A492",
-19024 => x"C0C0BFF990C0A499",
-19023 => x"C0C0BFF990C0A4B0",
-19022 => x"C0C0BFF990C0A4A4",
-19021 => x"C0C0BFF990C0A4F9",
-19020 => x"C0C0BFF990C0A4C0",
-19019 => x"C0C0BFF990C0F990",
-19018 => x"C0C0BFF990C0F980",
-19017 => x"C0C0BFF990C0F9F8",
-19016 => x"C0C0BFF990C0F982",
-19015 => x"C0C0BFF990C0F992",
-19014 => x"C0C0BFF990C0F999",
-19013 => x"C0C0BFF990C0F9B0",
-19012 => x"C0C0BFF990C0F9A4",
-19011 => x"C0C0BFF990C0F9F9",
-19010 => x"C0C0BFF990C0F9C0",
-19009 => x"C0C0BFF990C0C090",
-19008 => x"C0C0BFF990C0C080",
-19007 => x"C0C0BFF990C0C0F8",
-19006 => x"C0C0BFF990C0C082",
-19005 => x"C0C0BFF990C0C092",
-19004 => x"C0C0BFF990C0C099",
-19003 => x"C0C0BFF990C0C0B0",
-19002 => x"C0C0BFF990C0C0A4",
-19001 => x"C0C0BFF990C0C0F9",
-19000 => x"C0C0BFF990C0C0C0",
-18999 => x"C0C0BFF980909090",
-18998 => x"C0C0BFF980909080",
-18997 => x"C0C0BFF9809090F8",
-18996 => x"C0C0BFF980909082",
-18995 => x"C0C0BFF980909092",
-18994 => x"C0C0BFF980909099",
-18993 => x"C0C0BFF9809090B0",
-18992 => x"C0C0BFF9809090A4",
-18991 => x"C0C0BFF9809090F9",
-18990 => x"C0C0BFF9809090C0",
-18989 => x"C0C0BFF980908090",
-18988 => x"C0C0BFF980908080",
-18987 => x"C0C0BFF9809080F8",
-18986 => x"C0C0BFF980908082",
-18985 => x"C0C0BFF980908092",
-18984 => x"C0C0BFF980908099",
-18983 => x"C0C0BFF9809080B0",
-18982 => x"C0C0BFF9809080A4",
-18981 => x"C0C0BFF9809080F9",
-18980 => x"C0C0BFF9809080C0",
-18979 => x"C0C0BFF98090F890",
-18978 => x"C0C0BFF98090F880",
-18977 => x"C0C0BFF98090F8F8",
-18976 => x"C0C0BFF98090F882",
-18975 => x"C0C0BFF98090F892",
-18974 => x"C0C0BFF98090F899",
-18973 => x"C0C0BFF98090F8B0",
-18972 => x"C0C0BFF98090F8A4",
-18971 => x"C0C0BFF98090F8F9",
-18970 => x"C0C0BFF98090F8C0",
-18969 => x"C0C0BFF980908290",
-18968 => x"C0C0BFF980908280",
-18967 => x"C0C0BFF9809082F8",
-18966 => x"C0C0BFF980908282",
-18965 => x"C0C0BFF980908292",
-18964 => x"C0C0BFF980908299",
-18963 => x"C0C0BFF9809082B0",
-18962 => x"C0C0BFF9809082A4",
-18961 => x"C0C0BFF9809082F9",
-18960 => x"C0C0BFF9809082C0",
-18959 => x"C0C0BFF980909290",
-18958 => x"C0C0BFF980909280",
-18957 => x"C0C0BFF9809092F8",
-18956 => x"C0C0BFF980909282",
-18955 => x"C0C0BFF980909292",
-18954 => x"C0C0BFF980909299",
-18953 => x"C0C0BFF9809092B0",
-18952 => x"C0C0BFF9809092A4",
-18951 => x"C0C0BFF9809092F9",
-18950 => x"C0C0BFF9809092C0",
-18949 => x"C0C0BFF980909990",
-18948 => x"C0C0BFF980909980",
-18947 => x"C0C0BFF9809099F8",
-18946 => x"C0C0BFF980909982",
-18945 => x"C0C0BFF980909992",
-18944 => x"C0C0BFF980909999",
-18943 => x"C0C0BFF9809099B0",
-18942 => x"C0C0BFF9809099A4",
-18941 => x"C0C0BFF9809099F9",
-18940 => x"C0C0BFF9809099C0",
-18939 => x"C0C0BFF98090B090",
-18938 => x"C0C0BFF98090B080",
-18937 => x"C0C0BFF98090B0F8",
-18936 => x"C0C0BFF98090B082",
-18935 => x"C0C0BFF98090B092",
-18934 => x"C0C0BFF98090B099",
-18933 => x"C0C0BFF98090B0B0",
-18932 => x"C0C0BFF98090B0A4",
-18931 => x"C0C0BFF98090B0F9",
-18930 => x"C0C0BFF98090B0C0",
-18929 => x"C0C0BFF98090A490",
-18928 => x"C0C0BFF98090A480",
-18927 => x"C0C0BFF98090A4F8",
-18926 => x"C0C0BFF98090A482",
-18925 => x"C0C0BFF98090A492",
-18924 => x"C0C0BFF98090A499",
-18923 => x"C0C0BFF98090A4B0",
-18922 => x"C0C0BFF98090A4A4",
-18921 => x"C0C0BFF98090A4F9",
-18920 => x"C0C0BFF98090A4C0",
-18919 => x"C0C0BFF98090F990",
-18918 => x"C0C0BFF98090F980",
-18917 => x"C0C0BFF98090F9F8",
-18916 => x"C0C0BFF98090F982",
-18915 => x"C0C0BFF98090F992",
-18914 => x"C0C0BFF98090F999",
-18913 => x"C0C0BFF98090F9B0",
-18912 => x"C0C0BFF98090F9A4",
-18911 => x"C0C0BFF98090F9F9",
-18910 => x"C0C0BFF98090F9C0",
-18909 => x"C0C0BFF98090C090",
-18908 => x"C0C0BFF98090C080",
-18907 => x"C0C0BFF98090C0F8",
-18906 => x"C0C0BFF98090C082",
-18905 => x"C0C0BFF98090C092",
-18904 => x"C0C0BFF98090C099",
-18903 => x"C0C0BFF98090C0B0",
-18902 => x"C0C0BFF98090C0A4",
-18901 => x"C0C0BFF98090C0F9",
-18900 => x"C0C0BFF98090C0C0",
-18899 => x"C0C0BFF980809090",
-18898 => x"C0C0BFF980809080",
-18897 => x"C0C0BFF9808090F8",
-18896 => x"C0C0BFF980809082",
-18895 => x"C0C0BFF980809092",
-18894 => x"C0C0BFF980809099",
-18893 => x"C0C0BFF9808090B0",
-18892 => x"C0C0BFF9808090A4",
-18891 => x"C0C0BFF9808090F9",
-18890 => x"C0C0BFF9808090C0",
-18889 => x"C0C0BFF980808090",
-18888 => x"C0C0BFF980808080",
-18887 => x"C0C0BFF9808080F8",
-18886 => x"C0C0BFF980808082",
-18885 => x"C0C0BFF980808092",
-18884 => x"C0C0BFF980808099",
-18883 => x"C0C0BFF9808080B0",
-18882 => x"C0C0BFF9808080A4",
-18881 => x"C0C0BFF9808080F9",
-18880 => x"C0C0BFF9808080C0",
-18879 => x"C0C0BFF98080F890",
-18878 => x"C0C0BFF98080F880",
-18877 => x"C0C0BFF98080F8F8",
-18876 => x"C0C0BFF98080F882",
-18875 => x"C0C0BFF98080F892",
-18874 => x"C0C0BFF98080F899",
-18873 => x"C0C0BFF98080F8B0",
-18872 => x"C0C0BFF98080F8A4",
-18871 => x"C0C0BFF98080F8F9",
-18870 => x"C0C0BFF98080F8C0",
-18869 => x"C0C0BFF980808290",
-18868 => x"C0C0BFF980808280",
-18867 => x"C0C0BFF9808082F8",
-18866 => x"C0C0BFF980808282",
-18865 => x"C0C0BFF980808292",
-18864 => x"C0C0BFF980808299",
-18863 => x"C0C0BFF9808082B0",
-18862 => x"C0C0BFF9808082A4",
-18861 => x"C0C0BFF9808082F9",
-18860 => x"C0C0BFF9808082C0",
-18859 => x"C0C0BFF980809290",
-18858 => x"C0C0BFF980809280",
-18857 => x"C0C0BFF9808092F8",
-18856 => x"C0C0BFF980809282",
-18855 => x"C0C0BFF980809292",
-18854 => x"C0C0BFF980809299",
-18853 => x"C0C0BFF9808092B0",
-18852 => x"C0C0BFF9808092A4",
-18851 => x"C0C0BFF9808092F9",
-18850 => x"C0C0BFF9808092C0",
-18849 => x"C0C0BFF980809990",
-18848 => x"C0C0BFF980809980",
-18847 => x"C0C0BFF9808099F8",
-18846 => x"C0C0BFF980809982",
-18845 => x"C0C0BFF980809992",
-18844 => x"C0C0BFF980809999",
-18843 => x"C0C0BFF9808099B0",
-18842 => x"C0C0BFF9808099A4",
-18841 => x"C0C0BFF9808099F9",
-18840 => x"C0C0BFF9808099C0",
-18839 => x"C0C0BFF98080B090",
-18838 => x"C0C0BFF98080B080",
-18837 => x"C0C0BFF98080B0F8",
-18836 => x"C0C0BFF98080B082",
-18835 => x"C0C0BFF98080B092",
-18834 => x"C0C0BFF98080B099",
-18833 => x"C0C0BFF98080B0B0",
-18832 => x"C0C0BFF98080B0A4",
-18831 => x"C0C0BFF98080B0F9",
-18830 => x"C0C0BFF98080B0C0",
-18829 => x"C0C0BFF98080A490",
-18828 => x"C0C0BFF98080A480",
-18827 => x"C0C0BFF98080A4F8",
-18826 => x"C0C0BFF98080A482",
-18825 => x"C0C0BFF98080A492",
-18824 => x"C0C0BFF98080A499",
-18823 => x"C0C0BFF98080A4B0",
-18822 => x"C0C0BFF98080A4A4",
-18821 => x"C0C0BFF98080A4F9",
-18820 => x"C0C0BFF98080A4C0",
-18819 => x"C0C0BFF98080F990",
-18818 => x"C0C0BFF98080F980",
-18817 => x"C0C0BFF98080F9F8",
-18816 => x"C0C0BFF98080F982",
-18815 => x"C0C0BFF98080F992",
-18814 => x"C0C0BFF98080F999",
-18813 => x"C0C0BFF98080F9B0",
-18812 => x"C0C0BFF98080F9A4",
-18811 => x"C0C0BFF98080F9F9",
-18810 => x"C0C0BFF98080F9C0",
-18809 => x"C0C0BFF98080C090",
-18808 => x"C0C0BFF98080C080",
-18807 => x"C0C0BFF98080C0F8",
-18806 => x"C0C0BFF98080C082",
-18805 => x"C0C0BFF98080C092",
-18804 => x"C0C0BFF98080C099",
-18803 => x"C0C0BFF98080C0B0",
-18802 => x"C0C0BFF98080C0A4",
-18801 => x"C0C0BFF98080C0F9",
-18800 => x"C0C0BFF98080C0C0",
-18799 => x"C0C0BFF980F89090",
-18798 => x"C0C0BFF980F89080",
-18797 => x"C0C0BFF980F890F8",
-18796 => x"C0C0BFF980F89082",
-18795 => x"C0C0BFF980F89092",
-18794 => x"C0C0BFF980F89099",
-18793 => x"C0C0BFF980F890B0",
-18792 => x"C0C0BFF980F890A4",
-18791 => x"C0C0BFF980F890F9",
-18790 => x"C0C0BFF980F890C0",
-18789 => x"C0C0BFF980F88090",
-18788 => x"C0C0BFF980F88080",
-18787 => x"C0C0BFF980F880F8",
-18786 => x"C0C0BFF980F88082",
-18785 => x"C0C0BFF980F88092",
-18784 => x"C0C0BFF980F88099",
-18783 => x"C0C0BFF980F880B0",
-18782 => x"C0C0BFF980F880A4",
-18781 => x"C0C0BFF980F880F9",
-18780 => x"C0C0BFF980F880C0",
-18779 => x"C0C0BFF980F8F890",
-18778 => x"C0C0BFF980F8F880",
-18777 => x"C0C0BFF980F8F8F8",
-18776 => x"C0C0BFF980F8F882",
-18775 => x"C0C0BFF980F8F892",
-18774 => x"C0C0BFF980F8F899",
-18773 => x"C0C0BFF980F8F8B0",
-18772 => x"C0C0BFF980F8F8A4",
-18771 => x"C0C0BFF980F8F8F9",
-18770 => x"C0C0BFF980F8F8C0",
-18769 => x"C0C0BFF980F88290",
-18768 => x"C0C0BFF980F88280",
-18767 => x"C0C0BFF980F882F8",
-18766 => x"C0C0BFF980F88282",
-18765 => x"C0C0BFF980F88292",
-18764 => x"C0C0BFF980F88299",
-18763 => x"C0C0BFF980F882B0",
-18762 => x"C0C0BFF980F882A4",
-18761 => x"C0C0BFF980F882F9",
-18760 => x"C0C0BFF980F882C0",
-18759 => x"C0C0BFF980F89290",
-18758 => x"C0C0BFF980F89280",
-18757 => x"C0C0BFF980F892F8",
-18756 => x"C0C0BFF980F89282",
-18755 => x"C0C0BFF980F89292",
-18754 => x"C0C0BFF980F89299",
-18753 => x"C0C0BFF980F892B0",
-18752 => x"C0C0BFF980F892A4",
-18751 => x"C0C0BFF980F892F9",
-18750 => x"C0C0BFF980F892C0",
-18749 => x"C0C0BFF980F89990",
-18748 => x"C0C0BFF980F89980",
-18747 => x"C0C0BFF980F899F8",
-18746 => x"C0C0BFF980F89982",
-18745 => x"C0C0BFF980F89992",
-18744 => x"C0C0BFF980F89999",
-18743 => x"C0C0BFF980F899B0",
-18742 => x"C0C0BFF980F899A4",
-18741 => x"C0C0BFF980F899F9",
-18740 => x"C0C0BFF980F899C0",
-18739 => x"C0C0BFF980F8B090",
-18738 => x"C0C0BFF980F8B080",
-18737 => x"C0C0BFF980F8B0F8",
-18736 => x"C0C0BFF980F8B082",
-18735 => x"C0C0BFF980F8B092",
-18734 => x"C0C0BFF980F8B099",
-18733 => x"C0C0BFF980F8B0B0",
-18732 => x"C0C0BFF980F8B0A4",
-18731 => x"C0C0BFF980F8B0F9",
-18730 => x"C0C0BFF980F8B0C0",
-18729 => x"C0C0BFF980F8A490",
-18728 => x"C0C0BFF980F8A480",
-18727 => x"C0C0BFF980F8A4F8",
-18726 => x"C0C0BFF980F8A482",
-18725 => x"C0C0BFF980F8A492",
-18724 => x"C0C0BFF980F8A499",
-18723 => x"C0C0BFF980F8A4B0",
-18722 => x"C0C0BFF980F8A4A4",
-18721 => x"C0C0BFF980F8A4F9",
-18720 => x"C0C0BFF980F8A4C0",
-18719 => x"C0C0BFF980F8F990",
-18718 => x"C0C0BFF980F8F980",
-18717 => x"C0C0BFF980F8F9F8",
-18716 => x"C0C0BFF980F8F982",
-18715 => x"C0C0BFF980F8F992",
-18714 => x"C0C0BFF980F8F999",
-18713 => x"C0C0BFF980F8F9B0",
-18712 => x"C0C0BFF980F8F9A4",
-18711 => x"C0C0BFF980F8F9F9",
-18710 => x"C0C0BFF980F8F9C0",
-18709 => x"C0C0BFF980F8C090",
-18708 => x"C0C0BFF980F8C080",
-18707 => x"C0C0BFF980F8C0F8",
-18706 => x"C0C0BFF980F8C082",
-18705 => x"C0C0BFF980F8C092",
-18704 => x"C0C0BFF980F8C099",
-18703 => x"C0C0BFF980F8C0B0",
-18702 => x"C0C0BFF980F8C0A4",
-18701 => x"C0C0BFF980F8C0F9",
-18700 => x"C0C0BFF980F8C0C0",
-18699 => x"C0C0BFF980829090",
-18698 => x"C0C0BFF980829080",
-18697 => x"C0C0BFF9808290F8",
-18696 => x"C0C0BFF980829082",
-18695 => x"C0C0BFF980829092",
-18694 => x"C0C0BFF980829099",
-18693 => x"C0C0BFF9808290B0",
-18692 => x"C0C0BFF9808290A4",
-18691 => x"C0C0BFF9808290F9",
-18690 => x"C0C0BFF9808290C0",
-18689 => x"C0C0BFF980828090",
-18688 => x"C0C0BFF980828080",
-18687 => x"C0C0BFF9808280F8",
-18686 => x"C0C0BFF980828082",
-18685 => x"C0C0BFF980828092",
-18684 => x"C0C0BFF980828099",
-18683 => x"C0C0BFF9808280B0",
-18682 => x"C0C0BFF9808280A4",
-18681 => x"C0C0BFF9808280F9",
-18680 => x"C0C0BFF9808280C0",
-18679 => x"C0C0BFF98082F890",
-18678 => x"C0C0BFF98082F880",
-18677 => x"C0C0BFF98082F8F8",
-18676 => x"C0C0BFF98082F882",
-18675 => x"C0C0BFF98082F892",
-18674 => x"C0C0BFF98082F899",
-18673 => x"C0C0BFF98082F8B0",
-18672 => x"C0C0BFF98082F8A4",
-18671 => x"C0C0BFF98082F8F9",
-18670 => x"C0C0BFF98082F8C0",
-18669 => x"C0C0BFF980828290",
-18668 => x"C0C0BFF980828280",
-18667 => x"C0C0BFF9808282F8",
-18666 => x"C0C0BFF980828282",
-18665 => x"C0C0BFF980828292",
-18664 => x"C0C0BFF980828299",
-18663 => x"C0C0BFF9808282B0",
-18662 => x"C0C0BFF9808282A4",
-18661 => x"C0C0BFF9808282F9",
-18660 => x"C0C0BFF9808282C0",
-18659 => x"C0C0BFF980829290",
-18658 => x"C0C0BFF980829280",
-18657 => x"C0C0BFF9808292F8",
-18656 => x"C0C0BFF980829282",
-18655 => x"C0C0BFF980829292",
-18654 => x"C0C0BFF980829299",
-18653 => x"C0C0BFF9808292B0",
-18652 => x"C0C0BFF9808292A4",
-18651 => x"C0C0BFF9808292F9",
-18650 => x"C0C0BFF9808292C0",
-18649 => x"C0C0BFF980829990",
-18648 => x"C0C0BFF980829980",
-18647 => x"C0C0BFF9808299F8",
-18646 => x"C0C0BFF980829982",
-18645 => x"C0C0BFF980829992",
-18644 => x"C0C0BFF980829999",
-18643 => x"C0C0BFF9808299B0",
-18642 => x"C0C0BFF9808299A4",
-18641 => x"C0C0BFF9808299F9",
-18640 => x"C0C0BFF9808299C0",
-18639 => x"C0C0BFF98082B090",
-18638 => x"C0C0BFF98082B080",
-18637 => x"C0C0BFF98082B0F8",
-18636 => x"C0C0BFF98082B082",
-18635 => x"C0C0BFF98082B092",
-18634 => x"C0C0BFF98082B099",
-18633 => x"C0C0BFF98082B0B0",
-18632 => x"C0C0BFF98082B0A4",
-18631 => x"C0C0BFF98082B0F9",
-18630 => x"C0C0BFF98082B0C0",
-18629 => x"C0C0BFF98082A490",
-18628 => x"C0C0BFF98082A480",
-18627 => x"C0C0BFF98082A4F8",
-18626 => x"C0C0BFF98082A482",
-18625 => x"C0C0BFF98082A492",
-18624 => x"C0C0BFF98082A499",
-18623 => x"C0C0BFF98082A4B0",
-18622 => x"C0C0BFF98082A4A4",
-18621 => x"C0C0BFF98082A4F9",
-18620 => x"C0C0BFF98082A4C0",
-18619 => x"C0C0BFF98082F990",
-18618 => x"C0C0BFF98082F980",
-18617 => x"C0C0BFF98082F9F8",
-18616 => x"C0C0BFF98082F982",
-18615 => x"C0C0BFF98082F992",
-18614 => x"C0C0BFF98082F999",
-18613 => x"C0C0BFF98082F9B0",
-18612 => x"C0C0BFF98082F9A4",
-18611 => x"C0C0BFF98082F9F9",
-18610 => x"C0C0BFF98082F9C0",
-18609 => x"C0C0BFF98082C090",
-18608 => x"C0C0BFF98082C080",
-18607 => x"C0C0BFF98082C0F8",
-18606 => x"C0C0BFF98082C082",
-18605 => x"C0C0BFF98082C092",
-18604 => x"C0C0BFF98082C099",
-18603 => x"C0C0BFF98082C0B0",
-18602 => x"C0C0BFF98082C0A4",
-18601 => x"C0C0BFF98082C0F9",
-18600 => x"C0C0BFF98082C0C0",
-18599 => x"C0C0BFF980929090",
-18598 => x"C0C0BFF980929080",
-18597 => x"C0C0BFF9809290F8",
-18596 => x"C0C0BFF980929082",
-18595 => x"C0C0BFF980929092",
-18594 => x"C0C0BFF980929099",
-18593 => x"C0C0BFF9809290B0",
-18592 => x"C0C0BFF9809290A4",
-18591 => x"C0C0BFF9809290F9",
-18590 => x"C0C0BFF9809290C0",
-18589 => x"C0C0BFF980928090",
-18588 => x"C0C0BFF980928080",
-18587 => x"C0C0BFF9809280F8",
-18586 => x"C0C0BFF980928082",
-18585 => x"C0C0BFF980928092",
-18584 => x"C0C0BFF980928099",
-18583 => x"C0C0BFF9809280B0",
-18582 => x"C0C0BFF9809280A4",
-18581 => x"C0C0BFF9809280F9",
-18580 => x"C0C0BFF9809280C0",
-18579 => x"C0C0BFF98092F890",
-18578 => x"C0C0BFF98092F880",
-18577 => x"C0C0BFF98092F8F8",
-18576 => x"C0C0BFF98092F882",
-18575 => x"C0C0BFF98092F892",
-18574 => x"C0C0BFF98092F899",
-18573 => x"C0C0BFF98092F8B0",
-18572 => x"C0C0BFF98092F8A4",
-18571 => x"C0C0BFF98092F8F9",
-18570 => x"C0C0BFF98092F8C0",
-18569 => x"C0C0BFF980928290",
-18568 => x"C0C0BFF980928280",
-18567 => x"C0C0BFF9809282F8",
-18566 => x"C0C0BFF980928282",
-18565 => x"C0C0BFF980928292",
-18564 => x"C0C0BFF980928299",
-18563 => x"C0C0BFF9809282B0",
-18562 => x"C0C0BFF9809282A4",
-18561 => x"C0C0BFF9809282F9",
-18560 => x"C0C0BFF9809282C0",
-18559 => x"C0C0BFF980929290",
-18558 => x"C0C0BFF980929280",
-18557 => x"C0C0BFF9809292F8",
-18556 => x"C0C0BFF980929282",
-18555 => x"C0C0BFF980929292",
-18554 => x"C0C0BFF980929299",
-18553 => x"C0C0BFF9809292B0",
-18552 => x"C0C0BFF9809292A4",
-18551 => x"C0C0BFF9809292F9",
-18550 => x"C0C0BFF9809292C0",
-18549 => x"C0C0BFF980929990",
-18548 => x"C0C0BFF980929980",
-18547 => x"C0C0BFF9809299F8",
-18546 => x"C0C0BFF980929982",
-18545 => x"C0C0BFF980929992",
-18544 => x"C0C0BFF980929999",
-18543 => x"C0C0BFF9809299B0",
-18542 => x"C0C0BFF9809299A4",
-18541 => x"C0C0BFF9809299F9",
-18540 => x"C0C0BFF9809299C0",
-18539 => x"C0C0BFF98092B090",
-18538 => x"C0C0BFF98092B080",
-18537 => x"C0C0BFF98092B0F8",
-18536 => x"C0C0BFF98092B082",
-18535 => x"C0C0BFF98092B092",
-18534 => x"C0C0BFF98092B099",
-18533 => x"C0C0BFF98092B0B0",
-18532 => x"C0C0BFF98092B0A4",
-18531 => x"C0C0BFF98092B0F9",
-18530 => x"C0C0BFF98092B0C0",
-18529 => x"C0C0BFF98092A490",
-18528 => x"C0C0BFF98092A480",
-18527 => x"C0C0BFF98092A4F8",
-18526 => x"C0C0BFF98092A482",
-18525 => x"C0C0BFF98092A492",
-18524 => x"C0C0BFF98092A499",
-18523 => x"C0C0BFF98092A4B0",
-18522 => x"C0C0BFF98092A4A4",
-18521 => x"C0C0BFF98092A4F9",
-18520 => x"C0C0BFF98092A4C0",
-18519 => x"C0C0BFF98092F990",
-18518 => x"C0C0BFF98092F980",
-18517 => x"C0C0BFF98092F9F8",
-18516 => x"C0C0BFF98092F982",
-18515 => x"C0C0BFF98092F992",
-18514 => x"C0C0BFF98092F999",
-18513 => x"C0C0BFF98092F9B0",
-18512 => x"C0C0BFF98092F9A4",
-18511 => x"C0C0BFF98092F9F9",
-18510 => x"C0C0BFF98092F9C0",
-18509 => x"C0C0BFF98092C090",
-18508 => x"C0C0BFF98092C080",
-18507 => x"C0C0BFF98092C0F8",
-18506 => x"C0C0BFF98092C082",
-18505 => x"C0C0BFF98092C092",
-18504 => x"C0C0BFF98092C099",
-18503 => x"C0C0BFF98092C0B0",
-18502 => x"C0C0BFF98092C0A4",
-18501 => x"C0C0BFF98092C0F9",
-18500 => x"C0C0BFF98092C0C0",
-18499 => x"C0C0BFF980999090",
-18498 => x"C0C0BFF980999080",
-18497 => x"C0C0BFF9809990F8",
-18496 => x"C0C0BFF980999082",
-18495 => x"C0C0BFF980999092",
-18494 => x"C0C0BFF980999099",
-18493 => x"C0C0BFF9809990B0",
-18492 => x"C0C0BFF9809990A4",
-18491 => x"C0C0BFF9809990F9",
-18490 => x"C0C0BFF9809990C0",
-18489 => x"C0C0BFF980998090",
-18488 => x"C0C0BFF980998080",
-18487 => x"C0C0BFF9809980F8",
-18486 => x"C0C0BFF980998082",
-18485 => x"C0C0BFF980998092",
-18484 => x"C0C0BFF980998099",
-18483 => x"C0C0BFF9809980B0",
-18482 => x"C0C0BFF9809980A4",
-18481 => x"C0C0BFF9809980F9",
-18480 => x"C0C0BFF9809980C0",
-18479 => x"C0C0BFF98099F890",
-18478 => x"C0C0BFF98099F880",
-18477 => x"C0C0BFF98099F8F8",
-18476 => x"C0C0BFF98099F882",
-18475 => x"C0C0BFF98099F892",
-18474 => x"C0C0BFF98099F899",
-18473 => x"C0C0BFF98099F8B0",
-18472 => x"C0C0BFF98099F8A4",
-18471 => x"C0C0BFF98099F8F9",
-18470 => x"C0C0BFF98099F8C0",
-18469 => x"C0C0BFF980998290",
-18468 => x"C0C0BFF980998280",
-18467 => x"C0C0BFF9809982F8",
-18466 => x"C0C0BFF980998282",
-18465 => x"C0C0BFF980998292",
-18464 => x"C0C0BFF980998299",
-18463 => x"C0C0BFF9809982B0",
-18462 => x"C0C0BFF9809982A4",
-18461 => x"C0C0BFF9809982F9",
-18460 => x"C0C0BFF9809982C0",
-18459 => x"C0C0BFF980999290",
-18458 => x"C0C0BFF980999280",
-18457 => x"C0C0BFF9809992F8",
-18456 => x"C0C0BFF980999282",
-18455 => x"C0C0BFF980999292",
-18454 => x"C0C0BFF980999299",
-18453 => x"C0C0BFF9809992B0",
-18452 => x"C0C0BFF9809992A4",
-18451 => x"C0C0BFF9809992F9",
-18450 => x"C0C0BFF9809992C0",
-18449 => x"C0C0BFF980999990",
-18448 => x"C0C0BFF980999980",
-18447 => x"C0C0BFF9809999F8",
-18446 => x"C0C0BFF980999982",
-18445 => x"C0C0BFF980999992",
-18444 => x"C0C0BFF980999999",
-18443 => x"C0C0BFF9809999B0",
-18442 => x"C0C0BFF9809999A4",
-18441 => x"C0C0BFF9809999F9",
-18440 => x"C0C0BFF9809999C0",
-18439 => x"C0C0BFF98099B090",
-18438 => x"C0C0BFF98099B080",
-18437 => x"C0C0BFF98099B0F8",
-18436 => x"C0C0BFF98099B082",
-18435 => x"C0C0BFF98099B092",
-18434 => x"C0C0BFF98099B099",
-18433 => x"C0C0BFF98099B0B0",
-18432 => x"C0C0BFF98099B0A4",
-18431 => x"C0C0BFF98099B0F9",
-18430 => x"C0C0BFF98099B0C0",
-18429 => x"C0C0BFF98099A490",
-18428 => x"C0C0BFF98099A480",
-18427 => x"C0C0BFF98099A4F8",
-18426 => x"C0C0BFF98099A482",
-18425 => x"C0C0BFF98099A492",
-18424 => x"C0C0BFF98099A499",
-18423 => x"C0C0BFF98099A4B0",
-18422 => x"C0C0BFF98099A4A4",
-18421 => x"C0C0BFF98099A4F9",
-18420 => x"C0C0BFF98099A4C0",
-18419 => x"C0C0BFF98099F990",
-18418 => x"C0C0BFF98099F980",
-18417 => x"C0C0BFF98099F9F8",
-18416 => x"C0C0BFF98099F982",
-18415 => x"C0C0BFF98099F992",
-18414 => x"C0C0BFF98099F999",
-18413 => x"C0C0BFF98099F9B0",
-18412 => x"C0C0BFF98099F9A4",
-18411 => x"C0C0BFF98099F9F9",
-18410 => x"C0C0BFF98099F9C0",
-18409 => x"C0C0BFF98099C090",
-18408 => x"C0C0BFF98099C080",
-18407 => x"C0C0BFF98099C0F8",
-18406 => x"C0C0BFF98099C082",
-18405 => x"C0C0BFF98099C092",
-18404 => x"C0C0BFF98099C099",
-18403 => x"C0C0BFF98099C0B0",
-18402 => x"C0C0BFF98099C0A4",
-18401 => x"C0C0BFF98099C0F9",
-18400 => x"C0C0BFF98099C0C0",
-18399 => x"C0C0BFF980B09090",
-18398 => x"C0C0BFF980B09080",
-18397 => x"C0C0BFF980B090F8",
-18396 => x"C0C0BFF980B09082",
-18395 => x"C0C0BFF980B09092",
-18394 => x"C0C0BFF980B09099",
-18393 => x"C0C0BFF980B090B0",
-18392 => x"C0C0BFF980B090A4",
-18391 => x"C0C0BFF980B090F9",
-18390 => x"C0C0BFF980B090C0",
-18389 => x"C0C0BFF980B08090",
-18388 => x"C0C0BFF980B08080",
-18387 => x"C0C0BFF980B080F8",
-18386 => x"C0C0BFF980B08082",
-18385 => x"C0C0BFF980B08092",
-18384 => x"C0C0BFF980B08099",
-18383 => x"C0C0BFF980B080B0",
-18382 => x"C0C0BFF980B080A4",
-18381 => x"C0C0BFF980B080F9",
-18380 => x"C0C0BFF980B080C0",
-18379 => x"C0C0BFF980B0F890",
-18378 => x"C0C0BFF980B0F880",
-18377 => x"C0C0BFF980B0F8F8",
-18376 => x"C0C0BFF980B0F882",
-18375 => x"C0C0BFF980B0F892",
-18374 => x"C0C0BFF980B0F899",
-18373 => x"C0C0BFF980B0F8B0",
-18372 => x"C0C0BFF980B0F8A4",
-18371 => x"C0C0BFF980B0F8F9",
-18370 => x"C0C0BFF980B0F8C0",
-18369 => x"C0C0BFF980B08290",
-18368 => x"C0C0BFF980B08280",
-18367 => x"C0C0BFF980B082F8",
-18366 => x"C0C0BFF980B08282",
-18365 => x"C0C0BFF980B08292",
-18364 => x"C0C0BFF980B08299",
-18363 => x"C0C0BFF980B082B0",
-18362 => x"C0C0BFF980B082A4",
-18361 => x"C0C0BFF980B082F9",
-18360 => x"C0C0BFF980B082C0",
-18359 => x"C0C0BFF980B09290",
-18358 => x"C0C0BFF980B09280",
-18357 => x"C0C0BFF980B092F8",
-18356 => x"C0C0BFF980B09282",
-18355 => x"C0C0BFF980B09292",
-18354 => x"C0C0BFF980B09299",
-18353 => x"C0C0BFF980B092B0",
-18352 => x"C0C0BFF980B092A4",
-18351 => x"C0C0BFF980B092F9",
-18350 => x"C0C0BFF980B092C0",
-18349 => x"C0C0BFF980B09990",
-18348 => x"C0C0BFF980B09980",
-18347 => x"C0C0BFF980B099F8",
-18346 => x"C0C0BFF980B09982",
-18345 => x"C0C0BFF980B09992",
-18344 => x"C0C0BFF980B09999",
-18343 => x"C0C0BFF980B099B0",
-18342 => x"C0C0BFF980B099A4",
-18341 => x"C0C0BFF980B099F9",
-18340 => x"C0C0BFF980B099C0",
-18339 => x"C0C0BFF980B0B090",
-18338 => x"C0C0BFF980B0B080",
-18337 => x"C0C0BFF980B0B0F8",
-18336 => x"C0C0BFF980B0B082",
-18335 => x"C0C0BFF980B0B092",
-18334 => x"C0C0BFF980B0B099",
-18333 => x"C0C0BFF980B0B0B0",
-18332 => x"C0C0BFF980B0B0A4",
-18331 => x"C0C0BFF980B0B0F9",
-18330 => x"C0C0BFF980B0B0C0",
-18329 => x"C0C0BFF980B0A490",
-18328 => x"C0C0BFF980B0A480",
-18327 => x"C0C0BFF980B0A4F8",
-18326 => x"C0C0BFF980B0A482",
-18325 => x"C0C0BFF980B0A492",
-18324 => x"C0C0BFF980B0A499",
-18323 => x"C0C0BFF980B0A4B0",
-18322 => x"C0C0BFF980B0A4A4",
-18321 => x"C0C0BFF980B0A4F9",
-18320 => x"C0C0BFF980B0A4C0",
-18319 => x"C0C0BFF980B0F990",
-18318 => x"C0C0BFF980B0F980",
-18317 => x"C0C0BFF980B0F9F8",
-18316 => x"C0C0BFF980B0F982",
-18315 => x"C0C0BFF980B0F992",
-18314 => x"C0C0BFF980B0F999",
-18313 => x"C0C0BFF980B0F9B0",
-18312 => x"C0C0BFF980B0F9A4",
-18311 => x"C0C0BFF980B0F9F9",
-18310 => x"C0C0BFF980B0F9C0",
-18309 => x"C0C0BFF980B0C090",
-18308 => x"C0C0BFF980B0C080",
-18307 => x"C0C0BFF980B0C0F8",
-18306 => x"C0C0BFF980B0C082",
-18305 => x"C0C0BFF980B0C092",
-18304 => x"C0C0BFF980B0C099",
-18303 => x"C0C0BFF980B0C0B0",
-18302 => x"C0C0BFF980B0C0A4",
-18301 => x"C0C0BFF980B0C0F9",
-18300 => x"C0C0BFF980B0C0C0",
-18299 => x"C0C0BFF980A49090",
-18298 => x"C0C0BFF980A49080",
-18297 => x"C0C0BFF980A490F8",
-18296 => x"C0C0BFF980A49082",
-18295 => x"C0C0BFF980A49092",
-18294 => x"C0C0BFF980A49099",
-18293 => x"C0C0BFF980A490B0",
-18292 => x"C0C0BFF980A490A4",
-18291 => x"C0C0BFF980A490F9",
-18290 => x"C0C0BFF980A490C0",
-18289 => x"C0C0BFF980A48090",
-18288 => x"C0C0BFF980A48080",
-18287 => x"C0C0BFF980A480F8",
-18286 => x"C0C0BFF980A48082",
-18285 => x"C0C0BFF980A48092",
-18284 => x"C0C0BFF980A48099",
-18283 => x"C0C0BFF980A480B0",
-18282 => x"C0C0BFF980A480A4",
-18281 => x"C0C0BFF980A480F9",
-18280 => x"C0C0BFF980A480C0",
-18279 => x"C0C0BFF980A4F890",
-18278 => x"C0C0BFF980A4F880",
-18277 => x"C0C0BFF980A4F8F8",
-18276 => x"C0C0BFF980A4F882",
-18275 => x"C0C0BFF980A4F892",
-18274 => x"C0C0BFF980A4F899",
-18273 => x"C0C0BFF980A4F8B0",
-18272 => x"C0C0BFF980A4F8A4",
-18271 => x"C0C0BFF980A4F8F9",
-18270 => x"C0C0BFF980A4F8C0",
-18269 => x"C0C0BFF980A48290",
-18268 => x"C0C0BFF980A48280",
-18267 => x"C0C0BFF980A482F8",
-18266 => x"C0C0BFF980A48282",
-18265 => x"C0C0BFF980A48292",
-18264 => x"C0C0BFF980A48299",
-18263 => x"C0C0BFF980A482B0",
-18262 => x"C0C0BFF980A482A4",
-18261 => x"C0C0BFF980A482F9",
-18260 => x"C0C0BFF980A482C0",
-18259 => x"C0C0BFF980A49290",
-18258 => x"C0C0BFF980A49280",
-18257 => x"C0C0BFF980A492F8",
-18256 => x"C0C0BFF980A49282",
-18255 => x"C0C0BFF980A49292",
-18254 => x"C0C0BFF980A49299",
-18253 => x"C0C0BFF980A492B0",
-18252 => x"C0C0BFF980A492A4",
-18251 => x"C0C0BFF980A492F9",
-18250 => x"C0C0BFF980A492C0",
-18249 => x"C0C0BFF980A49990",
-18248 => x"C0C0BFF980A49980",
-18247 => x"C0C0BFF980A499F8",
-18246 => x"C0C0BFF980A49982",
-18245 => x"C0C0BFF980A49992",
-18244 => x"C0C0BFF980A49999",
-18243 => x"C0C0BFF980A499B0",
-18242 => x"C0C0BFF980A499A4",
-18241 => x"C0C0BFF980A499F9",
-18240 => x"C0C0BFF980A499C0",
-18239 => x"C0C0BFF980A4B090",
-18238 => x"C0C0BFF980A4B080",
-18237 => x"C0C0BFF980A4B0F8",
-18236 => x"C0C0BFF980A4B082",
-18235 => x"C0C0BFF980A4B092",
-18234 => x"C0C0BFF980A4B099",
-18233 => x"C0C0BFF980A4B0B0",
-18232 => x"C0C0BFF980A4B0A4",
-18231 => x"C0C0BFF980A4B0F9",
-18230 => x"C0C0BFF980A4B0C0",
-18229 => x"C0C0BFF980A4A490",
-18228 => x"C0C0BFF980A4A480",
-18227 => x"C0C0BFF980A4A4F8",
-18226 => x"C0C0BFF980A4A482",
-18225 => x"C0C0BFF980A4A492",
-18224 => x"C0C0BFF980A4A499",
-18223 => x"C0C0BFF980A4A4B0",
-18222 => x"C0C0BFF980A4A4A4",
-18221 => x"C0C0BFF980A4A4F9",
-18220 => x"C0C0BFF980A4A4C0",
-18219 => x"C0C0BFF980A4F990",
-18218 => x"C0C0BFF980A4F980",
-18217 => x"C0C0BFF980A4F9F8",
-18216 => x"C0C0BFF980A4F982",
-18215 => x"C0C0BFF980A4F992",
-18214 => x"C0C0BFF980A4F999",
-18213 => x"C0C0BFF980A4F9B0",
-18212 => x"C0C0BFF980A4F9A4",
-18211 => x"C0C0BFF980A4F9F9",
-18210 => x"C0C0BFF980A4F9C0",
-18209 => x"C0C0BFF980A4C090",
-18208 => x"C0C0BFF980A4C080",
-18207 => x"C0C0BFF980A4C0F8",
-18206 => x"C0C0BFF980A4C082",
-18205 => x"C0C0BFF980A4C092",
-18204 => x"C0C0BFF980A4C099",
-18203 => x"C0C0BFF980A4C0B0",
-18202 => x"C0C0BFF980A4C0A4",
-18201 => x"C0C0BFF980A4C0F9",
-18200 => x"C0C0BFF980A4C0C0",
-18199 => x"C0C0BFF980F99090",
-18198 => x"C0C0BFF980F99080",
-18197 => x"C0C0BFF980F990F8",
-18196 => x"C0C0BFF980F99082",
-18195 => x"C0C0BFF980F99092",
-18194 => x"C0C0BFF980F99099",
-18193 => x"C0C0BFF980F990B0",
-18192 => x"C0C0BFF980F990A4",
-18191 => x"C0C0BFF980F990F9",
-18190 => x"C0C0BFF980F990C0",
-18189 => x"C0C0BFF980F98090",
-18188 => x"C0C0BFF980F98080",
-18187 => x"C0C0BFF980F980F8",
-18186 => x"C0C0BFF980F98082",
-18185 => x"C0C0BFF980F98092",
-18184 => x"C0C0BFF980F98099",
-18183 => x"C0C0BFF980F980B0",
-18182 => x"C0C0BFF980F980A4",
-18181 => x"C0C0BFF980F980F9",
-18180 => x"C0C0BFF980F980C0",
-18179 => x"C0C0BFF980F9F890",
-18178 => x"C0C0BFF980F9F880",
-18177 => x"C0C0BFF980F9F8F8",
-18176 => x"C0C0BFF980F9F882",
-18175 => x"C0C0BFF980F9F892",
-18174 => x"C0C0BFF980F9F899",
-18173 => x"C0C0BFF980F9F8B0",
-18172 => x"C0C0BFF980F9F8A4",
-18171 => x"C0C0BFF980F9F8F9",
-18170 => x"C0C0BFF980F9F8C0",
-18169 => x"C0C0BFF980F98290",
-18168 => x"C0C0BFF980F98280",
-18167 => x"C0C0BFF980F982F8",
-18166 => x"C0C0BFF980F98282",
-18165 => x"C0C0BFF980F98292",
-18164 => x"C0C0BFF980F98299",
-18163 => x"C0C0BFF980F982B0",
-18162 => x"C0C0BFF980F982A4",
-18161 => x"C0C0BFF980F982F9",
-18160 => x"C0C0BFF980F982C0",
-18159 => x"C0C0BFF980F99290",
-18158 => x"C0C0BFF980F99280",
-18157 => x"C0C0BFF980F992F8",
-18156 => x"C0C0BFF980F99282",
-18155 => x"C0C0BFF980F99292",
-18154 => x"C0C0BFF980F99299",
-18153 => x"C0C0BFF980F992B0",
-18152 => x"C0C0BFF980F992A4",
-18151 => x"C0C0BFF980F992F9",
-18150 => x"C0C0BFF980F992C0",
-18149 => x"C0C0BFF980F99990",
-18148 => x"C0C0BFF980F99980",
-18147 => x"C0C0BFF980F999F8",
-18146 => x"C0C0BFF980F99982",
-18145 => x"C0C0BFF980F99992",
-18144 => x"C0C0BFF980F99999",
-18143 => x"C0C0BFF980F999B0",
-18142 => x"C0C0BFF980F999A4",
-18141 => x"C0C0BFF980F999F9",
-18140 => x"C0C0BFF980F999C0",
-18139 => x"C0C0BFF980F9B090",
-18138 => x"C0C0BFF980F9B080",
-18137 => x"C0C0BFF980F9B0F8",
-18136 => x"C0C0BFF980F9B082",
-18135 => x"C0C0BFF980F9B092",
-18134 => x"C0C0BFF980F9B099",
-18133 => x"C0C0BFF980F9B0B0",
-18132 => x"C0C0BFF980F9B0A4",
-18131 => x"C0C0BFF980F9B0F9",
-18130 => x"C0C0BFF980F9B0C0",
-18129 => x"C0C0BFF980F9A490",
-18128 => x"C0C0BFF980F9A480",
-18127 => x"C0C0BFF980F9A4F8",
-18126 => x"C0C0BFF980F9A482",
-18125 => x"C0C0BFF980F9A492",
-18124 => x"C0C0BFF980F9A499",
-18123 => x"C0C0BFF980F9A4B0",
-18122 => x"C0C0BFF980F9A4A4",
-18121 => x"C0C0BFF980F9A4F9",
-18120 => x"C0C0BFF980F9A4C0",
-18119 => x"C0C0BFF980F9F990",
-18118 => x"C0C0BFF980F9F980",
-18117 => x"C0C0BFF980F9F9F8",
-18116 => x"C0C0BFF980F9F982",
-18115 => x"C0C0BFF980F9F992",
-18114 => x"C0C0BFF980F9F999",
-18113 => x"C0C0BFF980F9F9B0",
-18112 => x"C0C0BFF980F9F9A4",
-18111 => x"C0C0BFF980F9F9F9",
-18110 => x"C0C0BFF980F9F9C0",
-18109 => x"C0C0BFF980F9C090",
-18108 => x"C0C0BFF980F9C080",
-18107 => x"C0C0BFF980F9C0F8",
-18106 => x"C0C0BFF980F9C082",
-18105 => x"C0C0BFF980F9C092",
-18104 => x"C0C0BFF980F9C099",
-18103 => x"C0C0BFF980F9C0B0",
-18102 => x"C0C0BFF980F9C0A4",
-18101 => x"C0C0BFF980F9C0F9",
-18100 => x"C0C0BFF980F9C0C0",
-18099 => x"C0C0BFF980C09090",
-18098 => x"C0C0BFF980C09080",
-18097 => x"C0C0BFF980C090F8",
-18096 => x"C0C0BFF980C09082",
-18095 => x"C0C0BFF980C09092",
-18094 => x"C0C0BFF980C09099",
-18093 => x"C0C0BFF980C090B0",
-18092 => x"C0C0BFF980C090A4",
-18091 => x"C0C0BFF980C090F9",
-18090 => x"C0C0BFF980C090C0",
-18089 => x"C0C0BFF980C08090",
-18088 => x"C0C0BFF980C08080",
-18087 => x"C0C0BFF980C080F8",
-18086 => x"C0C0BFF980C08082",
-18085 => x"C0C0BFF980C08092",
-18084 => x"C0C0BFF980C08099",
-18083 => x"C0C0BFF980C080B0",
-18082 => x"C0C0BFF980C080A4",
-18081 => x"C0C0BFF980C080F9",
-18080 => x"C0C0BFF980C080C0",
-18079 => x"C0C0BFF980C0F890",
-18078 => x"C0C0BFF980C0F880",
-18077 => x"C0C0BFF980C0F8F8",
-18076 => x"C0C0BFF980C0F882",
-18075 => x"C0C0BFF980C0F892",
-18074 => x"C0C0BFF980C0F899",
-18073 => x"C0C0BFF980C0F8B0",
-18072 => x"C0C0BFF980C0F8A4",
-18071 => x"C0C0BFF980C0F8F9",
-18070 => x"C0C0BFF980C0F8C0",
-18069 => x"C0C0BFF980C08290",
-18068 => x"C0C0BFF980C08280",
-18067 => x"C0C0BFF980C082F8",
-18066 => x"C0C0BFF980C08282",
-18065 => x"C0C0BFF980C08292",
-18064 => x"C0C0BFF980C08299",
-18063 => x"C0C0BFF980C082B0",
-18062 => x"C0C0BFF980C082A4",
-18061 => x"C0C0BFF980C082F9",
-18060 => x"C0C0BFF980C082C0",
-18059 => x"C0C0BFF980C09290",
-18058 => x"C0C0BFF980C09280",
-18057 => x"C0C0BFF980C092F8",
-18056 => x"C0C0BFF980C09282",
-18055 => x"C0C0BFF980C09292",
-18054 => x"C0C0BFF980C09299",
-18053 => x"C0C0BFF980C092B0",
-18052 => x"C0C0BFF980C092A4",
-18051 => x"C0C0BFF980C092F9",
-18050 => x"C0C0BFF980C092C0",
-18049 => x"C0C0BFF980C09990",
-18048 => x"C0C0BFF980C09980",
-18047 => x"C0C0BFF980C099F8",
-18046 => x"C0C0BFF980C09982",
-18045 => x"C0C0BFF980C09992",
-18044 => x"C0C0BFF980C09999",
-18043 => x"C0C0BFF980C099B0",
-18042 => x"C0C0BFF980C099A4",
-18041 => x"C0C0BFF980C099F9",
-18040 => x"C0C0BFF980C099C0",
-18039 => x"C0C0BFF980C0B090",
-18038 => x"C0C0BFF980C0B080",
-18037 => x"C0C0BFF980C0B0F8",
-18036 => x"C0C0BFF980C0B082",
-18035 => x"C0C0BFF980C0B092",
-18034 => x"C0C0BFF980C0B099",
-18033 => x"C0C0BFF980C0B0B0",
-18032 => x"C0C0BFF980C0B0A4",
-18031 => x"C0C0BFF980C0B0F9",
-18030 => x"C0C0BFF980C0B0C0",
-18029 => x"C0C0BFF980C0A490",
-18028 => x"C0C0BFF980C0A480",
-18027 => x"C0C0BFF980C0A4F8",
-18026 => x"C0C0BFF980C0A482",
-18025 => x"C0C0BFF980C0A492",
-18024 => x"C0C0BFF980C0A499",
-18023 => x"C0C0BFF980C0A4B0",
-18022 => x"C0C0BFF980C0A4A4",
-18021 => x"C0C0BFF980C0A4F9",
-18020 => x"C0C0BFF980C0A4C0",
-18019 => x"C0C0BFF980C0F990",
-18018 => x"C0C0BFF980C0F980",
-18017 => x"C0C0BFF980C0F9F8",
-18016 => x"C0C0BFF980C0F982",
-18015 => x"C0C0BFF980C0F992",
-18014 => x"C0C0BFF980C0F999",
-18013 => x"C0C0BFF980C0F9B0",
-18012 => x"C0C0BFF980C0F9A4",
-18011 => x"C0C0BFF980C0F9F9",
-18010 => x"C0C0BFF980C0F9C0",
-18009 => x"C0C0BFF980C0C090",
-18008 => x"C0C0BFF980C0C080",
-18007 => x"C0C0BFF980C0C0F8",
-18006 => x"C0C0BFF980C0C082",
-18005 => x"C0C0BFF980C0C092",
-18004 => x"C0C0BFF980C0C099",
-18003 => x"C0C0BFF980C0C0B0",
-18002 => x"C0C0BFF980C0C0A4",
-18001 => x"C0C0BFF980C0C0F9",
-18000 => x"C0C0BFF980C0C0C0",
-17999 => x"C0C0BFF9F8909090",
-17998 => x"C0C0BFF9F8909080",
-17997 => x"C0C0BFF9F89090F8",
-17996 => x"C0C0BFF9F8909082",
-17995 => x"C0C0BFF9F8909092",
-17994 => x"C0C0BFF9F8909099",
-17993 => x"C0C0BFF9F89090B0",
-17992 => x"C0C0BFF9F89090A4",
-17991 => x"C0C0BFF9F89090F9",
-17990 => x"C0C0BFF9F89090C0",
-17989 => x"C0C0BFF9F8908090",
-17988 => x"C0C0BFF9F8908080",
-17987 => x"C0C0BFF9F89080F8",
-17986 => x"C0C0BFF9F8908082",
-17985 => x"C0C0BFF9F8908092",
-17984 => x"C0C0BFF9F8908099",
-17983 => x"C0C0BFF9F89080B0",
-17982 => x"C0C0BFF9F89080A4",
-17981 => x"C0C0BFF9F89080F9",
-17980 => x"C0C0BFF9F89080C0",
-17979 => x"C0C0BFF9F890F890",
-17978 => x"C0C0BFF9F890F880",
-17977 => x"C0C0BFF9F890F8F8",
-17976 => x"C0C0BFF9F890F882",
-17975 => x"C0C0BFF9F890F892",
-17974 => x"C0C0BFF9F890F899",
-17973 => x"C0C0BFF9F890F8B0",
-17972 => x"C0C0BFF9F890F8A4",
-17971 => x"C0C0BFF9F890F8F9",
-17970 => x"C0C0BFF9F890F8C0",
-17969 => x"C0C0BFF9F8908290",
-17968 => x"C0C0BFF9F8908280",
-17967 => x"C0C0BFF9F89082F8",
-17966 => x"C0C0BFF9F8908282",
-17965 => x"C0C0BFF9F8908292",
-17964 => x"C0C0BFF9F8908299",
-17963 => x"C0C0BFF9F89082B0",
-17962 => x"C0C0BFF9F89082A4",
-17961 => x"C0C0BFF9F89082F9",
-17960 => x"C0C0BFF9F89082C0",
-17959 => x"C0C0BFF9F8909290",
-17958 => x"C0C0BFF9F8909280",
-17957 => x"C0C0BFF9F89092F8",
-17956 => x"C0C0BFF9F8909282",
-17955 => x"C0C0BFF9F8909292",
-17954 => x"C0C0BFF9F8909299",
-17953 => x"C0C0BFF9F89092B0",
-17952 => x"C0C0BFF9F89092A4",
-17951 => x"C0C0BFF9F89092F9",
-17950 => x"C0C0BFF9F89092C0",
-17949 => x"C0C0BFF9F8909990",
-17948 => x"C0C0BFF9F8909980",
-17947 => x"C0C0BFF9F89099F8",
-17946 => x"C0C0BFF9F8909982",
-17945 => x"C0C0BFF9F8909992",
-17944 => x"C0C0BFF9F8909999",
-17943 => x"C0C0BFF9F89099B0",
-17942 => x"C0C0BFF9F89099A4",
-17941 => x"C0C0BFF9F89099F9",
-17940 => x"C0C0BFF9F89099C0",
-17939 => x"C0C0BFF9F890B090",
-17938 => x"C0C0BFF9F890B080",
-17937 => x"C0C0BFF9F890B0F8",
-17936 => x"C0C0BFF9F890B082",
-17935 => x"C0C0BFF9F890B092",
-17934 => x"C0C0BFF9F890B099",
-17933 => x"C0C0BFF9F890B0B0",
-17932 => x"C0C0BFF9F890B0A4",
-17931 => x"C0C0BFF9F890B0F9",
-17930 => x"C0C0BFF9F890B0C0",
-17929 => x"C0C0BFF9F890A490",
-17928 => x"C0C0BFF9F890A480",
-17927 => x"C0C0BFF9F890A4F8",
-17926 => x"C0C0BFF9F890A482",
-17925 => x"C0C0BFF9F890A492",
-17924 => x"C0C0BFF9F890A499",
-17923 => x"C0C0BFF9F890A4B0",
-17922 => x"C0C0BFF9F890A4A4",
-17921 => x"C0C0BFF9F890A4F9",
-17920 => x"C0C0BFF9F890A4C0",
-17919 => x"C0C0BFF9F890F990",
-17918 => x"C0C0BFF9F890F980",
-17917 => x"C0C0BFF9F890F9F8",
-17916 => x"C0C0BFF9F890F982",
-17915 => x"C0C0BFF9F890F992",
-17914 => x"C0C0BFF9F890F999",
-17913 => x"C0C0BFF9F890F9B0",
-17912 => x"C0C0BFF9F890F9A4",
-17911 => x"C0C0BFF9F890F9F9",
-17910 => x"C0C0BFF9F890F9C0",
-17909 => x"C0C0BFF9F890C090",
-17908 => x"C0C0BFF9F890C080",
-17907 => x"C0C0BFF9F890C0F8",
-17906 => x"C0C0BFF9F890C082",
-17905 => x"C0C0BFF9F890C092",
-17904 => x"C0C0BFF9F890C099",
-17903 => x"C0C0BFF9F890C0B0",
-17902 => x"C0C0BFF9F890C0A4",
-17901 => x"C0C0BFF9F890C0F9",
-17900 => x"C0C0BFF9F890C0C0",
-17899 => x"C0C0BFF9F8809090",
-17898 => x"C0C0BFF9F8809080",
-17897 => x"C0C0BFF9F88090F8",
-17896 => x"C0C0BFF9F8809082",
-17895 => x"C0C0BFF9F8809092",
-17894 => x"C0C0BFF9F8809099",
-17893 => x"C0C0BFF9F88090B0",
-17892 => x"C0C0BFF9F88090A4",
-17891 => x"C0C0BFF9F88090F9",
-17890 => x"C0C0BFF9F88090C0",
-17889 => x"C0C0BFF9F8808090",
-17888 => x"C0C0BFF9F8808080",
-17887 => x"C0C0BFF9F88080F8",
-17886 => x"C0C0BFF9F8808082",
-17885 => x"C0C0BFF9F8808092",
-17884 => x"C0C0BFF9F8808099",
-17883 => x"C0C0BFF9F88080B0",
-17882 => x"C0C0BFF9F88080A4",
-17881 => x"C0C0BFF9F88080F9",
-17880 => x"C0C0BFF9F88080C0",
-17879 => x"C0C0BFF9F880F890",
-17878 => x"C0C0BFF9F880F880",
-17877 => x"C0C0BFF9F880F8F8",
-17876 => x"C0C0BFF9F880F882",
-17875 => x"C0C0BFF9F880F892",
-17874 => x"C0C0BFF9F880F899",
-17873 => x"C0C0BFF9F880F8B0",
-17872 => x"C0C0BFF9F880F8A4",
-17871 => x"C0C0BFF9F880F8F9",
-17870 => x"C0C0BFF9F880F8C0",
-17869 => x"C0C0BFF9F8808290",
-17868 => x"C0C0BFF9F8808280",
-17867 => x"C0C0BFF9F88082F8",
-17866 => x"C0C0BFF9F8808282",
-17865 => x"C0C0BFF9F8808292",
-17864 => x"C0C0BFF9F8808299",
-17863 => x"C0C0BFF9F88082B0",
-17862 => x"C0C0BFF9F88082A4",
-17861 => x"C0C0BFF9F88082F9",
-17860 => x"C0C0BFF9F88082C0",
-17859 => x"C0C0BFF9F8809290",
-17858 => x"C0C0BFF9F8809280",
-17857 => x"C0C0BFF9F88092F8",
-17856 => x"C0C0BFF9F8809282",
-17855 => x"C0C0BFF9F8809292",
-17854 => x"C0C0BFF9F8809299",
-17853 => x"C0C0BFF9F88092B0",
-17852 => x"C0C0BFF9F88092A4",
-17851 => x"C0C0BFF9F88092F9",
-17850 => x"C0C0BFF9F88092C0",
-17849 => x"C0C0BFF9F8809990",
-17848 => x"C0C0BFF9F8809980",
-17847 => x"C0C0BFF9F88099F8",
-17846 => x"C0C0BFF9F8809982",
-17845 => x"C0C0BFF9F8809992",
-17844 => x"C0C0BFF9F8809999",
-17843 => x"C0C0BFF9F88099B0",
-17842 => x"C0C0BFF9F88099A4",
-17841 => x"C0C0BFF9F88099F9",
-17840 => x"C0C0BFF9F88099C0",
-17839 => x"C0C0BFF9F880B090",
-17838 => x"C0C0BFF9F880B080",
-17837 => x"C0C0BFF9F880B0F8",
-17836 => x"C0C0BFF9F880B082",
-17835 => x"C0C0BFF9F880B092",
-17834 => x"C0C0BFF9F880B099",
-17833 => x"C0C0BFF9F880B0B0",
-17832 => x"C0C0BFF9F880B0A4",
-17831 => x"C0C0BFF9F880B0F9",
-17830 => x"C0C0BFF9F880B0C0",
-17829 => x"C0C0BFF9F880A490",
-17828 => x"C0C0BFF9F880A480",
-17827 => x"C0C0BFF9F880A4F8",
-17826 => x"C0C0BFF9F880A482",
-17825 => x"C0C0BFF9F880A492",
-17824 => x"C0C0BFF9F880A499",
-17823 => x"C0C0BFF9F880A4B0",
-17822 => x"C0C0BFF9F880A4A4",
-17821 => x"C0C0BFF9F880A4F9",
-17820 => x"C0C0BFF9F880A4C0",
-17819 => x"C0C0BFF9F880F990",
-17818 => x"C0C0BFF9F880F980",
-17817 => x"C0C0BFF9F880F9F8",
-17816 => x"C0C0BFF9F880F982",
-17815 => x"C0C0BFF9F880F992",
-17814 => x"C0C0BFF9F880F999",
-17813 => x"C0C0BFF9F880F9B0",
-17812 => x"C0C0BFF9F880F9A4",
-17811 => x"C0C0BFF9F880F9F9",
-17810 => x"C0C0BFF9F880F9C0",
-17809 => x"C0C0BFF9F880C090",
-17808 => x"C0C0BFF9F880C080",
-17807 => x"C0C0BFF9F880C0F8",
-17806 => x"C0C0BFF9F880C082",
-17805 => x"C0C0BFF9F880C092",
-17804 => x"C0C0BFF9F880C099",
-17803 => x"C0C0BFF9F880C0B0",
-17802 => x"C0C0BFF9F880C0A4",
-17801 => x"C0C0BFF9F880C0F9",
-17800 => x"C0C0BFF9F880C0C0",
-17799 => x"C0C0BFF9F8F89090",
-17798 => x"C0C0BFF9F8F89080",
-17797 => x"C0C0BFF9F8F890F8",
-17796 => x"C0C0BFF9F8F89082",
-17795 => x"C0C0BFF9F8F89092",
-17794 => x"C0C0BFF9F8F89099",
-17793 => x"C0C0BFF9F8F890B0",
-17792 => x"C0C0BFF9F8F890A4",
-17791 => x"C0C0BFF9F8F890F9",
-17790 => x"C0C0BFF9F8F890C0",
-17789 => x"C0C0BFF9F8F88090",
-17788 => x"C0C0BFF9F8F88080",
-17787 => x"C0C0BFF9F8F880F8",
-17786 => x"C0C0BFF9F8F88082",
-17785 => x"C0C0BFF9F8F88092",
-17784 => x"C0C0BFF9F8F88099",
-17783 => x"C0C0BFF9F8F880B0",
-17782 => x"C0C0BFF9F8F880A4",
-17781 => x"C0C0BFF9F8F880F9",
-17780 => x"C0C0BFF9F8F880C0",
-17779 => x"C0C0BFF9F8F8F890",
-17778 => x"C0C0BFF9F8F8F880",
-17777 => x"C0C0BFF9F8F8F8F8",
-17776 => x"C0C0BFF9F8F8F882",
-17775 => x"C0C0BFF9F8F8F892",
-17774 => x"C0C0BFF9F8F8F899",
-17773 => x"C0C0BFF9F8F8F8B0",
-17772 => x"C0C0BFF9F8F8F8A4",
-17771 => x"C0C0BFF9F8F8F8F9",
-17770 => x"C0C0BFF9F8F8F8C0",
-17769 => x"C0C0BFF9F8F88290",
-17768 => x"C0C0BFF9F8F88280",
-17767 => x"C0C0BFF9F8F882F8",
-17766 => x"C0C0BFF9F8F88282",
-17765 => x"C0C0BFF9F8F88292",
-17764 => x"C0C0BFF9F8F88299",
-17763 => x"C0C0BFF9F8F882B0",
-17762 => x"C0C0BFF9F8F882A4",
-17761 => x"C0C0BFF9F8F882F9",
-17760 => x"C0C0BFF9F8F882C0",
-17759 => x"C0C0BFF9F8F89290",
-17758 => x"C0C0BFF9F8F89280",
-17757 => x"C0C0BFF9F8F892F8",
-17756 => x"C0C0BFF9F8F89282",
-17755 => x"C0C0BFF9F8F89292",
-17754 => x"C0C0BFF9F8F89299",
-17753 => x"C0C0BFF9F8F892B0",
-17752 => x"C0C0BFF9F8F892A4",
-17751 => x"C0C0BFF9F8F892F9",
-17750 => x"C0C0BFF9F8F892C0",
-17749 => x"C0C0BFF9F8F89990",
-17748 => x"C0C0BFF9F8F89980",
-17747 => x"C0C0BFF9F8F899F8",
-17746 => x"C0C0BFF9F8F89982",
-17745 => x"C0C0BFF9F8F89992",
-17744 => x"C0C0BFF9F8F89999",
-17743 => x"C0C0BFF9F8F899B0",
-17742 => x"C0C0BFF9F8F899A4",
-17741 => x"C0C0BFF9F8F899F9",
-17740 => x"C0C0BFF9F8F899C0",
-17739 => x"C0C0BFF9F8F8B090",
-17738 => x"C0C0BFF9F8F8B080",
-17737 => x"C0C0BFF9F8F8B0F8",
-17736 => x"C0C0BFF9F8F8B082",
-17735 => x"C0C0BFF9F8F8B092",
-17734 => x"C0C0BFF9F8F8B099",
-17733 => x"C0C0BFF9F8F8B0B0",
-17732 => x"C0C0BFF9F8F8B0A4",
-17731 => x"C0C0BFF9F8F8B0F9",
-17730 => x"C0C0BFF9F8F8B0C0",
-17729 => x"C0C0BFF9F8F8A490",
-17728 => x"C0C0BFF9F8F8A480",
-17727 => x"C0C0BFF9F8F8A4F8",
-17726 => x"C0C0BFF9F8F8A482",
-17725 => x"C0C0BFF9F8F8A492",
-17724 => x"C0C0BFF9F8F8A499",
-17723 => x"C0C0BFF9F8F8A4B0",
-17722 => x"C0C0BFF9F8F8A4A4",
-17721 => x"C0C0BFF9F8F8A4F9",
-17720 => x"C0C0BFF9F8F8A4C0",
-17719 => x"C0C0BFF9F8F8F990",
-17718 => x"C0C0BFF9F8F8F980",
-17717 => x"C0C0BFF9F8F8F9F8",
-17716 => x"C0C0BFF9F8F8F982",
-17715 => x"C0C0BFF9F8F8F992",
-17714 => x"C0C0BFF9F8F8F999",
-17713 => x"C0C0BFF9F8F8F9B0",
-17712 => x"C0C0BFF9F8F8F9A4",
-17711 => x"C0C0BFF9F8F8F9F9",
-17710 => x"C0C0BFF9F8F8F9C0",
-17709 => x"C0C0BFF9F8F8C090",
-17708 => x"C0C0BFF9F8F8C080",
-17707 => x"C0C0BFF9F8F8C0F8",
-17706 => x"C0C0BFF9F8F8C082",
-17705 => x"C0C0BFF9F8F8C092",
-17704 => x"C0C0BFF9F8F8C099",
-17703 => x"C0C0BFF9F8F8C0B0",
-17702 => x"C0C0BFF9F8F8C0A4",
-17701 => x"C0C0BFF9F8F8C0F9",
-17700 => x"C0C0BFF9F8F8C0C0",
-17699 => x"C0C0BFF9F8829090",
-17698 => x"C0C0BFF9F8829080",
-17697 => x"C0C0BFF9F88290F8",
-17696 => x"C0C0BFF9F8829082",
-17695 => x"C0C0BFF9F8829092",
-17694 => x"C0C0BFF9F8829099",
-17693 => x"C0C0BFF9F88290B0",
-17692 => x"C0C0BFF9F88290A4",
-17691 => x"C0C0BFF9F88290F9",
-17690 => x"C0C0BFF9F88290C0",
-17689 => x"C0C0BFF9F8828090",
-17688 => x"C0C0BFF9F8828080",
-17687 => x"C0C0BFF9F88280F8",
-17686 => x"C0C0BFF9F8828082",
-17685 => x"C0C0BFF9F8828092",
-17684 => x"C0C0BFF9F8828099",
-17683 => x"C0C0BFF9F88280B0",
-17682 => x"C0C0BFF9F88280A4",
-17681 => x"C0C0BFF9F88280F9",
-17680 => x"C0C0BFF9F88280C0",
-17679 => x"C0C0BFF9F882F890",
-17678 => x"C0C0BFF9F882F880",
-17677 => x"C0C0BFF9F882F8F8",
-17676 => x"C0C0BFF9F882F882",
-17675 => x"C0C0BFF9F882F892",
-17674 => x"C0C0BFF9F882F899",
-17673 => x"C0C0BFF9F882F8B0",
-17672 => x"C0C0BFF9F882F8A4",
-17671 => x"C0C0BFF9F882F8F9",
-17670 => x"C0C0BFF9F882F8C0",
-17669 => x"C0C0BFF9F8828290",
-17668 => x"C0C0BFF9F8828280",
-17667 => x"C0C0BFF9F88282F8",
-17666 => x"C0C0BFF9F8828282",
-17665 => x"C0C0BFF9F8828292",
-17664 => x"C0C0BFF9F8828299",
-17663 => x"C0C0BFF9F88282B0",
-17662 => x"C0C0BFF9F88282A4",
-17661 => x"C0C0BFF9F88282F9",
-17660 => x"C0C0BFF9F88282C0",
-17659 => x"C0C0BFF9F8829290",
-17658 => x"C0C0BFF9F8829280",
-17657 => x"C0C0BFF9F88292F8",
-17656 => x"C0C0BFF9F8829282",
-17655 => x"C0C0BFF9F8829292",
-17654 => x"C0C0BFF9F8829299",
-17653 => x"C0C0BFF9F88292B0",
-17652 => x"C0C0BFF9F88292A4",
-17651 => x"C0C0BFF9F88292F9",
-17650 => x"C0C0BFF9F88292C0",
-17649 => x"C0C0BFF9F8829990",
-17648 => x"C0C0BFF9F8829980",
-17647 => x"C0C0BFF9F88299F8",
-17646 => x"C0C0BFF9F8829982",
-17645 => x"C0C0BFF9F8829992",
-17644 => x"C0C0BFF9F8829999",
-17643 => x"C0C0BFF9F88299B0",
-17642 => x"C0C0BFF9F88299A4",
-17641 => x"C0C0BFF9F88299F9",
-17640 => x"C0C0BFF9F88299C0",
-17639 => x"C0C0BFF9F882B090",
-17638 => x"C0C0BFF9F882B080",
-17637 => x"C0C0BFF9F882B0F8",
-17636 => x"C0C0BFF9F882B082",
-17635 => x"C0C0BFF9F882B092",
-17634 => x"C0C0BFF9F882B099",
-17633 => x"C0C0BFF9F882B0B0",
-17632 => x"C0C0BFF9F882B0A4",
-17631 => x"C0C0BFF9F882B0F9",
-17630 => x"C0C0BFF9F882B0C0",
-17629 => x"C0C0BFF9F882A490",
-17628 => x"C0C0BFF9F882A480",
-17627 => x"C0C0BFF9F882A4F8",
-17626 => x"C0C0BFF9F882A482",
-17625 => x"C0C0BFF9F882A492",
-17624 => x"C0C0BFF9F882A499",
-17623 => x"C0C0BFF9F882A4B0",
-17622 => x"C0C0BFF9F882A4A4",
-17621 => x"C0C0BFF9F882A4F9",
-17620 => x"C0C0BFF9F882A4C0",
-17619 => x"C0C0BFF9F882F990",
-17618 => x"C0C0BFF9F882F980",
-17617 => x"C0C0BFF9F882F9F8",
-17616 => x"C0C0BFF9F882F982",
-17615 => x"C0C0BFF9F882F992",
-17614 => x"C0C0BFF9F882F999",
-17613 => x"C0C0BFF9F882F9B0",
-17612 => x"C0C0BFF9F882F9A4",
-17611 => x"C0C0BFF9F882F9F9",
-17610 => x"C0C0BFF9F882F9C0",
-17609 => x"C0C0BFF9F882C090",
-17608 => x"C0C0BFF9F882C080",
-17607 => x"C0C0BFF9F882C0F8",
-17606 => x"C0C0BFF9F882C082",
-17605 => x"C0C0BFF9F882C092",
-17604 => x"C0C0BFF9F882C099",
-17603 => x"C0C0BFF9F882C0B0",
-17602 => x"C0C0BFF9F882C0A4",
-17601 => x"C0C0BFF9F882C0F9",
-17600 => x"C0C0BFF9F882C0C0",
-17599 => x"C0C0BFF9F8929090",
-17598 => x"C0C0BFF9F8929080",
-17597 => x"C0C0BFF9F89290F8",
-17596 => x"C0C0BFF9F8929082",
-17595 => x"C0C0BFF9F8929092",
-17594 => x"C0C0BFF9F8929099",
-17593 => x"C0C0BFF9F89290B0",
-17592 => x"C0C0BFF9F89290A4",
-17591 => x"C0C0BFF9F89290F9",
-17590 => x"C0C0BFF9F89290C0",
-17589 => x"C0C0BFF9F8928090",
-17588 => x"C0C0BFF9F8928080",
-17587 => x"C0C0BFF9F89280F8",
-17586 => x"C0C0BFF9F8928082",
-17585 => x"C0C0BFF9F8928092",
-17584 => x"C0C0BFF9F8928099",
-17583 => x"C0C0BFF9F89280B0",
-17582 => x"C0C0BFF9F89280A4",
-17581 => x"C0C0BFF9F89280F9",
-17580 => x"C0C0BFF9F89280C0",
-17579 => x"C0C0BFF9F892F890",
-17578 => x"C0C0BFF9F892F880",
-17577 => x"C0C0BFF9F892F8F8",
-17576 => x"C0C0BFF9F892F882",
-17575 => x"C0C0BFF9F892F892",
-17574 => x"C0C0BFF9F892F899",
-17573 => x"C0C0BFF9F892F8B0",
-17572 => x"C0C0BFF9F892F8A4",
-17571 => x"C0C0BFF9F892F8F9",
-17570 => x"C0C0BFF9F892F8C0",
-17569 => x"C0C0BFF9F8928290",
-17568 => x"C0C0BFF9F8928280",
-17567 => x"C0C0BFF9F89282F8",
-17566 => x"C0C0BFF9F8928282",
-17565 => x"C0C0BFF9F8928292",
-17564 => x"C0C0BFF9F8928299",
-17563 => x"C0C0BFF9F89282B0",
-17562 => x"C0C0BFF9F89282A4",
-17561 => x"C0C0BFF9F89282F9",
-17560 => x"C0C0BFF9F89282C0",
-17559 => x"C0C0BFF9F8929290",
-17558 => x"C0C0BFF9F8929280",
-17557 => x"C0C0BFF9F89292F8",
-17556 => x"C0C0BFF9F8929282",
-17555 => x"C0C0BFF9F8929292",
-17554 => x"C0C0BFF9F8929299",
-17553 => x"C0C0BFF9F89292B0",
-17552 => x"C0C0BFF9F89292A4",
-17551 => x"C0C0BFF9F89292F9",
-17550 => x"C0C0BFF9F89292C0",
-17549 => x"C0C0BFF9F8929990",
-17548 => x"C0C0BFF9F8929980",
-17547 => x"C0C0BFF9F89299F8",
-17546 => x"C0C0BFF9F8929982",
-17545 => x"C0C0BFF9F8929992",
-17544 => x"C0C0BFF9F8929999",
-17543 => x"C0C0BFF9F89299B0",
-17542 => x"C0C0BFF9F89299A4",
-17541 => x"C0C0BFF9F89299F9",
-17540 => x"C0C0BFF9F89299C0",
-17539 => x"C0C0BFF9F892B090",
-17538 => x"C0C0BFF9F892B080",
-17537 => x"C0C0BFF9F892B0F8",
-17536 => x"C0C0BFF9F892B082",
-17535 => x"C0C0BFF9F892B092",
-17534 => x"C0C0BFF9F892B099",
-17533 => x"C0C0BFF9F892B0B0",
-17532 => x"C0C0BFF9F892B0A4",
-17531 => x"C0C0BFF9F892B0F9",
-17530 => x"C0C0BFF9F892B0C0",
-17529 => x"C0C0BFF9F892A490",
-17528 => x"C0C0BFF9F892A480",
-17527 => x"C0C0BFF9F892A4F8",
-17526 => x"C0C0BFF9F892A482",
-17525 => x"C0C0BFF9F892A492",
-17524 => x"C0C0BFF9F892A499",
-17523 => x"C0C0BFF9F892A4B0",
-17522 => x"C0C0BFF9F892A4A4",
-17521 => x"C0C0BFF9F892A4F9",
-17520 => x"C0C0BFF9F892A4C0",
-17519 => x"C0C0BFF9F892F990",
-17518 => x"C0C0BFF9F892F980",
-17517 => x"C0C0BFF9F892F9F8",
-17516 => x"C0C0BFF9F892F982",
-17515 => x"C0C0BFF9F892F992",
-17514 => x"C0C0BFF9F892F999",
-17513 => x"C0C0BFF9F892F9B0",
-17512 => x"C0C0BFF9F892F9A4",
-17511 => x"C0C0BFF9F892F9F9",
-17510 => x"C0C0BFF9F892F9C0",
-17509 => x"C0C0BFF9F892C090",
-17508 => x"C0C0BFF9F892C080",
-17507 => x"C0C0BFF9F892C0F8",
-17506 => x"C0C0BFF9F892C082",
-17505 => x"C0C0BFF9F892C092",
-17504 => x"C0C0BFF9F892C099",
-17503 => x"C0C0BFF9F892C0B0",
-17502 => x"C0C0BFF9F892C0A4",
-17501 => x"C0C0BFF9F892C0F9",
-17500 => x"C0C0BFF9F892C0C0",
-17499 => x"C0C0BFF9F8999090",
-17498 => x"C0C0BFF9F8999080",
-17497 => x"C0C0BFF9F89990F8",
-17496 => x"C0C0BFF9F8999082",
-17495 => x"C0C0BFF9F8999092",
-17494 => x"C0C0BFF9F8999099",
-17493 => x"C0C0BFF9F89990B0",
-17492 => x"C0C0BFF9F89990A4",
-17491 => x"C0C0BFF9F89990F9",
-17490 => x"C0C0BFF9F89990C0",
-17489 => x"C0C0BFF9F8998090",
-17488 => x"C0C0BFF9F8998080",
-17487 => x"C0C0BFF9F89980F8",
-17486 => x"C0C0BFF9F8998082",
-17485 => x"C0C0BFF9F8998092",
-17484 => x"C0C0BFF9F8998099",
-17483 => x"C0C0BFF9F89980B0",
-17482 => x"C0C0BFF9F89980A4",
-17481 => x"C0C0BFF9F89980F9",
-17480 => x"C0C0BFF9F89980C0",
-17479 => x"C0C0BFF9F899F890",
-17478 => x"C0C0BFF9F899F880",
-17477 => x"C0C0BFF9F899F8F8",
-17476 => x"C0C0BFF9F899F882",
-17475 => x"C0C0BFF9F899F892",
-17474 => x"C0C0BFF9F899F899",
-17473 => x"C0C0BFF9F899F8B0",
-17472 => x"C0C0BFF9F899F8A4",
-17471 => x"C0C0BFF9F899F8F9",
-17470 => x"C0C0BFF9F899F8C0",
-17469 => x"C0C0BFF9F8998290",
-17468 => x"C0C0BFF9F8998280",
-17467 => x"C0C0BFF9F89982F8",
-17466 => x"C0C0BFF9F8998282",
-17465 => x"C0C0BFF9F8998292",
-17464 => x"C0C0BFF9F8998299",
-17463 => x"C0C0BFF9F89982B0",
-17462 => x"C0C0BFF9F89982A4",
-17461 => x"C0C0BFF9F89982F9",
-17460 => x"C0C0BFF9F89982C0",
-17459 => x"C0C0BFF9F8999290",
-17458 => x"C0C0BFF9F8999280",
-17457 => x"C0C0BFF9F89992F8",
-17456 => x"C0C0BFF9F8999282",
-17455 => x"C0C0BFF9F8999292",
-17454 => x"C0C0BFF9F8999299",
-17453 => x"C0C0BFF9F89992B0",
-17452 => x"C0C0BFF9F89992A4",
-17451 => x"C0C0BFF9F89992F9",
-17450 => x"C0C0BFF9F89992C0",
-17449 => x"C0C0BFF9F8999990",
-17448 => x"C0C0BFF9F8999980",
-17447 => x"C0C0BFF9F89999F8",
-17446 => x"C0C0BFF9F8999982",
-17445 => x"C0C0BFF9F8999992",
-17444 => x"C0C0BFF9F8999999",
-17443 => x"C0C0BFF9F89999B0",
-17442 => x"C0C0BFF9F89999A4",
-17441 => x"C0C0BFF9F89999F9",
-17440 => x"C0C0BFF9F89999C0",
-17439 => x"C0C0BFF9F899B090",
-17438 => x"C0C0BFF9F899B080",
-17437 => x"C0C0BFF9F899B0F8",
-17436 => x"C0C0BFF9F899B082",
-17435 => x"C0C0BFF9F899B092",
-17434 => x"C0C0BFF9F899B099",
-17433 => x"C0C0BFF9F899B0B0",
-17432 => x"C0C0BFF9F899B0A4",
-17431 => x"C0C0BFF9F899B0F9",
-17430 => x"C0C0BFF9F899B0C0",
-17429 => x"C0C0BFF9F899A490",
-17428 => x"C0C0BFF9F899A480",
-17427 => x"C0C0BFF9F899A4F8",
-17426 => x"C0C0BFF9F899A482",
-17425 => x"C0C0BFF9F899A492",
-17424 => x"C0C0BFF9F899A499",
-17423 => x"C0C0BFF9F899A4B0",
-17422 => x"C0C0BFF9F899A4A4",
-17421 => x"C0C0BFF9F899A4F9",
-17420 => x"C0C0BFF9F899A4C0",
-17419 => x"C0C0BFF9F899F990",
-17418 => x"C0C0BFF9F899F980",
-17417 => x"C0C0BFF9F899F9F8",
-17416 => x"C0C0BFF9F899F982",
-17415 => x"C0C0BFF9F899F992",
-17414 => x"C0C0BFF9F899F999",
-17413 => x"C0C0BFF9F899F9B0",
-17412 => x"C0C0BFF9F899F9A4",
-17411 => x"C0C0BFF9F899F9F9",
-17410 => x"C0C0BFF9F899F9C0",
-17409 => x"C0C0BFF9F899C090",
-17408 => x"C0C0BFF9F899C080",
-17407 => x"C0C0BFF9F899C0F8",
-17406 => x"C0C0BFF9F899C082",
-17405 => x"C0C0BFF9F899C092",
-17404 => x"C0C0BFF9F899C099",
-17403 => x"C0C0BFF9F899C0B0",
-17402 => x"C0C0BFF9F899C0A4",
-17401 => x"C0C0BFF9F899C0F9",
-17400 => x"C0C0BFF9F899C0C0",
-17399 => x"C0C0BFF9F8B09090",
-17398 => x"C0C0BFF9F8B09080",
-17397 => x"C0C0BFF9F8B090F8",
-17396 => x"C0C0BFF9F8B09082",
-17395 => x"C0C0BFF9F8B09092",
-17394 => x"C0C0BFF9F8B09099",
-17393 => x"C0C0BFF9F8B090B0",
-17392 => x"C0C0BFF9F8B090A4",
-17391 => x"C0C0BFF9F8B090F9",
-17390 => x"C0C0BFF9F8B090C0",
-17389 => x"C0C0BFF9F8B08090",
-17388 => x"C0C0BFF9F8B08080",
-17387 => x"C0C0BFF9F8B080F8",
-17386 => x"C0C0BFF9F8B08082",
-17385 => x"C0C0BFF9F8B08092",
-17384 => x"C0C0BFF9F8B08099",
-17383 => x"C0C0BFF9F8B080B0",
-17382 => x"C0C0BFF9F8B080A4",
-17381 => x"C0C0BFF9F8B080F9",
-17380 => x"C0C0BFF9F8B080C0",
-17379 => x"C0C0BFF9F8B0F890",
-17378 => x"C0C0BFF9F8B0F880",
-17377 => x"C0C0BFF9F8B0F8F8",
-17376 => x"C0C0BFF9F8B0F882",
-17375 => x"C0C0BFF9F8B0F892",
-17374 => x"C0C0BFF9F8B0F899",
-17373 => x"C0C0BFF9F8B0F8B0",
-17372 => x"C0C0BFF9F8B0F8A4",
-17371 => x"C0C0BFF9F8B0F8F9",
-17370 => x"C0C0BFF9F8B0F8C0",
-17369 => x"C0C0BFF9F8B08290",
-17368 => x"C0C0BFF9F8B08280",
-17367 => x"C0C0BFF9F8B082F8",
-17366 => x"C0C0BFF9F8B08282",
-17365 => x"C0C0BFF9F8B08292",
-17364 => x"C0C0BFF9F8B08299",
-17363 => x"C0C0BFF9F8B082B0",
-17362 => x"C0C0BFF9F8B082A4",
-17361 => x"C0C0BFF9F8B082F9",
-17360 => x"C0C0BFF9F8B082C0",
-17359 => x"C0C0BFF9F8B09290",
-17358 => x"C0C0BFF9F8B09280",
-17357 => x"C0C0BFF9F8B092F8",
-17356 => x"C0C0BFF9F8B09282",
-17355 => x"C0C0BFF9F8B09292",
-17354 => x"C0C0BFF9F8B09299",
-17353 => x"C0C0BFF9F8B092B0",
-17352 => x"C0C0BFF9F8B092A4",
-17351 => x"C0C0BFF9F8B092F9",
-17350 => x"C0C0BFF9F8B092C0",
-17349 => x"C0C0BFF9F8B09990",
-17348 => x"C0C0BFF9F8B09980",
-17347 => x"C0C0BFF9F8B099F8",
-17346 => x"C0C0BFF9F8B09982",
-17345 => x"C0C0BFF9F8B09992",
-17344 => x"C0C0BFF9F8B09999",
-17343 => x"C0C0BFF9F8B099B0",
-17342 => x"C0C0BFF9F8B099A4",
-17341 => x"C0C0BFF9F8B099F9",
-17340 => x"C0C0BFF9F8B099C0",
-17339 => x"C0C0BFF9F8B0B090",
-17338 => x"C0C0BFF9F8B0B080",
-17337 => x"C0C0BFF9F8B0B0F8",
-17336 => x"C0C0BFF9F8B0B082",
-17335 => x"C0C0BFF9F8B0B092",
-17334 => x"C0C0BFF9F8B0B099",
-17333 => x"C0C0BFF9F8B0B0B0",
-17332 => x"C0C0BFF9F8B0B0A4",
-17331 => x"C0C0BFF9F8B0B0F9",
-17330 => x"C0C0BFF9F8B0B0C0",
-17329 => x"C0C0BFF9F8B0A490",
-17328 => x"C0C0BFF9F8B0A480",
-17327 => x"C0C0BFF9F8B0A4F8",
-17326 => x"C0C0BFF9F8B0A482",
-17325 => x"C0C0BFF9F8B0A492",
-17324 => x"C0C0BFF9F8B0A499",
-17323 => x"C0C0BFF9F8B0A4B0",
-17322 => x"C0C0BFF9F8B0A4A4",
-17321 => x"C0C0BFF9F8B0A4F9",
-17320 => x"C0C0BFF9F8B0A4C0",
-17319 => x"C0C0BFF9F8B0F990",
-17318 => x"C0C0BFF9F8B0F980",
-17317 => x"C0C0BFF9F8B0F9F8",
-17316 => x"C0C0BFF9F8B0F982",
-17315 => x"C0C0BFF9F8B0F992",
-17314 => x"C0C0BFF9F8B0F999",
-17313 => x"C0C0BFF9F8B0F9B0",
-17312 => x"C0C0BFF9F8B0F9A4",
-17311 => x"C0C0BFF9F8B0F9F9",
-17310 => x"C0C0BFF9F8B0F9C0",
-17309 => x"C0C0BFF9F8B0C090",
-17308 => x"C0C0BFF9F8B0C080",
-17307 => x"C0C0BFF9F8B0C0F8",
-17306 => x"C0C0BFF9F8B0C082",
-17305 => x"C0C0BFF9F8B0C092",
-17304 => x"C0C0BFF9F8B0C099",
-17303 => x"C0C0BFF9F8B0C0B0",
-17302 => x"C0C0BFF9F8B0C0A4",
-17301 => x"C0C0BFF9F8B0C0F9",
-17300 => x"C0C0BFF9F8B0C0C0",
-17299 => x"C0C0BFF9F8A49090",
-17298 => x"C0C0BFF9F8A49080",
-17297 => x"C0C0BFF9F8A490F8",
-17296 => x"C0C0BFF9F8A49082",
-17295 => x"C0C0BFF9F8A49092",
-17294 => x"C0C0BFF9F8A49099",
-17293 => x"C0C0BFF9F8A490B0",
-17292 => x"C0C0BFF9F8A490A4",
-17291 => x"C0C0BFF9F8A490F9",
-17290 => x"C0C0BFF9F8A490C0",
-17289 => x"C0C0BFF9F8A48090",
-17288 => x"C0C0BFF9F8A48080",
-17287 => x"C0C0BFF9F8A480F8",
-17286 => x"C0C0BFF9F8A48082",
-17285 => x"C0C0BFF9F8A48092",
-17284 => x"C0C0BFF9F8A48099",
-17283 => x"C0C0BFF9F8A480B0",
-17282 => x"C0C0BFF9F8A480A4",
-17281 => x"C0C0BFF9F8A480F9",
-17280 => x"C0C0BFF9F8A480C0",
-17279 => x"C0C0BFF9F8A4F890",
-17278 => x"C0C0BFF9F8A4F880",
-17277 => x"C0C0BFF9F8A4F8F8",
-17276 => x"C0C0BFF9F8A4F882",
-17275 => x"C0C0BFF9F8A4F892",
-17274 => x"C0C0BFF9F8A4F899",
-17273 => x"C0C0BFF9F8A4F8B0",
-17272 => x"C0C0BFF9F8A4F8A4",
-17271 => x"C0C0BFF9F8A4F8F9",
-17270 => x"C0C0BFF9F8A4F8C0",
-17269 => x"C0C0BFF9F8A48290",
-17268 => x"C0C0BFF9F8A48280",
-17267 => x"C0C0BFF9F8A482F8",
-17266 => x"C0C0BFF9F8A48282",
-17265 => x"C0C0BFF9F8A48292",
-17264 => x"C0C0BFF9F8A48299",
-17263 => x"C0C0BFF9F8A482B0",
-17262 => x"C0C0BFF9F8A482A4",
-17261 => x"C0C0BFF9F8A482F9",
-17260 => x"C0C0BFF9F8A482C0",
-17259 => x"C0C0BFF9F8A49290",
-17258 => x"C0C0BFF9F8A49280",
-17257 => x"C0C0BFF9F8A492F8",
-17256 => x"C0C0BFF9F8A49282",
-17255 => x"C0C0BFF9F8A49292",
-17254 => x"C0C0BFF9F8A49299",
-17253 => x"C0C0BFF9F8A492B0",
-17252 => x"C0C0BFF9F8A492A4",
-17251 => x"C0C0BFF9F8A492F9",
-17250 => x"C0C0BFF9F8A492C0",
-17249 => x"C0C0BFF9F8A49990",
-17248 => x"C0C0BFF9F8A49980",
-17247 => x"C0C0BFF9F8A499F8",
-17246 => x"C0C0BFF9F8A49982",
-17245 => x"C0C0BFF9F8A49992",
-17244 => x"C0C0BFF9F8A49999",
-17243 => x"C0C0BFF9F8A499B0",
-17242 => x"C0C0BFF9F8A499A4",
-17241 => x"C0C0BFF9F8A499F9",
-17240 => x"C0C0BFF9F8A499C0",
-17239 => x"C0C0BFF9F8A4B090",
-17238 => x"C0C0BFF9F8A4B080",
-17237 => x"C0C0BFF9F8A4B0F8",
-17236 => x"C0C0BFF9F8A4B082",
-17235 => x"C0C0BFF9F8A4B092",
-17234 => x"C0C0BFF9F8A4B099",
-17233 => x"C0C0BFF9F8A4B0B0",
-17232 => x"C0C0BFF9F8A4B0A4",
-17231 => x"C0C0BFF9F8A4B0F9",
-17230 => x"C0C0BFF9F8A4B0C0",
-17229 => x"C0C0BFF9F8A4A490",
-17228 => x"C0C0BFF9F8A4A480",
-17227 => x"C0C0BFF9F8A4A4F8",
-17226 => x"C0C0BFF9F8A4A482",
-17225 => x"C0C0BFF9F8A4A492",
-17224 => x"C0C0BFF9F8A4A499",
-17223 => x"C0C0BFF9F8A4A4B0",
-17222 => x"C0C0BFF9F8A4A4A4",
-17221 => x"C0C0BFF9F8A4A4F9",
-17220 => x"C0C0BFF9F8A4A4C0",
-17219 => x"C0C0BFF9F8A4F990",
-17218 => x"C0C0BFF9F8A4F980",
-17217 => x"C0C0BFF9F8A4F9F8",
-17216 => x"C0C0BFF9F8A4F982",
-17215 => x"C0C0BFF9F8A4F992",
-17214 => x"C0C0BFF9F8A4F999",
-17213 => x"C0C0BFF9F8A4F9B0",
-17212 => x"C0C0BFF9F8A4F9A4",
-17211 => x"C0C0BFF9F8A4F9F9",
-17210 => x"C0C0BFF9F8A4F9C0",
-17209 => x"C0C0BFF9F8A4C090",
-17208 => x"C0C0BFF9F8A4C080",
-17207 => x"C0C0BFF9F8A4C0F8",
-17206 => x"C0C0BFF9F8A4C082",
-17205 => x"C0C0BFF9F8A4C092",
-17204 => x"C0C0BFF9F8A4C099",
-17203 => x"C0C0BFF9F8A4C0B0",
-17202 => x"C0C0BFF9F8A4C0A4",
-17201 => x"C0C0BFF9F8A4C0F9",
-17200 => x"C0C0BFF9F8A4C0C0",
-17199 => x"C0C0BFF9F8F99090",
-17198 => x"C0C0BFF9F8F99080",
-17197 => x"C0C0BFF9F8F990F8",
-17196 => x"C0C0BFF9F8F99082",
-17195 => x"C0C0BFF9F8F99092",
-17194 => x"C0C0BFF9F8F99099",
-17193 => x"C0C0BFF9F8F990B0",
-17192 => x"C0C0BFF9F8F990A4",
-17191 => x"C0C0BFF9F8F990F9",
-17190 => x"C0C0BFF9F8F990C0",
-17189 => x"C0C0BFF9F8F98090",
-17188 => x"C0C0BFF9F8F98080",
-17187 => x"C0C0BFF9F8F980F8",
-17186 => x"C0C0BFF9F8F98082",
-17185 => x"C0C0BFF9F8F98092",
-17184 => x"C0C0BFF9F8F98099",
-17183 => x"C0C0BFF9F8F980B0",
-17182 => x"C0C0BFF9F8F980A4",
-17181 => x"C0C0BFF9F8F980F9",
-17180 => x"C0C0BFF9F8F980C0",
-17179 => x"C0C0BFF9F8F9F890",
-17178 => x"C0C0BFF9F8F9F880",
-17177 => x"C0C0BFF9F8F9F8F8",
-17176 => x"C0C0BFF9F8F9F882",
-17175 => x"C0C0BFF9F8F9F892",
-17174 => x"C0C0BFF9F8F9F899",
-17173 => x"C0C0BFF9F8F9F8B0",
-17172 => x"C0C0BFF9F8F9F8A4",
-17171 => x"C0C0BFF9F8F9F8F9",
-17170 => x"C0C0BFF9F8F9F8C0",
-17169 => x"C0C0BFF9F8F98290",
-17168 => x"C0C0BFF9F8F98280",
-17167 => x"C0C0BFF9F8F982F8",
-17166 => x"C0C0BFF9F8F98282",
-17165 => x"C0C0BFF9F8F98292",
-17164 => x"C0C0BFF9F8F98299",
-17163 => x"C0C0BFF9F8F982B0",
-17162 => x"C0C0BFF9F8F982A4",
-17161 => x"C0C0BFF9F8F982F9",
-17160 => x"C0C0BFF9F8F982C0",
-17159 => x"C0C0BFF9F8F99290",
-17158 => x"C0C0BFF9F8F99280",
-17157 => x"C0C0BFF9F8F992F8",
-17156 => x"C0C0BFF9F8F99282",
-17155 => x"C0C0BFF9F8F99292",
-17154 => x"C0C0BFF9F8F99299",
-17153 => x"C0C0BFF9F8F992B0",
-17152 => x"C0C0BFF9F8F992A4",
-17151 => x"C0C0BFF9F8F992F9",
-17150 => x"C0C0BFF9F8F992C0",
-17149 => x"C0C0BFF9F8F99990",
-17148 => x"C0C0BFF9F8F99980",
-17147 => x"C0C0BFF9F8F999F8",
-17146 => x"C0C0BFF9F8F99982",
-17145 => x"C0C0BFF9F8F99992",
-17144 => x"C0C0BFF9F8F99999",
-17143 => x"C0C0BFF9F8F999B0",
-17142 => x"C0C0BFF9F8F999A4",
-17141 => x"C0C0BFF9F8F999F9",
-17140 => x"C0C0BFF9F8F999C0",
-17139 => x"C0C0BFF9F8F9B090",
-17138 => x"C0C0BFF9F8F9B080",
-17137 => x"C0C0BFF9F8F9B0F8",
-17136 => x"C0C0BFF9F8F9B082",
-17135 => x"C0C0BFF9F8F9B092",
-17134 => x"C0C0BFF9F8F9B099",
-17133 => x"C0C0BFF9F8F9B0B0",
-17132 => x"C0C0BFF9F8F9B0A4",
-17131 => x"C0C0BFF9F8F9B0F9",
-17130 => x"C0C0BFF9F8F9B0C0",
-17129 => x"C0C0BFF9F8F9A490",
-17128 => x"C0C0BFF9F8F9A480",
-17127 => x"C0C0BFF9F8F9A4F8",
-17126 => x"C0C0BFF9F8F9A482",
-17125 => x"C0C0BFF9F8F9A492",
-17124 => x"C0C0BFF9F8F9A499",
-17123 => x"C0C0BFF9F8F9A4B0",
-17122 => x"C0C0BFF9F8F9A4A4",
-17121 => x"C0C0BFF9F8F9A4F9",
-17120 => x"C0C0BFF9F8F9A4C0",
-17119 => x"C0C0BFF9F8F9F990",
-17118 => x"C0C0BFF9F8F9F980",
-17117 => x"C0C0BFF9F8F9F9F8",
-17116 => x"C0C0BFF9F8F9F982",
-17115 => x"C0C0BFF9F8F9F992",
-17114 => x"C0C0BFF9F8F9F999",
-17113 => x"C0C0BFF9F8F9F9B0",
-17112 => x"C0C0BFF9F8F9F9A4",
-17111 => x"C0C0BFF9F8F9F9F9",
-17110 => x"C0C0BFF9F8F9F9C0",
-17109 => x"C0C0BFF9F8F9C090",
-17108 => x"C0C0BFF9F8F9C080",
-17107 => x"C0C0BFF9F8F9C0F8",
-17106 => x"C0C0BFF9F8F9C082",
-17105 => x"C0C0BFF9F8F9C092",
-17104 => x"C0C0BFF9F8F9C099",
-17103 => x"C0C0BFF9F8F9C0B0",
-17102 => x"C0C0BFF9F8F9C0A4",
-17101 => x"C0C0BFF9F8F9C0F9",
-17100 => x"C0C0BFF9F8F9C0C0",
-17099 => x"C0C0BFF9F8C09090",
-17098 => x"C0C0BFF9F8C09080",
-17097 => x"C0C0BFF9F8C090F8",
-17096 => x"C0C0BFF9F8C09082",
-17095 => x"C0C0BFF9F8C09092",
-17094 => x"C0C0BFF9F8C09099",
-17093 => x"C0C0BFF9F8C090B0",
-17092 => x"C0C0BFF9F8C090A4",
-17091 => x"C0C0BFF9F8C090F9",
-17090 => x"C0C0BFF9F8C090C0",
-17089 => x"C0C0BFF9F8C08090",
-17088 => x"C0C0BFF9F8C08080",
-17087 => x"C0C0BFF9F8C080F8",
-17086 => x"C0C0BFF9F8C08082",
-17085 => x"C0C0BFF9F8C08092",
-17084 => x"C0C0BFF9F8C08099",
-17083 => x"C0C0BFF9F8C080B0",
-17082 => x"C0C0BFF9F8C080A4",
-17081 => x"C0C0BFF9F8C080F9",
-17080 => x"C0C0BFF9F8C080C0",
-17079 => x"C0C0BFF9F8C0F890",
-17078 => x"C0C0BFF9F8C0F880",
-17077 => x"C0C0BFF9F8C0F8F8",
-17076 => x"C0C0BFF9F8C0F882",
-17075 => x"C0C0BFF9F8C0F892",
-17074 => x"C0C0BFF9F8C0F899",
-17073 => x"C0C0BFF9F8C0F8B0",
-17072 => x"C0C0BFF9F8C0F8A4",
-17071 => x"C0C0BFF9F8C0F8F9",
-17070 => x"C0C0BFF9F8C0F8C0",
-17069 => x"C0C0BFF9F8C08290",
-17068 => x"C0C0BFF9F8C08280",
-17067 => x"C0C0BFF9F8C082F8",
-17066 => x"C0C0BFF9F8C08282",
-17065 => x"C0C0BFF9F8C08292",
-17064 => x"C0C0BFF9F8C08299",
-17063 => x"C0C0BFF9F8C082B0",
-17062 => x"C0C0BFF9F8C082A4",
-17061 => x"C0C0BFF9F8C082F9",
-17060 => x"C0C0BFF9F8C082C0",
-17059 => x"C0C0BFF9F8C09290",
-17058 => x"C0C0BFF9F8C09280",
-17057 => x"C0C0BFF9F8C092F8",
-17056 => x"C0C0BFF9F8C09282",
-17055 => x"C0C0BFF9F8C09292",
-17054 => x"C0C0BFF9F8C09299",
-17053 => x"C0C0BFF9F8C092B0",
-17052 => x"C0C0BFF9F8C092A4",
-17051 => x"C0C0BFF9F8C092F9",
-17050 => x"C0C0BFF9F8C092C0",
-17049 => x"C0C0BFF9F8C09990",
-17048 => x"C0C0BFF9F8C09980",
-17047 => x"C0C0BFF9F8C099F8",
-17046 => x"C0C0BFF9F8C09982",
-17045 => x"C0C0BFF9F8C09992",
-17044 => x"C0C0BFF9F8C09999",
-17043 => x"C0C0BFF9F8C099B0",
-17042 => x"C0C0BFF9F8C099A4",
-17041 => x"C0C0BFF9F8C099F9",
-17040 => x"C0C0BFF9F8C099C0",
-17039 => x"C0C0BFF9F8C0B090",
-17038 => x"C0C0BFF9F8C0B080",
-17037 => x"C0C0BFF9F8C0B0F8",
-17036 => x"C0C0BFF9F8C0B082",
-17035 => x"C0C0BFF9F8C0B092",
-17034 => x"C0C0BFF9F8C0B099",
-17033 => x"C0C0BFF9F8C0B0B0",
-17032 => x"C0C0BFF9F8C0B0A4",
-17031 => x"C0C0BFF9F8C0B0F9",
-17030 => x"C0C0BFF9F8C0B0C0",
-17029 => x"C0C0BFF9F8C0A490",
-17028 => x"C0C0BFF9F8C0A480",
-17027 => x"C0C0BFF9F8C0A4F8",
-17026 => x"C0C0BFF9F8C0A482",
-17025 => x"C0C0BFF9F8C0A492",
-17024 => x"C0C0BFF9F8C0A499",
-17023 => x"C0C0BFF9F8C0A4B0",
-17022 => x"C0C0BFF9F8C0A4A4",
-17021 => x"C0C0BFF9F8C0A4F9",
-17020 => x"C0C0BFF9F8C0A4C0",
-17019 => x"C0C0BFF9F8C0F990",
-17018 => x"C0C0BFF9F8C0F980",
-17017 => x"C0C0BFF9F8C0F9F8",
-17016 => x"C0C0BFF9F8C0F982",
-17015 => x"C0C0BFF9F8C0F992",
-17014 => x"C0C0BFF9F8C0F999",
-17013 => x"C0C0BFF9F8C0F9B0",
-17012 => x"C0C0BFF9F8C0F9A4",
-17011 => x"C0C0BFF9F8C0F9F9",
-17010 => x"C0C0BFF9F8C0F9C0",
-17009 => x"C0C0BFF9F8C0C090",
-17008 => x"C0C0BFF9F8C0C080",
-17007 => x"C0C0BFF9F8C0C0F8",
-17006 => x"C0C0BFF9F8C0C082",
-17005 => x"C0C0BFF9F8C0C092",
-17004 => x"C0C0BFF9F8C0C099",
-17003 => x"C0C0BFF9F8C0C0B0",
-17002 => x"C0C0BFF9F8C0C0A4",
-17001 => x"C0C0BFF9F8C0C0F9",
-17000 => x"C0C0BFF9F8C0C0C0",
-16999 => x"C0C0BFF982909090",
-16998 => x"C0C0BFF982909080",
-16997 => x"C0C0BFF9829090F8",
-16996 => x"C0C0BFF982909082",
-16995 => x"C0C0BFF982909092",
-16994 => x"C0C0BFF982909099",
-16993 => x"C0C0BFF9829090B0",
-16992 => x"C0C0BFF9829090A4",
-16991 => x"C0C0BFF9829090F9",
-16990 => x"C0C0BFF9829090C0",
-16989 => x"C0C0BFF982908090",
-16988 => x"C0C0BFF982908080",
-16987 => x"C0C0BFF9829080F8",
-16986 => x"C0C0BFF982908082",
-16985 => x"C0C0BFF982908092",
-16984 => x"C0C0BFF982908099",
-16983 => x"C0C0BFF9829080B0",
-16982 => x"C0C0BFF9829080A4",
-16981 => x"C0C0BFF9829080F9",
-16980 => x"C0C0BFF9829080C0",
-16979 => x"C0C0BFF98290F890",
-16978 => x"C0C0BFF98290F880",
-16977 => x"C0C0BFF98290F8F8",
-16976 => x"C0C0BFF98290F882",
-16975 => x"C0C0BFF98290F892",
-16974 => x"C0C0BFF98290F899",
-16973 => x"C0C0BFF98290F8B0",
-16972 => x"C0C0BFF98290F8A4",
-16971 => x"C0C0BFF98290F8F9",
-16970 => x"C0C0BFF98290F8C0",
-16969 => x"C0C0BFF982908290",
-16968 => x"C0C0BFF982908280",
-16967 => x"C0C0BFF9829082F8",
-16966 => x"C0C0BFF982908282",
-16965 => x"C0C0BFF982908292",
-16964 => x"C0C0BFF982908299",
-16963 => x"C0C0BFF9829082B0",
-16962 => x"C0C0BFF9829082A4",
-16961 => x"C0C0BFF9829082F9",
-16960 => x"C0C0BFF9829082C0",
-16959 => x"C0C0BFF982909290",
-16958 => x"C0C0BFF982909280",
-16957 => x"C0C0BFF9829092F8",
-16956 => x"C0C0BFF982909282",
-16955 => x"C0C0BFF982909292",
-16954 => x"C0C0BFF982909299",
-16953 => x"C0C0BFF9829092B0",
-16952 => x"C0C0BFF9829092A4",
-16951 => x"C0C0BFF9829092F9",
-16950 => x"C0C0BFF9829092C0",
-16949 => x"C0C0BFF982909990",
-16948 => x"C0C0BFF982909980",
-16947 => x"C0C0BFF9829099F8",
-16946 => x"C0C0BFF982909982",
-16945 => x"C0C0BFF982909992",
-16944 => x"C0C0BFF982909999",
-16943 => x"C0C0BFF9829099B0",
-16942 => x"C0C0BFF9829099A4",
-16941 => x"C0C0BFF9829099F9",
-16940 => x"C0C0BFF9829099C0",
-16939 => x"C0C0BFF98290B090",
-16938 => x"C0C0BFF98290B080",
-16937 => x"C0C0BFF98290B0F8",
-16936 => x"C0C0BFF98290B082",
-16935 => x"C0C0BFF98290B092",
-16934 => x"C0C0BFF98290B099",
-16933 => x"C0C0BFF98290B0B0",
-16932 => x"C0C0BFF98290B0A4",
-16931 => x"C0C0BFF98290B0F9",
-16930 => x"C0C0BFF98290B0C0",
-16929 => x"C0C0BFF98290A490",
-16928 => x"C0C0BFF98290A480",
-16927 => x"C0C0BFF98290A4F8",
-16926 => x"C0C0BFF98290A482",
-16925 => x"C0C0BFF98290A492",
-16924 => x"C0C0BFF98290A499",
-16923 => x"C0C0BFF98290A4B0",
-16922 => x"C0C0BFF98290A4A4",
-16921 => x"C0C0BFF98290A4F9",
-16920 => x"C0C0BFF98290A4C0",
-16919 => x"C0C0BFF98290F990",
-16918 => x"C0C0BFF98290F980",
-16917 => x"C0C0BFF98290F9F8",
-16916 => x"C0C0BFF98290F982",
-16915 => x"C0C0BFF98290F992",
-16914 => x"C0C0BFF98290F999",
-16913 => x"C0C0BFF98290F9B0",
-16912 => x"C0C0BFF98290F9A4",
-16911 => x"C0C0BFF98290F9F9",
-16910 => x"C0C0BFF98290F9C0",
-16909 => x"C0C0BFF98290C090",
-16908 => x"C0C0BFF98290C080",
-16907 => x"C0C0BFF98290C0F8",
-16906 => x"C0C0BFF98290C082",
-16905 => x"C0C0BFF98290C092",
-16904 => x"C0C0BFF98290C099",
-16903 => x"C0C0BFF98290C0B0",
-16902 => x"C0C0BFF98290C0A4",
-16901 => x"C0C0BFF98290C0F9",
-16900 => x"C0C0BFF98290C0C0",
-16899 => x"C0C0BFF982809090",
-16898 => x"C0C0BFF982809080",
-16897 => x"C0C0BFF9828090F8",
-16896 => x"C0C0BFF982809082",
-16895 => x"C0C0BFF982809092",
-16894 => x"C0C0BFF982809099",
-16893 => x"C0C0BFF9828090B0",
-16892 => x"C0C0BFF9828090A4",
-16891 => x"C0C0BFF9828090F9",
-16890 => x"C0C0BFF9828090C0",
-16889 => x"C0C0BFF982808090",
-16888 => x"C0C0BFF982808080",
-16887 => x"C0C0BFF9828080F8",
-16886 => x"C0C0BFF982808082",
-16885 => x"C0C0BFF982808092",
-16884 => x"C0C0BFF982808099",
-16883 => x"C0C0BFF9828080B0",
-16882 => x"C0C0BFF9828080A4",
-16881 => x"C0C0BFF9828080F9",
-16880 => x"C0C0BFF9828080C0",
-16879 => x"C0C0BFF98280F890",
-16878 => x"C0C0BFF98280F880",
-16877 => x"C0C0BFF98280F8F8",
-16876 => x"C0C0BFF98280F882",
-16875 => x"C0C0BFF98280F892",
-16874 => x"C0C0BFF98280F899",
-16873 => x"C0C0BFF98280F8B0",
-16872 => x"C0C0BFF98280F8A4",
-16871 => x"C0C0BFF98280F8F9",
-16870 => x"C0C0BFF98280F8C0",
-16869 => x"C0C0BFF982808290",
-16868 => x"C0C0BFF982808280",
-16867 => x"C0C0BFF9828082F8",
-16866 => x"C0C0BFF982808282",
-16865 => x"C0C0BFF982808292",
-16864 => x"C0C0BFF982808299",
-16863 => x"C0C0BFF9828082B0",
-16862 => x"C0C0BFF9828082A4",
-16861 => x"C0C0BFF9828082F9",
-16860 => x"C0C0BFF9828082C0",
-16859 => x"C0C0BFF982809290",
-16858 => x"C0C0BFF982809280",
-16857 => x"C0C0BFF9828092F8",
-16856 => x"C0C0BFF982809282",
-16855 => x"C0C0BFF982809292",
-16854 => x"C0C0BFF982809299",
-16853 => x"C0C0BFF9828092B0",
-16852 => x"C0C0BFF9828092A4",
-16851 => x"C0C0BFF9828092F9",
-16850 => x"C0C0BFF9828092C0",
-16849 => x"C0C0BFF982809990",
-16848 => x"C0C0BFF982809980",
-16847 => x"C0C0BFF9828099F8",
-16846 => x"C0C0BFF982809982",
-16845 => x"C0C0BFF982809992",
-16844 => x"C0C0BFF982809999",
-16843 => x"C0C0BFF9828099B0",
-16842 => x"C0C0BFF9828099A4",
-16841 => x"C0C0BFF9828099F9",
-16840 => x"C0C0BFF9828099C0",
-16839 => x"C0C0BFF98280B090",
-16838 => x"C0C0BFF98280B080",
-16837 => x"C0C0BFF98280B0F8",
-16836 => x"C0C0BFF98280B082",
-16835 => x"C0C0BFF98280B092",
-16834 => x"C0C0BFF98280B099",
-16833 => x"C0C0BFF98280B0B0",
-16832 => x"C0C0BFF98280B0A4",
-16831 => x"C0C0BFF98280B0F9",
-16830 => x"C0C0BFF98280B0C0",
-16829 => x"C0C0BFF98280A490",
-16828 => x"C0C0BFF98280A480",
-16827 => x"C0C0BFF98280A4F8",
-16826 => x"C0C0BFF98280A482",
-16825 => x"C0C0BFF98280A492",
-16824 => x"C0C0BFF98280A499",
-16823 => x"C0C0BFF98280A4B0",
-16822 => x"C0C0BFF98280A4A4",
-16821 => x"C0C0BFF98280A4F9",
-16820 => x"C0C0BFF98280A4C0",
-16819 => x"C0C0BFF98280F990",
-16818 => x"C0C0BFF98280F980",
-16817 => x"C0C0BFF98280F9F8",
-16816 => x"C0C0BFF98280F982",
-16815 => x"C0C0BFF98280F992",
-16814 => x"C0C0BFF98280F999",
-16813 => x"C0C0BFF98280F9B0",
-16812 => x"C0C0BFF98280F9A4",
-16811 => x"C0C0BFF98280F9F9",
-16810 => x"C0C0BFF98280F9C0",
-16809 => x"C0C0BFF98280C090",
-16808 => x"C0C0BFF98280C080",
-16807 => x"C0C0BFF98280C0F8",
-16806 => x"C0C0BFF98280C082",
-16805 => x"C0C0BFF98280C092",
-16804 => x"C0C0BFF98280C099",
-16803 => x"C0C0BFF98280C0B0",
-16802 => x"C0C0BFF98280C0A4",
-16801 => x"C0C0BFF98280C0F9",
-16800 => x"C0C0BFF98280C0C0",
-16799 => x"C0C0BFF982F89090",
-16798 => x"C0C0BFF982F89080",
-16797 => x"C0C0BFF982F890F8",
-16796 => x"C0C0BFF982F89082",
-16795 => x"C0C0BFF982F89092",
-16794 => x"C0C0BFF982F89099",
-16793 => x"C0C0BFF982F890B0",
-16792 => x"C0C0BFF982F890A4",
-16791 => x"C0C0BFF982F890F9",
-16790 => x"C0C0BFF982F890C0",
-16789 => x"C0C0BFF982F88090",
-16788 => x"C0C0BFF982F88080",
-16787 => x"C0C0BFF982F880F8",
-16786 => x"C0C0BFF982F88082",
-16785 => x"C0C0BFF982F88092",
-16784 => x"C0C0BFF982F88099",
-16783 => x"C0C0BFF982F880B0",
-16782 => x"C0C0BFF982F880A4",
-16781 => x"C0C0BFF982F880F9",
-16780 => x"C0C0BFF982F880C0",
-16779 => x"C0C0BFF982F8F890",
-16778 => x"C0C0BFF982F8F880",
-16777 => x"C0C0BFF982F8F8F8",
-16776 => x"C0C0BFF982F8F882",
-16775 => x"C0C0BFF982F8F892",
-16774 => x"C0C0BFF982F8F899",
-16773 => x"C0C0BFF982F8F8B0",
-16772 => x"C0C0BFF982F8F8A4",
-16771 => x"C0C0BFF982F8F8F9",
-16770 => x"C0C0BFF982F8F8C0",
-16769 => x"C0C0BFF982F88290",
-16768 => x"C0C0BFF982F88280",
-16767 => x"C0C0BFF982F882F8",
-16766 => x"C0C0BFF982F88282",
-16765 => x"C0C0BFF982F88292",
-16764 => x"C0C0BFF982F88299",
-16763 => x"C0C0BFF982F882B0",
-16762 => x"C0C0BFF982F882A4",
-16761 => x"C0C0BFF982F882F9",
-16760 => x"C0C0BFF982F882C0",
-16759 => x"C0C0BFF982F89290",
-16758 => x"C0C0BFF982F89280",
-16757 => x"C0C0BFF982F892F8",
-16756 => x"C0C0BFF982F89282",
-16755 => x"C0C0BFF982F89292",
-16754 => x"C0C0BFF982F89299",
-16753 => x"C0C0BFF982F892B0",
-16752 => x"C0C0BFF982F892A4",
-16751 => x"C0C0BFF982F892F9",
-16750 => x"C0C0BFF982F892C0",
-16749 => x"C0C0BFF982F89990",
-16748 => x"C0C0BFF982F89980",
-16747 => x"C0C0BFF982F899F8",
-16746 => x"C0C0BFF982F89982",
-16745 => x"C0C0BFF982F89992",
-16744 => x"C0C0BFF982F89999",
-16743 => x"C0C0BFF982F899B0",
-16742 => x"C0C0BFF982F899A4",
-16741 => x"C0C0BFF982F899F9",
-16740 => x"C0C0BFF982F899C0",
-16739 => x"C0C0BFF982F8B090",
-16738 => x"C0C0BFF982F8B080",
-16737 => x"C0C0BFF982F8B0F8",
-16736 => x"C0C0BFF982F8B082",
-16735 => x"C0C0BFF982F8B092",
-16734 => x"C0C0BFF982F8B099",
-16733 => x"C0C0BFF982F8B0B0",
-16732 => x"C0C0BFF982F8B0A4",
-16731 => x"C0C0BFF982F8B0F9",
-16730 => x"C0C0BFF982F8B0C0",
-16729 => x"C0C0BFF982F8A490",
-16728 => x"C0C0BFF982F8A480",
-16727 => x"C0C0BFF982F8A4F8",
-16726 => x"C0C0BFF982F8A482",
-16725 => x"C0C0BFF982F8A492",
-16724 => x"C0C0BFF982F8A499",
-16723 => x"C0C0BFF982F8A4B0",
-16722 => x"C0C0BFF982F8A4A4",
-16721 => x"C0C0BFF982F8A4F9",
-16720 => x"C0C0BFF982F8A4C0",
-16719 => x"C0C0BFF982F8F990",
-16718 => x"C0C0BFF982F8F980",
-16717 => x"C0C0BFF982F8F9F8",
-16716 => x"C0C0BFF982F8F982",
-16715 => x"C0C0BFF982F8F992",
-16714 => x"C0C0BFF982F8F999",
-16713 => x"C0C0BFF982F8F9B0",
-16712 => x"C0C0BFF982F8F9A4",
-16711 => x"C0C0BFF982F8F9F9",
-16710 => x"C0C0BFF982F8F9C0",
-16709 => x"C0C0BFF982F8C090",
-16708 => x"C0C0BFF982F8C080",
-16707 => x"C0C0BFF982F8C0F8",
-16706 => x"C0C0BFF982F8C082",
-16705 => x"C0C0BFF982F8C092",
-16704 => x"C0C0BFF982F8C099",
-16703 => x"C0C0BFF982F8C0B0",
-16702 => x"C0C0BFF982F8C0A4",
-16701 => x"C0C0BFF982F8C0F9",
-16700 => x"C0C0BFF982F8C0C0",
-16699 => x"C0C0BFF982829090",
-16698 => x"C0C0BFF982829080",
-16697 => x"C0C0BFF9828290F8",
-16696 => x"C0C0BFF982829082",
-16695 => x"C0C0BFF982829092",
-16694 => x"C0C0BFF982829099",
-16693 => x"C0C0BFF9828290B0",
-16692 => x"C0C0BFF9828290A4",
-16691 => x"C0C0BFF9828290F9",
-16690 => x"C0C0BFF9828290C0",
-16689 => x"C0C0BFF982828090",
-16688 => x"C0C0BFF982828080",
-16687 => x"C0C0BFF9828280F8",
-16686 => x"C0C0BFF982828082",
-16685 => x"C0C0BFF982828092",
-16684 => x"C0C0BFF982828099",
-16683 => x"C0C0BFF9828280B0",
-16682 => x"C0C0BFF9828280A4",
-16681 => x"C0C0BFF9828280F9",
-16680 => x"C0C0BFF9828280C0",
-16679 => x"C0C0BFF98282F890",
-16678 => x"C0C0BFF98282F880",
-16677 => x"C0C0BFF98282F8F8",
-16676 => x"C0C0BFF98282F882",
-16675 => x"C0C0BFF98282F892",
-16674 => x"C0C0BFF98282F899",
-16673 => x"C0C0BFF98282F8B0",
-16672 => x"C0C0BFF98282F8A4",
-16671 => x"C0C0BFF98282F8F9",
-16670 => x"C0C0BFF98282F8C0",
-16669 => x"C0C0BFF982828290",
-16668 => x"C0C0BFF982828280",
-16667 => x"C0C0BFF9828282F8",
-16666 => x"C0C0BFF982828282",
-16665 => x"C0C0BFF982828292",
-16664 => x"C0C0BFF982828299",
-16663 => x"C0C0BFF9828282B0",
-16662 => x"C0C0BFF9828282A4",
-16661 => x"C0C0BFF9828282F9",
-16660 => x"C0C0BFF9828282C0",
-16659 => x"C0C0BFF982829290",
-16658 => x"C0C0BFF982829280",
-16657 => x"C0C0BFF9828292F8",
-16656 => x"C0C0BFF982829282",
-16655 => x"C0C0BFF982829292",
-16654 => x"C0C0BFF982829299",
-16653 => x"C0C0BFF9828292B0",
-16652 => x"C0C0BFF9828292A4",
-16651 => x"C0C0BFF9828292F9",
-16650 => x"C0C0BFF9828292C0",
-16649 => x"C0C0BFF982829990",
-16648 => x"C0C0BFF982829980",
-16647 => x"C0C0BFF9828299F8",
-16646 => x"C0C0BFF982829982",
-16645 => x"C0C0BFF982829992",
-16644 => x"C0C0BFF982829999",
-16643 => x"C0C0BFF9828299B0",
-16642 => x"C0C0BFF9828299A4",
-16641 => x"C0C0BFF9828299F9",
-16640 => x"C0C0BFF9828299C0",
-16639 => x"C0C0BFF98282B090",
-16638 => x"C0C0BFF98282B080",
-16637 => x"C0C0BFF98282B0F8",
-16636 => x"C0C0BFF98282B082",
-16635 => x"C0C0BFF98282B092",
-16634 => x"C0C0BFF98282B099",
-16633 => x"C0C0BFF98282B0B0",
-16632 => x"C0C0BFF98282B0A4",
-16631 => x"C0C0BFF98282B0F9",
-16630 => x"C0C0BFF98282B0C0",
-16629 => x"C0C0BFF98282A490",
-16628 => x"C0C0BFF98282A480",
-16627 => x"C0C0BFF98282A4F8",
-16626 => x"C0C0BFF98282A482",
-16625 => x"C0C0BFF98282A492",
-16624 => x"C0C0BFF98282A499",
-16623 => x"C0C0BFF98282A4B0",
-16622 => x"C0C0BFF98282A4A4",
-16621 => x"C0C0BFF98282A4F9",
-16620 => x"C0C0BFF98282A4C0",
-16619 => x"C0C0BFF98282F990",
-16618 => x"C0C0BFF98282F980",
-16617 => x"C0C0BFF98282F9F8",
-16616 => x"C0C0BFF98282F982",
-16615 => x"C0C0BFF98282F992",
-16614 => x"C0C0BFF98282F999",
-16613 => x"C0C0BFF98282F9B0",
-16612 => x"C0C0BFF98282F9A4",
-16611 => x"C0C0BFF98282F9F9",
-16610 => x"C0C0BFF98282F9C0",
-16609 => x"C0C0BFF98282C090",
-16608 => x"C0C0BFF98282C080",
-16607 => x"C0C0BFF98282C0F8",
-16606 => x"C0C0BFF98282C082",
-16605 => x"C0C0BFF98282C092",
-16604 => x"C0C0BFF98282C099",
-16603 => x"C0C0BFF98282C0B0",
-16602 => x"C0C0BFF98282C0A4",
-16601 => x"C0C0BFF98282C0F9",
-16600 => x"C0C0BFF98282C0C0",
-16599 => x"C0C0BFF982929090",
-16598 => x"C0C0BFF982929080",
-16597 => x"C0C0BFF9829290F8",
-16596 => x"C0C0BFF982929082",
-16595 => x"C0C0BFF982929092",
-16594 => x"C0C0BFF982929099",
-16593 => x"C0C0BFF9829290B0",
-16592 => x"C0C0BFF9829290A4",
-16591 => x"C0C0BFF9829290F9",
-16590 => x"C0C0BFF9829290C0",
-16589 => x"C0C0BFF982928090",
-16588 => x"C0C0BFF982928080",
-16587 => x"C0C0BFF9829280F8",
-16586 => x"C0C0BFF982928082",
-16585 => x"C0C0BFF982928092",
-16584 => x"C0C0BFF982928099",
-16583 => x"C0C0BFF9829280B0",
-16582 => x"C0C0BFF9829280A4",
-16581 => x"C0C0BFF9829280F9",
-16580 => x"C0C0BFF9829280C0",
-16579 => x"C0C0BFF98292F890",
-16578 => x"C0C0BFF98292F880",
-16577 => x"C0C0BFF98292F8F8",
-16576 => x"C0C0BFF98292F882",
-16575 => x"C0C0BFF98292F892",
-16574 => x"C0C0BFF98292F899",
-16573 => x"C0C0BFF98292F8B0",
-16572 => x"C0C0BFF98292F8A4",
-16571 => x"C0C0BFF98292F8F9",
-16570 => x"C0C0BFF98292F8C0",
-16569 => x"C0C0BFF982928290",
-16568 => x"C0C0BFF982928280",
-16567 => x"C0C0BFF9829282F8",
-16566 => x"C0C0BFF982928282",
-16565 => x"C0C0BFF982928292",
-16564 => x"C0C0BFF982928299",
-16563 => x"C0C0BFF9829282B0",
-16562 => x"C0C0BFF9829282A4",
-16561 => x"C0C0BFF9829282F9",
-16560 => x"C0C0BFF9829282C0",
-16559 => x"C0C0BFF982929290",
-16558 => x"C0C0BFF982929280",
-16557 => x"C0C0BFF9829292F8",
-16556 => x"C0C0BFF982929282",
-16555 => x"C0C0BFF982929292",
-16554 => x"C0C0BFF982929299",
-16553 => x"C0C0BFF9829292B0",
-16552 => x"C0C0BFF9829292A4",
-16551 => x"C0C0BFF9829292F9",
-16550 => x"C0C0BFF9829292C0",
-16549 => x"C0C0BFF982929990",
-16548 => x"C0C0BFF982929980",
-16547 => x"C0C0BFF9829299F8",
-16546 => x"C0C0BFF982929982",
-16545 => x"C0C0BFF982929992",
-16544 => x"C0C0BFF982929999",
-16543 => x"C0C0BFF9829299B0",
-16542 => x"C0C0BFF9829299A4",
-16541 => x"C0C0BFF9829299F9",
-16540 => x"C0C0BFF9829299C0",
-16539 => x"C0C0BFF98292B090",
-16538 => x"C0C0BFF98292B080",
-16537 => x"C0C0BFF98292B0F8",
-16536 => x"C0C0BFF98292B082",
-16535 => x"C0C0BFF98292B092",
-16534 => x"C0C0BFF98292B099",
-16533 => x"C0C0BFF98292B0B0",
-16532 => x"C0C0BFF98292B0A4",
-16531 => x"C0C0BFF98292B0F9",
-16530 => x"C0C0BFF98292B0C0",
-16529 => x"C0C0BFF98292A490",
-16528 => x"C0C0BFF98292A480",
-16527 => x"C0C0BFF98292A4F8",
-16526 => x"C0C0BFF98292A482",
-16525 => x"C0C0BFF98292A492",
-16524 => x"C0C0BFF98292A499",
-16523 => x"C0C0BFF98292A4B0",
-16522 => x"C0C0BFF98292A4A4",
-16521 => x"C0C0BFF98292A4F9",
-16520 => x"C0C0BFF98292A4C0",
-16519 => x"C0C0BFF98292F990",
-16518 => x"C0C0BFF98292F980",
-16517 => x"C0C0BFF98292F9F8",
-16516 => x"C0C0BFF98292F982",
-16515 => x"C0C0BFF98292F992",
-16514 => x"C0C0BFF98292F999",
-16513 => x"C0C0BFF98292F9B0",
-16512 => x"C0C0BFF98292F9A4",
-16511 => x"C0C0BFF98292F9F9",
-16510 => x"C0C0BFF98292F9C0",
-16509 => x"C0C0BFF98292C090",
-16508 => x"C0C0BFF98292C080",
-16507 => x"C0C0BFF98292C0F8",
-16506 => x"C0C0BFF98292C082",
-16505 => x"C0C0BFF98292C092",
-16504 => x"C0C0BFF98292C099",
-16503 => x"C0C0BFF98292C0B0",
-16502 => x"C0C0BFF98292C0A4",
-16501 => x"C0C0BFF98292C0F9",
-16500 => x"C0C0BFF98292C0C0",
-16499 => x"C0C0BFF982999090",
-16498 => x"C0C0BFF982999080",
-16497 => x"C0C0BFF9829990F8",
-16496 => x"C0C0BFF982999082",
-16495 => x"C0C0BFF982999092",
-16494 => x"C0C0BFF982999099",
-16493 => x"C0C0BFF9829990B0",
-16492 => x"C0C0BFF9829990A4",
-16491 => x"C0C0BFF9829990F9",
-16490 => x"C0C0BFF9829990C0",
-16489 => x"C0C0BFF982998090",
-16488 => x"C0C0BFF982998080",
-16487 => x"C0C0BFF9829980F8",
-16486 => x"C0C0BFF982998082",
-16485 => x"C0C0BFF982998092",
-16484 => x"C0C0BFF982998099",
-16483 => x"C0C0BFF9829980B0",
-16482 => x"C0C0BFF9829980A4",
-16481 => x"C0C0BFF9829980F9",
-16480 => x"C0C0BFF9829980C0",
-16479 => x"C0C0BFF98299F890",
-16478 => x"C0C0BFF98299F880",
-16477 => x"C0C0BFF98299F8F8",
-16476 => x"C0C0BFF98299F882",
-16475 => x"C0C0BFF98299F892",
-16474 => x"C0C0BFF98299F899",
-16473 => x"C0C0BFF98299F8B0",
-16472 => x"C0C0BFF98299F8A4",
-16471 => x"C0C0BFF98299F8F9",
-16470 => x"C0C0BFF98299F8C0",
-16469 => x"C0C0BFF982998290",
-16468 => x"C0C0BFF982998280",
-16467 => x"C0C0BFF9829982F8",
-16466 => x"C0C0BFF982998282",
-16465 => x"C0C0BFF982998292",
-16464 => x"C0C0BFF982998299",
-16463 => x"C0C0BFF9829982B0",
-16462 => x"C0C0BFF9829982A4",
-16461 => x"C0C0BFF9829982F9",
-16460 => x"C0C0BFF9829982C0",
-16459 => x"C0C0BFF982999290",
-16458 => x"C0C0BFF982999280",
-16457 => x"C0C0BFF9829992F8",
-16456 => x"C0C0BFF982999282",
-16455 => x"C0C0BFF982999292",
-16454 => x"C0C0BFF982999299",
-16453 => x"C0C0BFF9829992B0",
-16452 => x"C0C0BFF9829992A4",
-16451 => x"C0C0BFF9829992F9",
-16450 => x"C0C0BFF9829992C0",
-16449 => x"C0C0BFF982999990",
-16448 => x"C0C0BFF982999980",
-16447 => x"C0C0BFF9829999F8",
-16446 => x"C0C0BFF982999982",
-16445 => x"C0C0BFF982999992",
-16444 => x"C0C0BFF982999999",
-16443 => x"C0C0BFF9829999B0",
-16442 => x"C0C0BFF9829999A4",
-16441 => x"C0C0BFF9829999F9",
-16440 => x"C0C0BFF9829999C0",
-16439 => x"C0C0BFF98299B090",
-16438 => x"C0C0BFF98299B080",
-16437 => x"C0C0BFF98299B0F8",
-16436 => x"C0C0BFF98299B082",
-16435 => x"C0C0BFF98299B092",
-16434 => x"C0C0BFF98299B099",
-16433 => x"C0C0BFF98299B0B0",
-16432 => x"C0C0BFF98299B0A4",
-16431 => x"C0C0BFF98299B0F9",
-16430 => x"C0C0BFF98299B0C0",
-16429 => x"C0C0BFF98299A490",
-16428 => x"C0C0BFF98299A480",
-16427 => x"C0C0BFF98299A4F8",
-16426 => x"C0C0BFF98299A482",
-16425 => x"C0C0BFF98299A492",
-16424 => x"C0C0BFF98299A499",
-16423 => x"C0C0BFF98299A4B0",
-16422 => x"C0C0BFF98299A4A4",
-16421 => x"C0C0BFF98299A4F9",
-16420 => x"C0C0BFF98299A4C0",
-16419 => x"C0C0BFF98299F990",
-16418 => x"C0C0BFF98299F980",
-16417 => x"C0C0BFF98299F9F8",
-16416 => x"C0C0BFF98299F982",
-16415 => x"C0C0BFF98299F992",
-16414 => x"C0C0BFF98299F999",
-16413 => x"C0C0BFF98299F9B0",
-16412 => x"C0C0BFF98299F9A4",
-16411 => x"C0C0BFF98299F9F9",
-16410 => x"C0C0BFF98299F9C0",
-16409 => x"C0C0BFF98299C090",
-16408 => x"C0C0BFF98299C080",
-16407 => x"C0C0BFF98299C0F8",
-16406 => x"C0C0BFF98299C082",
-16405 => x"C0C0BFF98299C092",
-16404 => x"C0C0BFF98299C099",
-16403 => x"C0C0BFF98299C0B0",
-16402 => x"C0C0BFF98299C0A4",
-16401 => x"C0C0BFF98299C0F9",
-16400 => x"C0C0BFF98299C0C0",
-16399 => x"C0C0BFF982B09090",
-16398 => x"C0C0BFF982B09080",
-16397 => x"C0C0BFF982B090F8",
-16396 => x"C0C0BFF982B09082",
-16395 => x"C0C0BFF982B09092",
-16394 => x"C0C0BFF982B09099",
-16393 => x"C0C0BFF982B090B0",
-16392 => x"C0C0BFF982B090A4",
-16391 => x"C0C0BFF982B090F9",
-16390 => x"C0C0BFF982B090C0",
-16389 => x"C0C0BFF982B08090",
-16388 => x"C0C0BFF982B08080",
-16387 => x"C0C0BFF982B080F8",
-16386 => x"C0C0BFF982B08082",
-16385 => x"C0C0BFF982B08092",
-16384 => x"C0C0BFF982B08099",
-16383 => x"C0C0BFF982B080B0",
-16382 => x"C0C0BFF982B080A4",
-16381 => x"C0C0BFF982B080F9",
-16380 => x"C0C0BFF982B080C0",
-16379 => x"C0C0BFF982B0F890",
-16378 => x"C0C0BFF982B0F880",
-16377 => x"C0C0BFF982B0F8F8",
-16376 => x"C0C0BFF982B0F882",
-16375 => x"C0C0BFF982B0F892",
-16374 => x"C0C0BFF982B0F899",
-16373 => x"C0C0BFF982B0F8B0",
-16372 => x"C0C0BFF982B0F8A4",
-16371 => x"C0C0BFF982B0F8F9",
-16370 => x"C0C0BFF982B0F8C0",
-16369 => x"C0C0BFF982B08290",
-16368 => x"C0C0BFF982B08280",
-16367 => x"C0C0BFF982B082F8",
-16366 => x"C0C0BFF982B08282",
-16365 => x"C0C0BFF982B08292",
-16364 => x"C0C0BFF982B08299",
-16363 => x"C0C0BFF982B082B0",
-16362 => x"C0C0BFF982B082A4",
-16361 => x"C0C0BFF982B082F9",
-16360 => x"C0C0BFF982B082C0",
-16359 => x"C0C0BFF982B09290",
-16358 => x"C0C0BFF982B09280",
-16357 => x"C0C0BFF982B092F8",
-16356 => x"C0C0BFF982B09282",
-16355 => x"C0C0BFF982B09292",
-16354 => x"C0C0BFF982B09299",
-16353 => x"C0C0BFF982B092B0",
-16352 => x"C0C0BFF982B092A4",
-16351 => x"C0C0BFF982B092F9",
-16350 => x"C0C0BFF982B092C0",
-16349 => x"C0C0BFF982B09990",
-16348 => x"C0C0BFF982B09980",
-16347 => x"C0C0BFF982B099F8",
-16346 => x"C0C0BFF982B09982",
-16345 => x"C0C0BFF982B09992",
-16344 => x"C0C0BFF982B09999",
-16343 => x"C0C0BFF982B099B0",
-16342 => x"C0C0BFF982B099A4",
-16341 => x"C0C0BFF982B099F9",
-16340 => x"C0C0BFF982B099C0",
-16339 => x"C0C0BFF982B0B090",
-16338 => x"C0C0BFF982B0B080",
-16337 => x"C0C0BFF982B0B0F8",
-16336 => x"C0C0BFF982B0B082",
-16335 => x"C0C0BFF982B0B092",
-16334 => x"C0C0BFF982B0B099",
-16333 => x"C0C0BFF982B0B0B0",
-16332 => x"C0C0BFF982B0B0A4",
-16331 => x"C0C0BFF982B0B0F9",
-16330 => x"C0C0BFF982B0B0C0",
-16329 => x"C0C0BFF982B0A490",
-16328 => x"C0C0BFF982B0A480",
-16327 => x"C0C0BFF982B0A4F8",
-16326 => x"C0C0BFF982B0A482",
-16325 => x"C0C0BFF982B0A492",
-16324 => x"C0C0BFF982B0A499",
-16323 => x"C0C0BFF982B0A4B0",
-16322 => x"C0C0BFF982B0A4A4",
-16321 => x"C0C0BFF982B0A4F9",
-16320 => x"C0C0BFF982B0A4C0",
-16319 => x"C0C0BFF982B0F990",
-16318 => x"C0C0BFF982B0F980",
-16317 => x"C0C0BFF982B0F9F8",
-16316 => x"C0C0BFF982B0F982",
-16315 => x"C0C0BFF982B0F992",
-16314 => x"C0C0BFF982B0F999",
-16313 => x"C0C0BFF982B0F9B0",
-16312 => x"C0C0BFF982B0F9A4",
-16311 => x"C0C0BFF982B0F9F9",
-16310 => x"C0C0BFF982B0F9C0",
-16309 => x"C0C0BFF982B0C090",
-16308 => x"C0C0BFF982B0C080",
-16307 => x"C0C0BFF982B0C0F8",
-16306 => x"C0C0BFF982B0C082",
-16305 => x"C0C0BFF982B0C092",
-16304 => x"C0C0BFF982B0C099",
-16303 => x"C0C0BFF982B0C0B0",
-16302 => x"C0C0BFF982B0C0A4",
-16301 => x"C0C0BFF982B0C0F9",
-16300 => x"C0C0BFF982B0C0C0",
-16299 => x"C0C0BFF982A49090",
-16298 => x"C0C0BFF982A49080",
-16297 => x"C0C0BFF982A490F8",
-16296 => x"C0C0BFF982A49082",
-16295 => x"C0C0BFF982A49092",
-16294 => x"C0C0BFF982A49099",
-16293 => x"C0C0BFF982A490B0",
-16292 => x"C0C0BFF982A490A4",
-16291 => x"C0C0BFF982A490F9",
-16290 => x"C0C0BFF982A490C0",
-16289 => x"C0C0BFF982A48090",
-16288 => x"C0C0BFF982A48080",
-16287 => x"C0C0BFF982A480F8",
-16286 => x"C0C0BFF982A48082",
-16285 => x"C0C0BFF982A48092",
-16284 => x"C0C0BFF982A48099",
-16283 => x"C0C0BFF982A480B0",
-16282 => x"C0C0BFF982A480A4",
-16281 => x"C0C0BFF982A480F9",
-16280 => x"C0C0BFF982A480C0",
-16279 => x"C0C0BFF982A4F890",
-16278 => x"C0C0BFF982A4F880",
-16277 => x"C0C0BFF982A4F8F8",
-16276 => x"C0C0BFF982A4F882",
-16275 => x"C0C0BFF982A4F892",
-16274 => x"C0C0BFF982A4F899",
-16273 => x"C0C0BFF982A4F8B0",
-16272 => x"C0C0BFF982A4F8A4",
-16271 => x"C0C0BFF982A4F8F9",
-16270 => x"C0C0BFF982A4F8C0",
-16269 => x"C0C0BFF982A48290",
-16268 => x"C0C0BFF982A48280",
-16267 => x"C0C0BFF982A482F8",
-16266 => x"C0C0BFF982A48282",
-16265 => x"C0C0BFF982A48292",
-16264 => x"C0C0BFF982A48299",
-16263 => x"C0C0BFF982A482B0",
-16262 => x"C0C0BFF982A482A4",
-16261 => x"C0C0BFF982A482F9",
-16260 => x"C0C0BFF982A482C0",
-16259 => x"C0C0BFF982A49290",
-16258 => x"C0C0BFF982A49280",
-16257 => x"C0C0BFF982A492F8",
-16256 => x"C0C0BFF982A49282",
-16255 => x"C0C0BFF982A49292",
-16254 => x"C0C0BFF982A49299",
-16253 => x"C0C0BFF982A492B0",
-16252 => x"C0C0BFF982A492A4",
-16251 => x"C0C0BFF982A492F9",
-16250 => x"C0C0BFF982A492C0",
-16249 => x"C0C0BFF982A49990",
-16248 => x"C0C0BFF982A49980",
-16247 => x"C0C0BFF982A499F8",
-16246 => x"C0C0BFF982A49982",
-16245 => x"C0C0BFF982A49992",
-16244 => x"C0C0BFF982A49999",
-16243 => x"C0C0BFF982A499B0",
-16242 => x"C0C0BFF982A499A4",
-16241 => x"C0C0BFF982A499F9",
-16240 => x"C0C0BFF982A499C0",
-16239 => x"C0C0BFF982A4B090",
-16238 => x"C0C0BFF982A4B080",
-16237 => x"C0C0BFF982A4B0F8",
-16236 => x"C0C0BFF982A4B082",
-16235 => x"C0C0BFF982A4B092",
-16234 => x"C0C0BFF982A4B099",
-16233 => x"C0C0BFF982A4B0B0",
-16232 => x"C0C0BFF982A4B0A4",
-16231 => x"C0C0BFF982A4B0F9",
-16230 => x"C0C0BFF982A4B0C0",
-16229 => x"C0C0BFF982A4A490",
-16228 => x"C0C0BFF982A4A480",
-16227 => x"C0C0BFF982A4A4F8",
-16226 => x"C0C0BFF982A4A482",
-16225 => x"C0C0BFF982A4A492",
-16224 => x"C0C0BFF982A4A499",
-16223 => x"C0C0BFF982A4A4B0",
-16222 => x"C0C0BFF982A4A4A4",
-16221 => x"C0C0BFF982A4A4F9",
-16220 => x"C0C0BFF982A4A4C0",
-16219 => x"C0C0BFF982A4F990",
-16218 => x"C0C0BFF982A4F980",
-16217 => x"C0C0BFF982A4F9F8",
-16216 => x"C0C0BFF982A4F982",
-16215 => x"C0C0BFF982A4F992",
-16214 => x"C0C0BFF982A4F999",
-16213 => x"C0C0BFF982A4F9B0",
-16212 => x"C0C0BFF982A4F9A4",
-16211 => x"C0C0BFF982A4F9F9",
-16210 => x"C0C0BFF982A4F9C0",
-16209 => x"C0C0BFF982A4C090",
-16208 => x"C0C0BFF982A4C080",
-16207 => x"C0C0BFF982A4C0F8",
-16206 => x"C0C0BFF982A4C082",
-16205 => x"C0C0BFF982A4C092",
-16204 => x"C0C0BFF982A4C099",
-16203 => x"C0C0BFF982A4C0B0",
-16202 => x"C0C0BFF982A4C0A4",
-16201 => x"C0C0BFF982A4C0F9",
-16200 => x"C0C0BFF982A4C0C0",
-16199 => x"C0C0BFF982F99090",
-16198 => x"C0C0BFF982F99080",
-16197 => x"C0C0BFF982F990F8",
-16196 => x"C0C0BFF982F99082",
-16195 => x"C0C0BFF982F99092",
-16194 => x"C0C0BFF982F99099",
-16193 => x"C0C0BFF982F990B0",
-16192 => x"C0C0BFF982F990A4",
-16191 => x"C0C0BFF982F990F9",
-16190 => x"C0C0BFF982F990C0",
-16189 => x"C0C0BFF982F98090",
-16188 => x"C0C0BFF982F98080",
-16187 => x"C0C0BFF982F980F8",
-16186 => x"C0C0BFF982F98082",
-16185 => x"C0C0BFF982F98092",
-16184 => x"C0C0BFF982F98099",
-16183 => x"C0C0BFF982F980B0",
-16182 => x"C0C0BFF982F980A4",
-16181 => x"C0C0BFF982F980F9",
-16180 => x"C0C0BFF982F980C0",
-16179 => x"C0C0BFF982F9F890",
-16178 => x"C0C0BFF982F9F880",
-16177 => x"C0C0BFF982F9F8F8",
-16176 => x"C0C0BFF982F9F882",
-16175 => x"C0C0BFF982F9F892",
-16174 => x"C0C0BFF982F9F899",
-16173 => x"C0C0BFF982F9F8B0",
-16172 => x"C0C0BFF982F9F8A4",
-16171 => x"C0C0BFF982F9F8F9",
-16170 => x"C0C0BFF982F9F8C0",
-16169 => x"C0C0BFF982F98290",
-16168 => x"C0C0BFF982F98280",
-16167 => x"C0C0BFF982F982F8",
-16166 => x"C0C0BFF982F98282",
-16165 => x"C0C0BFF982F98292",
-16164 => x"C0C0BFF982F98299",
-16163 => x"C0C0BFF982F982B0",
-16162 => x"C0C0BFF982F982A4",
-16161 => x"C0C0BFF982F982F9",
-16160 => x"C0C0BFF982F982C0",
-16159 => x"C0C0BFF982F99290",
-16158 => x"C0C0BFF982F99280",
-16157 => x"C0C0BFF982F992F8",
-16156 => x"C0C0BFF982F99282",
-16155 => x"C0C0BFF982F99292",
-16154 => x"C0C0BFF982F99299",
-16153 => x"C0C0BFF982F992B0",
-16152 => x"C0C0BFF982F992A4",
-16151 => x"C0C0BFF982F992F9",
-16150 => x"C0C0BFF982F992C0",
-16149 => x"C0C0BFF982F99990",
-16148 => x"C0C0BFF982F99980",
-16147 => x"C0C0BFF982F999F8",
-16146 => x"C0C0BFF982F99982",
-16145 => x"C0C0BFF982F99992",
-16144 => x"C0C0BFF982F99999",
-16143 => x"C0C0BFF982F999B0",
-16142 => x"C0C0BFF982F999A4",
-16141 => x"C0C0BFF982F999F9",
-16140 => x"C0C0BFF982F999C0",
-16139 => x"C0C0BFF982F9B090",
-16138 => x"C0C0BFF982F9B080",
-16137 => x"C0C0BFF982F9B0F8",
-16136 => x"C0C0BFF982F9B082",
-16135 => x"C0C0BFF982F9B092",
-16134 => x"C0C0BFF982F9B099",
-16133 => x"C0C0BFF982F9B0B0",
-16132 => x"C0C0BFF982F9B0A4",
-16131 => x"C0C0BFF982F9B0F9",
-16130 => x"C0C0BFF982F9B0C0",
-16129 => x"C0C0BFF982F9A490",
-16128 => x"C0C0BFF982F9A480",
-16127 => x"C0C0BFF982F9A4F8",
-16126 => x"C0C0BFF982F9A482",
-16125 => x"C0C0BFF982F9A492",
-16124 => x"C0C0BFF982F9A499",
-16123 => x"C0C0BFF982F9A4B0",
-16122 => x"C0C0BFF982F9A4A4",
-16121 => x"C0C0BFF982F9A4F9",
-16120 => x"C0C0BFF982F9A4C0",
-16119 => x"C0C0BFF982F9F990",
-16118 => x"C0C0BFF982F9F980",
-16117 => x"C0C0BFF982F9F9F8",
-16116 => x"C0C0BFF982F9F982",
-16115 => x"C0C0BFF982F9F992",
-16114 => x"C0C0BFF982F9F999",
-16113 => x"C0C0BFF982F9F9B0",
-16112 => x"C0C0BFF982F9F9A4",
-16111 => x"C0C0BFF982F9F9F9",
-16110 => x"C0C0BFF982F9F9C0",
-16109 => x"C0C0BFF982F9C090",
-16108 => x"C0C0BFF982F9C080",
-16107 => x"C0C0BFF982F9C0F8",
-16106 => x"C0C0BFF982F9C082",
-16105 => x"C0C0BFF982F9C092",
-16104 => x"C0C0BFF982F9C099",
-16103 => x"C0C0BFF982F9C0B0",
-16102 => x"C0C0BFF982F9C0A4",
-16101 => x"C0C0BFF982F9C0F9",
-16100 => x"C0C0BFF982F9C0C0",
-16099 => x"C0C0BFF982C09090",
-16098 => x"C0C0BFF982C09080",
-16097 => x"C0C0BFF982C090F8",
-16096 => x"C0C0BFF982C09082",
-16095 => x"C0C0BFF982C09092",
-16094 => x"C0C0BFF982C09099",
-16093 => x"C0C0BFF982C090B0",
-16092 => x"C0C0BFF982C090A4",
-16091 => x"C0C0BFF982C090F9",
-16090 => x"C0C0BFF982C090C0",
-16089 => x"C0C0BFF982C08090",
-16088 => x"C0C0BFF982C08080",
-16087 => x"C0C0BFF982C080F8",
-16086 => x"C0C0BFF982C08082",
-16085 => x"C0C0BFF982C08092",
-16084 => x"C0C0BFF982C08099",
-16083 => x"C0C0BFF982C080B0",
-16082 => x"C0C0BFF982C080A4",
-16081 => x"C0C0BFF982C080F9",
-16080 => x"C0C0BFF982C080C0",
-16079 => x"C0C0BFF982C0F890",
-16078 => x"C0C0BFF982C0F880",
-16077 => x"C0C0BFF982C0F8F8",
-16076 => x"C0C0BFF982C0F882",
-16075 => x"C0C0BFF982C0F892",
-16074 => x"C0C0BFF982C0F899",
-16073 => x"C0C0BFF982C0F8B0",
-16072 => x"C0C0BFF982C0F8A4",
-16071 => x"C0C0BFF982C0F8F9",
-16070 => x"C0C0BFF982C0F8C0",
-16069 => x"C0C0BFF982C08290",
-16068 => x"C0C0BFF982C08280",
-16067 => x"C0C0BFF982C082F8",
-16066 => x"C0C0BFF982C08282",
-16065 => x"C0C0BFF982C08292",
-16064 => x"C0C0BFF982C08299",
-16063 => x"C0C0BFF982C082B0",
-16062 => x"C0C0BFF982C082A4",
-16061 => x"C0C0BFF982C082F9",
-16060 => x"C0C0BFF982C082C0",
-16059 => x"C0C0BFF982C09290",
-16058 => x"C0C0BFF982C09280",
-16057 => x"C0C0BFF982C092F8",
-16056 => x"C0C0BFF982C09282",
-16055 => x"C0C0BFF982C09292",
-16054 => x"C0C0BFF982C09299",
-16053 => x"C0C0BFF982C092B0",
-16052 => x"C0C0BFF982C092A4",
-16051 => x"C0C0BFF982C092F9",
-16050 => x"C0C0BFF982C092C0",
-16049 => x"C0C0BFF982C09990",
-16048 => x"C0C0BFF982C09980",
-16047 => x"C0C0BFF982C099F8",
-16046 => x"C0C0BFF982C09982",
-16045 => x"C0C0BFF982C09992",
-16044 => x"C0C0BFF982C09999",
-16043 => x"C0C0BFF982C099B0",
-16042 => x"C0C0BFF982C099A4",
-16041 => x"C0C0BFF982C099F9",
-16040 => x"C0C0BFF982C099C0",
-16039 => x"C0C0BFF982C0B090",
-16038 => x"C0C0BFF982C0B080",
-16037 => x"C0C0BFF982C0B0F8",
-16036 => x"C0C0BFF982C0B082",
-16035 => x"C0C0BFF982C0B092",
-16034 => x"C0C0BFF982C0B099",
-16033 => x"C0C0BFF982C0B0B0",
-16032 => x"C0C0BFF982C0B0A4",
-16031 => x"C0C0BFF982C0B0F9",
-16030 => x"C0C0BFF982C0B0C0",
-16029 => x"C0C0BFF982C0A490",
-16028 => x"C0C0BFF982C0A480",
-16027 => x"C0C0BFF982C0A4F8",
-16026 => x"C0C0BFF982C0A482",
-16025 => x"C0C0BFF982C0A492",
-16024 => x"C0C0BFF982C0A499",
-16023 => x"C0C0BFF982C0A4B0",
-16022 => x"C0C0BFF982C0A4A4",
-16021 => x"C0C0BFF982C0A4F9",
-16020 => x"C0C0BFF982C0A4C0",
-16019 => x"C0C0BFF982C0F990",
-16018 => x"C0C0BFF982C0F980",
-16017 => x"C0C0BFF982C0F9F8",
-16016 => x"C0C0BFF982C0F982",
-16015 => x"C0C0BFF982C0F992",
-16014 => x"C0C0BFF982C0F999",
-16013 => x"C0C0BFF982C0F9B0",
-16012 => x"C0C0BFF982C0F9A4",
-16011 => x"C0C0BFF982C0F9F9",
-16010 => x"C0C0BFF982C0F9C0",
-16009 => x"C0C0BFF982C0C090",
-16008 => x"C0C0BFF982C0C080",
-16007 => x"C0C0BFF982C0C0F8",
-16006 => x"C0C0BFF982C0C082",
-16005 => x"C0C0BFF982C0C092",
-16004 => x"C0C0BFF982C0C099",
-16003 => x"C0C0BFF982C0C0B0",
-16002 => x"C0C0BFF982C0C0A4",
-16001 => x"C0C0BFF982C0C0F9",
-16000 => x"C0C0BFF982C0C0C0",
-15999 => x"C0C0BFF992909090",
-15998 => x"C0C0BFF992909080",
-15997 => x"C0C0BFF9929090F8",
-15996 => x"C0C0BFF992909082",
-15995 => x"C0C0BFF992909092",
-15994 => x"C0C0BFF992909099",
-15993 => x"C0C0BFF9929090B0",
-15992 => x"C0C0BFF9929090A4",
-15991 => x"C0C0BFF9929090F9",
-15990 => x"C0C0BFF9929090C0",
-15989 => x"C0C0BFF992908090",
-15988 => x"C0C0BFF992908080",
-15987 => x"C0C0BFF9929080F8",
-15986 => x"C0C0BFF992908082",
-15985 => x"C0C0BFF992908092",
-15984 => x"C0C0BFF992908099",
-15983 => x"C0C0BFF9929080B0",
-15982 => x"C0C0BFF9929080A4",
-15981 => x"C0C0BFF9929080F9",
-15980 => x"C0C0BFF9929080C0",
-15979 => x"C0C0BFF99290F890",
-15978 => x"C0C0BFF99290F880",
-15977 => x"C0C0BFF99290F8F8",
-15976 => x"C0C0BFF99290F882",
-15975 => x"C0C0BFF99290F892",
-15974 => x"C0C0BFF99290F899",
-15973 => x"C0C0BFF99290F8B0",
-15972 => x"C0C0BFF99290F8A4",
-15971 => x"C0C0BFF99290F8F9",
-15970 => x"C0C0BFF99290F8C0",
-15969 => x"C0C0BFF992908290",
-15968 => x"C0C0BFF992908280",
-15967 => x"C0C0BFF9929082F8",
-15966 => x"C0C0BFF992908282",
-15965 => x"C0C0BFF992908292",
-15964 => x"C0C0BFF992908299",
-15963 => x"C0C0BFF9929082B0",
-15962 => x"C0C0BFF9929082A4",
-15961 => x"C0C0BFF9929082F9",
-15960 => x"C0C0BFF9929082C0",
-15959 => x"C0C0BFF992909290",
-15958 => x"C0C0BFF992909280",
-15957 => x"C0C0BFF9929092F8",
-15956 => x"C0C0BFF992909282",
-15955 => x"C0C0BFF992909292",
-15954 => x"C0C0BFF992909299",
-15953 => x"C0C0BFF9929092B0",
-15952 => x"C0C0BFF9929092A4",
-15951 => x"C0C0BFF9929092F9",
-15950 => x"C0C0BFF9929092C0",
-15949 => x"C0C0BFF992909990",
-15948 => x"C0C0BFF992909980",
-15947 => x"C0C0BFF9929099F8",
-15946 => x"C0C0BFF992909982",
-15945 => x"C0C0BFF992909992",
-15944 => x"C0C0BFF992909999",
-15943 => x"C0C0BFF9929099B0",
-15942 => x"C0C0BFF9929099A4",
-15941 => x"C0C0BFF9929099F9",
-15940 => x"C0C0BFF9929099C0",
-15939 => x"C0C0BFF99290B090",
-15938 => x"C0C0BFF99290B080",
-15937 => x"C0C0BFF99290B0F8",
-15936 => x"C0C0BFF99290B082",
-15935 => x"C0C0BFF99290B092",
-15934 => x"C0C0BFF99290B099",
-15933 => x"C0C0BFF99290B0B0",
-15932 => x"C0C0BFF99290B0A4",
-15931 => x"C0C0BFF99290B0F9",
-15930 => x"C0C0BFF99290B0C0",
-15929 => x"C0C0BFF99290A490",
-15928 => x"C0C0BFF99290A480",
-15927 => x"C0C0BFF99290A4F8",
-15926 => x"C0C0BFF99290A482",
-15925 => x"C0C0BFF99290A492",
-15924 => x"C0C0BFF99290A499",
-15923 => x"C0C0BFF99290A4B0",
-15922 => x"C0C0BFF99290A4A4",
-15921 => x"C0C0BFF99290A4F9",
-15920 => x"C0C0BFF99290A4C0",
-15919 => x"C0C0BFF99290F990",
-15918 => x"C0C0BFF99290F980",
-15917 => x"C0C0BFF99290F9F8",
-15916 => x"C0C0BFF99290F982",
-15915 => x"C0C0BFF99290F992",
-15914 => x"C0C0BFF99290F999",
-15913 => x"C0C0BFF99290F9B0",
-15912 => x"C0C0BFF99290F9A4",
-15911 => x"C0C0BFF99290F9F9",
-15910 => x"C0C0BFF99290F9C0",
-15909 => x"C0C0BFF99290C090",
-15908 => x"C0C0BFF99290C080",
-15907 => x"C0C0BFF99290C0F8",
-15906 => x"C0C0BFF99290C082",
-15905 => x"C0C0BFF99290C092",
-15904 => x"C0C0BFF99290C099",
-15903 => x"C0C0BFF99290C0B0",
-15902 => x"C0C0BFF99290C0A4",
-15901 => x"C0C0BFF99290C0F9",
-15900 => x"C0C0BFF99290C0C0",
-15899 => x"C0C0BFF992809090",
-15898 => x"C0C0BFF992809080",
-15897 => x"C0C0BFF9928090F8",
-15896 => x"C0C0BFF992809082",
-15895 => x"C0C0BFF992809092",
-15894 => x"C0C0BFF992809099",
-15893 => x"C0C0BFF9928090B0",
-15892 => x"C0C0BFF9928090A4",
-15891 => x"C0C0BFF9928090F9",
-15890 => x"C0C0BFF9928090C0",
-15889 => x"C0C0BFF992808090",
-15888 => x"C0C0BFF992808080",
-15887 => x"C0C0BFF9928080F8",
-15886 => x"C0C0BFF992808082",
-15885 => x"C0C0BFF992808092",
-15884 => x"C0C0BFF992808099",
-15883 => x"C0C0BFF9928080B0",
-15882 => x"C0C0BFF9928080A4",
-15881 => x"C0C0BFF9928080F9",
-15880 => x"C0C0BFF9928080C0",
-15879 => x"C0C0BFF99280F890",
-15878 => x"C0C0BFF99280F880",
-15877 => x"C0C0BFF99280F8F8",
-15876 => x"C0C0BFF99280F882",
-15875 => x"C0C0BFF99280F892",
-15874 => x"C0C0BFF99280F899",
-15873 => x"C0C0BFF99280F8B0",
-15872 => x"C0C0BFF99280F8A4",
-15871 => x"C0C0BFF99280F8F9",
-15870 => x"C0C0BFF99280F8C0",
-15869 => x"C0C0BFF992808290",
-15868 => x"C0C0BFF992808280",
-15867 => x"C0C0BFF9928082F8",
-15866 => x"C0C0BFF992808282",
-15865 => x"C0C0BFF992808292",
-15864 => x"C0C0BFF992808299",
-15863 => x"C0C0BFF9928082B0",
-15862 => x"C0C0BFF9928082A4",
-15861 => x"C0C0BFF9928082F9",
-15860 => x"C0C0BFF9928082C0",
-15859 => x"C0C0BFF992809290",
-15858 => x"C0C0BFF992809280",
-15857 => x"C0C0BFF9928092F8",
-15856 => x"C0C0BFF992809282",
-15855 => x"C0C0BFF992809292",
-15854 => x"C0C0BFF992809299",
-15853 => x"C0C0BFF9928092B0",
-15852 => x"C0C0BFF9928092A4",
-15851 => x"C0C0BFF9928092F9",
-15850 => x"C0C0BFF9928092C0",
-15849 => x"C0C0BFF992809990",
-15848 => x"C0C0BFF992809980",
-15847 => x"C0C0BFF9928099F8",
-15846 => x"C0C0BFF992809982",
-15845 => x"C0C0BFF992809992",
-15844 => x"C0C0BFF992809999",
-15843 => x"C0C0BFF9928099B0",
-15842 => x"C0C0BFF9928099A4",
-15841 => x"C0C0BFF9928099F9",
-15840 => x"C0C0BFF9928099C0",
-15839 => x"C0C0BFF99280B090",
-15838 => x"C0C0BFF99280B080",
-15837 => x"C0C0BFF99280B0F8",
-15836 => x"C0C0BFF99280B082",
-15835 => x"C0C0BFF99280B092",
-15834 => x"C0C0BFF99280B099",
-15833 => x"C0C0BFF99280B0B0",
-15832 => x"C0C0BFF99280B0A4",
-15831 => x"C0C0BFF99280B0F9",
-15830 => x"C0C0BFF99280B0C0",
-15829 => x"C0C0BFF99280A490",
-15828 => x"C0C0BFF99280A480",
-15827 => x"C0C0BFF99280A4F8",
-15826 => x"C0C0BFF99280A482",
-15825 => x"C0C0BFF99280A492",
-15824 => x"C0C0BFF99280A499",
-15823 => x"C0C0BFF99280A4B0",
-15822 => x"C0C0BFF99280A4A4",
-15821 => x"C0C0BFF99280A4F9",
-15820 => x"C0C0BFF99280A4C0",
-15819 => x"C0C0BFF99280F990",
-15818 => x"C0C0BFF99280F980",
-15817 => x"C0C0BFF99280F9F8",
-15816 => x"C0C0BFF99280F982",
-15815 => x"C0C0BFF99280F992",
-15814 => x"C0C0BFF99280F999",
-15813 => x"C0C0BFF99280F9B0",
-15812 => x"C0C0BFF99280F9A4",
-15811 => x"C0C0BFF99280F9F9",
-15810 => x"C0C0BFF99280F9C0",
-15809 => x"C0C0BFF99280C090",
-15808 => x"C0C0BFF99280C080",
-15807 => x"C0C0BFF99280C0F8",
-15806 => x"C0C0BFF99280C082",
-15805 => x"C0C0BFF99280C092",
-15804 => x"C0C0BFF99280C099",
-15803 => x"C0C0BFF99280C0B0",
-15802 => x"C0C0BFF99280C0A4",
-15801 => x"C0C0BFF99280C0F9",
-15800 => x"C0C0BFF99280C0C0",
-15799 => x"C0C0BFF992F89090",
-15798 => x"C0C0BFF992F89080",
-15797 => x"C0C0BFF992F890F8",
-15796 => x"C0C0BFF992F89082",
-15795 => x"C0C0BFF992F89092",
-15794 => x"C0C0BFF992F89099",
-15793 => x"C0C0BFF992F890B0",
-15792 => x"C0C0BFF992F890A4",
-15791 => x"C0C0BFF992F890F9",
-15790 => x"C0C0BFF992F890C0",
-15789 => x"C0C0BFF992F88090",
-15788 => x"C0C0BFF992F88080",
-15787 => x"C0C0BFF992F880F8",
-15786 => x"C0C0BFF992F88082",
-15785 => x"C0C0BFF992F88092",
-15784 => x"C0C0BFF992F88099",
-15783 => x"C0C0BFF992F880B0",
-15782 => x"C0C0BFF992F880A4",
-15781 => x"C0C0BFF992F880F9",
-15780 => x"C0C0BFF992F880C0",
-15779 => x"C0C0BFF992F8F890",
-15778 => x"C0C0BFF992F8F880",
-15777 => x"C0C0BFF992F8F8F8",
-15776 => x"C0C0BFF992F8F882",
-15775 => x"C0C0BFF992F8F892",
-15774 => x"C0C0BFF992F8F899",
-15773 => x"C0C0BFF992F8F8B0",
-15772 => x"C0C0BFF992F8F8A4",
-15771 => x"C0C0BFF992F8F8F9",
-15770 => x"C0C0BFF992F8F8C0",
-15769 => x"C0C0BFF992F88290",
-15768 => x"C0C0BFF992F88280",
-15767 => x"C0C0BFF992F882F8",
-15766 => x"C0C0BFF992F88282",
-15765 => x"C0C0BFF992F88292",
-15764 => x"C0C0BFF992F88299",
-15763 => x"C0C0BFF992F882B0",
-15762 => x"C0C0BFF992F882A4",
-15761 => x"C0C0BFF992F882F9",
-15760 => x"C0C0BFF992F882C0",
-15759 => x"C0C0BFF992F89290",
-15758 => x"C0C0BFF992F89280",
-15757 => x"C0C0BFF992F892F8",
-15756 => x"C0C0BFF992F89282",
-15755 => x"C0C0BFF992F89292",
-15754 => x"C0C0BFF992F89299",
-15753 => x"C0C0BFF992F892B0",
-15752 => x"C0C0BFF992F892A4",
-15751 => x"C0C0BFF992F892F9",
-15750 => x"C0C0BFF992F892C0",
-15749 => x"C0C0BFF992F89990",
-15748 => x"C0C0BFF992F89980",
-15747 => x"C0C0BFF992F899F8",
-15746 => x"C0C0BFF992F89982",
-15745 => x"C0C0BFF992F89992",
-15744 => x"C0C0BFF992F89999",
-15743 => x"C0C0BFF992F899B0",
-15742 => x"C0C0BFF992F899A4",
-15741 => x"C0C0BFF992F899F9",
-15740 => x"C0C0BFF992F899C0",
-15739 => x"C0C0BFF992F8B090",
-15738 => x"C0C0BFF992F8B080",
-15737 => x"C0C0BFF992F8B0F8",
-15736 => x"C0C0BFF992F8B082",
-15735 => x"C0C0BFF992F8B092",
-15734 => x"C0C0BFF992F8B099",
-15733 => x"C0C0BFF992F8B0B0",
-15732 => x"C0C0BFF992F8B0A4",
-15731 => x"C0C0BFF992F8B0F9",
-15730 => x"C0C0BFF992F8B0C0",
-15729 => x"C0C0BFF992F8A490",
-15728 => x"C0C0BFF992F8A480",
-15727 => x"C0C0BFF992F8A4F8",
-15726 => x"C0C0BFF992F8A482",
-15725 => x"C0C0BFF992F8A492",
-15724 => x"C0C0BFF992F8A499",
-15723 => x"C0C0BFF992F8A4B0",
-15722 => x"C0C0BFF992F8A4A4",
-15721 => x"C0C0BFF992F8A4F9",
-15720 => x"C0C0BFF992F8A4C0",
-15719 => x"C0C0BFF992F8F990",
-15718 => x"C0C0BFF992F8F980",
-15717 => x"C0C0BFF992F8F9F8",
-15716 => x"C0C0BFF992F8F982",
-15715 => x"C0C0BFF992F8F992",
-15714 => x"C0C0BFF992F8F999",
-15713 => x"C0C0BFF992F8F9B0",
-15712 => x"C0C0BFF992F8F9A4",
-15711 => x"C0C0BFF992F8F9F9",
-15710 => x"C0C0BFF992F8F9C0",
-15709 => x"C0C0BFF992F8C090",
-15708 => x"C0C0BFF992F8C080",
-15707 => x"C0C0BFF992F8C0F8",
-15706 => x"C0C0BFF992F8C082",
-15705 => x"C0C0BFF992F8C092",
-15704 => x"C0C0BFF992F8C099",
-15703 => x"C0C0BFF992F8C0B0",
-15702 => x"C0C0BFF992F8C0A4",
-15701 => x"C0C0BFF992F8C0F9",
-15700 => x"C0C0BFF992F8C0C0",
-15699 => x"C0C0BFF992829090",
-15698 => x"C0C0BFF992829080",
-15697 => x"C0C0BFF9928290F8",
-15696 => x"C0C0BFF992829082",
-15695 => x"C0C0BFF992829092",
-15694 => x"C0C0BFF992829099",
-15693 => x"C0C0BFF9928290B0",
-15692 => x"C0C0BFF9928290A4",
-15691 => x"C0C0BFF9928290F9",
-15690 => x"C0C0BFF9928290C0",
-15689 => x"C0C0BFF992828090",
-15688 => x"C0C0BFF992828080",
-15687 => x"C0C0BFF9928280F8",
-15686 => x"C0C0BFF992828082",
-15685 => x"C0C0BFF992828092",
-15684 => x"C0C0BFF992828099",
-15683 => x"C0C0BFF9928280B0",
-15682 => x"C0C0BFF9928280A4",
-15681 => x"C0C0BFF9928280F9",
-15680 => x"C0C0BFF9928280C0",
-15679 => x"C0C0BFF99282F890",
-15678 => x"C0C0BFF99282F880",
-15677 => x"C0C0BFF99282F8F8",
-15676 => x"C0C0BFF99282F882",
-15675 => x"C0C0BFF99282F892",
-15674 => x"C0C0BFF99282F899",
-15673 => x"C0C0BFF99282F8B0",
-15672 => x"C0C0BFF99282F8A4",
-15671 => x"C0C0BFF99282F8F9",
-15670 => x"C0C0BFF99282F8C0",
-15669 => x"C0C0BFF992828290",
-15668 => x"C0C0BFF992828280",
-15667 => x"C0C0BFF9928282F8",
-15666 => x"C0C0BFF992828282",
-15665 => x"C0C0BFF992828292",
-15664 => x"C0C0BFF992828299",
-15663 => x"C0C0BFF9928282B0",
-15662 => x"C0C0BFF9928282A4",
-15661 => x"C0C0BFF9928282F9",
-15660 => x"C0C0BFF9928282C0",
-15659 => x"C0C0BFF992829290",
-15658 => x"C0C0BFF992829280",
-15657 => x"C0C0BFF9928292F8",
-15656 => x"C0C0BFF992829282",
-15655 => x"C0C0BFF992829292",
-15654 => x"C0C0BFF992829299",
-15653 => x"C0C0BFF9928292B0",
-15652 => x"C0C0BFF9928292A4",
-15651 => x"C0C0BFF9928292F9",
-15650 => x"C0C0BFF9928292C0",
-15649 => x"C0C0BFF992829990",
-15648 => x"C0C0BFF992829980",
-15647 => x"C0C0BFF9928299F8",
-15646 => x"C0C0BFF992829982",
-15645 => x"C0C0BFF992829992",
-15644 => x"C0C0BFF992829999",
-15643 => x"C0C0BFF9928299B0",
-15642 => x"C0C0BFF9928299A4",
-15641 => x"C0C0BFF9928299F9",
-15640 => x"C0C0BFF9928299C0",
-15639 => x"C0C0BFF99282B090",
-15638 => x"C0C0BFF99282B080",
-15637 => x"C0C0BFF99282B0F8",
-15636 => x"C0C0BFF99282B082",
-15635 => x"C0C0BFF99282B092",
-15634 => x"C0C0BFF99282B099",
-15633 => x"C0C0BFF99282B0B0",
-15632 => x"C0C0BFF99282B0A4",
-15631 => x"C0C0BFF99282B0F9",
-15630 => x"C0C0BFF99282B0C0",
-15629 => x"C0C0BFF99282A490",
-15628 => x"C0C0BFF99282A480",
-15627 => x"C0C0BFF99282A4F8",
-15626 => x"C0C0BFF99282A482",
-15625 => x"C0C0BFF99282A492",
-15624 => x"C0C0BFF99282A499",
-15623 => x"C0C0BFF99282A4B0",
-15622 => x"C0C0BFF99282A4A4",
-15621 => x"C0C0BFF99282A4F9",
-15620 => x"C0C0BFF99282A4C0",
-15619 => x"C0C0BFF99282F990",
-15618 => x"C0C0BFF99282F980",
-15617 => x"C0C0BFF99282F9F8",
-15616 => x"C0C0BFF99282F982",
-15615 => x"C0C0BFF99282F992",
-15614 => x"C0C0BFF99282F999",
-15613 => x"C0C0BFF99282F9B0",
-15612 => x"C0C0BFF99282F9A4",
-15611 => x"C0C0BFF99282F9F9",
-15610 => x"C0C0BFF99282F9C0",
-15609 => x"C0C0BFF99282C090",
-15608 => x"C0C0BFF99282C080",
-15607 => x"C0C0BFF99282C0F8",
-15606 => x"C0C0BFF99282C082",
-15605 => x"C0C0BFF99282C092",
-15604 => x"C0C0BFF99282C099",
-15603 => x"C0C0BFF99282C0B0",
-15602 => x"C0C0BFF99282C0A4",
-15601 => x"C0C0BFF99282C0F9",
-15600 => x"C0C0BFF99282C0C0",
-15599 => x"C0C0BFF992929090",
-15598 => x"C0C0BFF992929080",
-15597 => x"C0C0BFF9929290F8",
-15596 => x"C0C0BFF992929082",
-15595 => x"C0C0BFF992929092",
-15594 => x"C0C0BFF992929099",
-15593 => x"C0C0BFF9929290B0",
-15592 => x"C0C0BFF9929290A4",
-15591 => x"C0C0BFF9929290F9",
-15590 => x"C0C0BFF9929290C0",
-15589 => x"C0C0BFF992928090",
-15588 => x"C0C0BFF992928080",
-15587 => x"C0C0BFF9929280F8",
-15586 => x"C0C0BFF992928082",
-15585 => x"C0C0BFF992928092",
-15584 => x"C0C0BFF992928099",
-15583 => x"C0C0BFF9929280B0",
-15582 => x"C0C0BFF9929280A4",
-15581 => x"C0C0BFF9929280F9",
-15580 => x"C0C0BFF9929280C0",
-15579 => x"C0C0BFF99292F890",
-15578 => x"C0C0BFF99292F880",
-15577 => x"C0C0BFF99292F8F8",
-15576 => x"C0C0BFF99292F882",
-15575 => x"C0C0BFF99292F892",
-15574 => x"C0C0BFF99292F899",
-15573 => x"C0C0BFF99292F8B0",
-15572 => x"C0C0BFF99292F8A4",
-15571 => x"C0C0BFF99292F8F9",
-15570 => x"C0C0BFF99292F8C0",
-15569 => x"C0C0BFF992928290",
-15568 => x"C0C0BFF992928280",
-15567 => x"C0C0BFF9929282F8",
-15566 => x"C0C0BFF992928282",
-15565 => x"C0C0BFF992928292",
-15564 => x"C0C0BFF992928299",
-15563 => x"C0C0BFF9929282B0",
-15562 => x"C0C0BFF9929282A4",
-15561 => x"C0C0BFF9929282F9",
-15560 => x"C0C0BFF9929282C0",
-15559 => x"C0C0BFF992929290",
-15558 => x"C0C0BFF992929280",
-15557 => x"C0C0BFF9929292F8",
-15556 => x"C0C0BFF992929282",
-15555 => x"C0C0BFF992929292",
-15554 => x"C0C0BFF992929299",
-15553 => x"C0C0BFF9929292B0",
-15552 => x"C0C0BFF9929292A4",
-15551 => x"C0C0BFF9929292F9",
-15550 => x"C0C0BFF9929292C0",
-15549 => x"C0C0BFF992929990",
-15548 => x"C0C0BFF992929980",
-15547 => x"C0C0BFF9929299F8",
-15546 => x"C0C0BFF992929982",
-15545 => x"C0C0BFF992929992",
-15544 => x"C0C0BFF992929999",
-15543 => x"C0C0BFF9929299B0",
-15542 => x"C0C0BFF9929299A4",
-15541 => x"C0C0BFF9929299F9",
-15540 => x"C0C0BFF9929299C0",
-15539 => x"C0C0BFF99292B090",
-15538 => x"C0C0BFF99292B080",
-15537 => x"C0C0BFF99292B0F8",
-15536 => x"C0C0BFF99292B082",
-15535 => x"C0C0BFF99292B092",
-15534 => x"C0C0BFF99292B099",
-15533 => x"C0C0BFF99292B0B0",
-15532 => x"C0C0BFF99292B0A4",
-15531 => x"C0C0BFF99292B0F9",
-15530 => x"C0C0BFF99292B0C0",
-15529 => x"C0C0BFF99292A490",
-15528 => x"C0C0BFF99292A480",
-15527 => x"C0C0BFF99292A4F8",
-15526 => x"C0C0BFF99292A482",
-15525 => x"C0C0BFF99292A492",
-15524 => x"C0C0BFF99292A499",
-15523 => x"C0C0BFF99292A4B0",
-15522 => x"C0C0BFF99292A4A4",
-15521 => x"C0C0BFF99292A4F9",
-15520 => x"C0C0BFF99292A4C0",
-15519 => x"C0C0BFF99292F990",
-15518 => x"C0C0BFF99292F980",
-15517 => x"C0C0BFF99292F9F8",
-15516 => x"C0C0BFF99292F982",
-15515 => x"C0C0BFF99292F992",
-15514 => x"C0C0BFF99292F999",
-15513 => x"C0C0BFF99292F9B0",
-15512 => x"C0C0BFF99292F9A4",
-15511 => x"C0C0BFF99292F9F9",
-15510 => x"C0C0BFF99292F9C0",
-15509 => x"C0C0BFF99292C090",
-15508 => x"C0C0BFF99292C080",
-15507 => x"C0C0BFF99292C0F8",
-15506 => x"C0C0BFF99292C082",
-15505 => x"C0C0BFF99292C092",
-15504 => x"C0C0BFF99292C099",
-15503 => x"C0C0BFF99292C0B0",
-15502 => x"C0C0BFF99292C0A4",
-15501 => x"C0C0BFF99292C0F9",
-15500 => x"C0C0BFF99292C0C0",
-15499 => x"C0C0BFF992999090",
-15498 => x"C0C0BFF992999080",
-15497 => x"C0C0BFF9929990F8",
-15496 => x"C0C0BFF992999082",
-15495 => x"C0C0BFF992999092",
-15494 => x"C0C0BFF992999099",
-15493 => x"C0C0BFF9929990B0",
-15492 => x"C0C0BFF9929990A4",
-15491 => x"C0C0BFF9929990F9",
-15490 => x"C0C0BFF9929990C0",
-15489 => x"C0C0BFF992998090",
-15488 => x"C0C0BFF992998080",
-15487 => x"C0C0BFF9929980F8",
-15486 => x"C0C0BFF992998082",
-15485 => x"C0C0BFF992998092",
-15484 => x"C0C0BFF992998099",
-15483 => x"C0C0BFF9929980B0",
-15482 => x"C0C0BFF9929980A4",
-15481 => x"C0C0BFF9929980F9",
-15480 => x"C0C0BFF9929980C0",
-15479 => x"C0C0BFF99299F890",
-15478 => x"C0C0BFF99299F880",
-15477 => x"C0C0BFF99299F8F8",
-15476 => x"C0C0BFF99299F882",
-15475 => x"C0C0BFF99299F892",
-15474 => x"C0C0BFF99299F899",
-15473 => x"C0C0BFF99299F8B0",
-15472 => x"C0C0BFF99299F8A4",
-15471 => x"C0C0BFF99299F8F9",
-15470 => x"C0C0BFF99299F8C0",
-15469 => x"C0C0BFF992998290",
-15468 => x"C0C0BFF992998280",
-15467 => x"C0C0BFF9929982F8",
-15466 => x"C0C0BFF992998282",
-15465 => x"C0C0BFF992998292",
-15464 => x"C0C0BFF992998299",
-15463 => x"C0C0BFF9929982B0",
-15462 => x"C0C0BFF9929982A4",
-15461 => x"C0C0BFF9929982F9",
-15460 => x"C0C0BFF9929982C0",
-15459 => x"C0C0BFF992999290",
-15458 => x"C0C0BFF992999280",
-15457 => x"C0C0BFF9929992F8",
-15456 => x"C0C0BFF992999282",
-15455 => x"C0C0BFF992999292",
-15454 => x"C0C0BFF992999299",
-15453 => x"C0C0BFF9929992B0",
-15452 => x"C0C0BFF9929992A4",
-15451 => x"C0C0BFF9929992F9",
-15450 => x"C0C0BFF9929992C0",
-15449 => x"C0C0BFF992999990",
-15448 => x"C0C0BFF992999980",
-15447 => x"C0C0BFF9929999F8",
-15446 => x"C0C0BFF992999982",
-15445 => x"C0C0BFF992999992",
-15444 => x"C0C0BFF992999999",
-15443 => x"C0C0BFF9929999B0",
-15442 => x"C0C0BFF9929999A4",
-15441 => x"C0C0BFF9929999F9",
-15440 => x"C0C0BFF9929999C0",
-15439 => x"C0C0BFF99299B090",
-15438 => x"C0C0BFF99299B080",
-15437 => x"C0C0BFF99299B0F8",
-15436 => x"C0C0BFF99299B082",
-15435 => x"C0C0BFF99299B092",
-15434 => x"C0C0BFF99299B099",
-15433 => x"C0C0BFF99299B0B0",
-15432 => x"C0C0BFF99299B0A4",
-15431 => x"C0C0BFF99299B0F9",
-15430 => x"C0C0BFF99299B0C0",
-15429 => x"C0C0BFF99299A490",
-15428 => x"C0C0BFF99299A480",
-15427 => x"C0C0BFF99299A4F8",
-15426 => x"C0C0BFF99299A482",
-15425 => x"C0C0BFF99299A492",
-15424 => x"C0C0BFF99299A499",
-15423 => x"C0C0BFF99299A4B0",
-15422 => x"C0C0BFF99299A4A4",
-15421 => x"C0C0BFF99299A4F9",
-15420 => x"C0C0BFF99299A4C0",
-15419 => x"C0C0BFF99299F990",
-15418 => x"C0C0BFF99299F980",
-15417 => x"C0C0BFF99299F9F8",
-15416 => x"C0C0BFF99299F982",
-15415 => x"C0C0BFF99299F992",
-15414 => x"C0C0BFF99299F999",
-15413 => x"C0C0BFF99299F9B0",
-15412 => x"C0C0BFF99299F9A4",
-15411 => x"C0C0BFF99299F9F9",
-15410 => x"C0C0BFF99299F9C0",
-15409 => x"C0C0BFF99299C090",
-15408 => x"C0C0BFF99299C080",
-15407 => x"C0C0BFF99299C0F8",
-15406 => x"C0C0BFF99299C082",
-15405 => x"C0C0BFF99299C092",
-15404 => x"C0C0BFF99299C099",
-15403 => x"C0C0BFF99299C0B0",
-15402 => x"C0C0BFF99299C0A4",
-15401 => x"C0C0BFF99299C0F9",
-15400 => x"C0C0BFF99299C0C0",
-15399 => x"C0C0BFF992B09090",
-15398 => x"C0C0BFF992B09080",
-15397 => x"C0C0BFF992B090F8",
-15396 => x"C0C0BFF992B09082",
-15395 => x"C0C0BFF992B09092",
-15394 => x"C0C0BFF992B09099",
-15393 => x"C0C0BFF992B090B0",
-15392 => x"C0C0BFF992B090A4",
-15391 => x"C0C0BFF992B090F9",
-15390 => x"C0C0BFF992B090C0",
-15389 => x"C0C0BFF992B08090",
-15388 => x"C0C0BFF992B08080",
-15387 => x"C0C0BFF992B080F8",
-15386 => x"C0C0BFF992B08082",
-15385 => x"C0C0BFF992B08092",
-15384 => x"C0C0BFF992B08099",
-15383 => x"C0C0BFF992B080B0",
-15382 => x"C0C0BFF992B080A4",
-15381 => x"C0C0BFF992B080F9",
-15380 => x"C0C0BFF992B080C0",
-15379 => x"C0C0BFF992B0F890",
-15378 => x"C0C0BFF992B0F880",
-15377 => x"C0C0BFF992B0F8F8",
-15376 => x"C0C0BFF992B0F882",
-15375 => x"C0C0BFF992B0F892",
-15374 => x"C0C0BFF992B0F899",
-15373 => x"C0C0BFF992B0F8B0",
-15372 => x"C0C0BFF992B0F8A4",
-15371 => x"C0C0BFF992B0F8F9",
-15370 => x"C0C0BFF992B0F8C0",
-15369 => x"C0C0BFF992B08290",
-15368 => x"C0C0BFF992B08280",
-15367 => x"C0C0BFF992B082F8",
-15366 => x"C0C0BFF992B08282",
-15365 => x"C0C0BFF992B08292",
-15364 => x"C0C0BFF992B08299",
-15363 => x"C0C0BFF992B082B0",
-15362 => x"C0C0BFF992B082A4",
-15361 => x"C0C0BFF992B082F9",
-15360 => x"C0C0BFF992B082C0",
-15359 => x"C0C0BFF992B09290",
-15358 => x"C0C0BFF992B09280",
-15357 => x"C0C0BFF992B092F8",
-15356 => x"C0C0BFF992B09282",
-15355 => x"C0C0BFF992B09292",
-15354 => x"C0C0BFF992B09299",
-15353 => x"C0C0BFF992B092B0",
-15352 => x"C0C0BFF992B092A4",
-15351 => x"C0C0BFF992B092F9",
-15350 => x"C0C0BFF992B092C0",
-15349 => x"C0C0BFF992B09990",
-15348 => x"C0C0BFF992B09980",
-15347 => x"C0C0BFF992B099F8",
-15346 => x"C0C0BFF992B09982",
-15345 => x"C0C0BFF992B09992",
-15344 => x"C0C0BFF992B09999",
-15343 => x"C0C0BFF992B099B0",
-15342 => x"C0C0BFF992B099A4",
-15341 => x"C0C0BFF992B099F9",
-15340 => x"C0C0BFF992B099C0",
-15339 => x"C0C0BFF992B0B090",
-15338 => x"C0C0BFF992B0B080",
-15337 => x"C0C0BFF992B0B0F8",
-15336 => x"C0C0BFF992B0B082",
-15335 => x"C0C0BFF992B0B092",
-15334 => x"C0C0BFF992B0B099",
-15333 => x"C0C0BFF992B0B0B0",
-15332 => x"C0C0BFF992B0B0A4",
-15331 => x"C0C0BFF992B0B0F9",
-15330 => x"C0C0BFF992B0B0C0",
-15329 => x"C0C0BFF992B0A490",
-15328 => x"C0C0BFF992B0A480",
-15327 => x"C0C0BFF992B0A4F8",
-15326 => x"C0C0BFF992B0A482",
-15325 => x"C0C0BFF992B0A492",
-15324 => x"C0C0BFF992B0A499",
-15323 => x"C0C0BFF992B0A4B0",
-15322 => x"C0C0BFF992B0A4A4",
-15321 => x"C0C0BFF992B0A4F9",
-15320 => x"C0C0BFF992B0A4C0",
-15319 => x"C0C0BFF992B0F990",
-15318 => x"C0C0BFF992B0F980",
-15317 => x"C0C0BFF992B0F9F8",
-15316 => x"C0C0BFF992B0F982",
-15315 => x"C0C0BFF992B0F992",
-15314 => x"C0C0BFF992B0F999",
-15313 => x"C0C0BFF992B0F9B0",
-15312 => x"C0C0BFF992B0F9A4",
-15311 => x"C0C0BFF992B0F9F9",
-15310 => x"C0C0BFF992B0F9C0",
-15309 => x"C0C0BFF992B0C090",
-15308 => x"C0C0BFF992B0C080",
-15307 => x"C0C0BFF992B0C0F8",
-15306 => x"C0C0BFF992B0C082",
-15305 => x"C0C0BFF992B0C092",
-15304 => x"C0C0BFF992B0C099",
-15303 => x"C0C0BFF992B0C0B0",
-15302 => x"C0C0BFF992B0C0A4",
-15301 => x"C0C0BFF992B0C0F9",
-15300 => x"C0C0BFF992B0C0C0",
-15299 => x"C0C0BFF992A49090",
-15298 => x"C0C0BFF992A49080",
-15297 => x"C0C0BFF992A490F8",
-15296 => x"C0C0BFF992A49082",
-15295 => x"C0C0BFF992A49092",
-15294 => x"C0C0BFF992A49099",
-15293 => x"C0C0BFF992A490B0",
-15292 => x"C0C0BFF992A490A4",
-15291 => x"C0C0BFF992A490F9",
-15290 => x"C0C0BFF992A490C0",
-15289 => x"C0C0BFF992A48090",
-15288 => x"C0C0BFF992A48080",
-15287 => x"C0C0BFF992A480F8",
-15286 => x"C0C0BFF992A48082",
-15285 => x"C0C0BFF992A48092",
-15284 => x"C0C0BFF992A48099",
-15283 => x"C0C0BFF992A480B0",
-15282 => x"C0C0BFF992A480A4",
-15281 => x"C0C0BFF992A480F9",
-15280 => x"C0C0BFF992A480C0",
-15279 => x"C0C0BFF992A4F890",
-15278 => x"C0C0BFF992A4F880",
-15277 => x"C0C0BFF992A4F8F8",
-15276 => x"C0C0BFF992A4F882",
-15275 => x"C0C0BFF992A4F892",
-15274 => x"C0C0BFF992A4F899",
-15273 => x"C0C0BFF992A4F8B0",
-15272 => x"C0C0BFF992A4F8A4",
-15271 => x"C0C0BFF992A4F8F9",
-15270 => x"C0C0BFF992A4F8C0",
-15269 => x"C0C0BFF992A48290",
-15268 => x"C0C0BFF992A48280",
-15267 => x"C0C0BFF992A482F8",
-15266 => x"C0C0BFF992A48282",
-15265 => x"C0C0BFF992A48292",
-15264 => x"C0C0BFF992A48299",
-15263 => x"C0C0BFF992A482B0",
-15262 => x"C0C0BFF992A482A4",
-15261 => x"C0C0BFF992A482F9",
-15260 => x"C0C0BFF992A482C0",
-15259 => x"C0C0BFF992A49290",
-15258 => x"C0C0BFF992A49280",
-15257 => x"C0C0BFF992A492F8",
-15256 => x"C0C0BFF992A49282",
-15255 => x"C0C0BFF992A49292",
-15254 => x"C0C0BFF992A49299",
-15253 => x"C0C0BFF992A492B0",
-15252 => x"C0C0BFF992A492A4",
-15251 => x"C0C0BFF992A492F9",
-15250 => x"C0C0BFF992A492C0",
-15249 => x"C0C0BFF992A49990",
-15248 => x"C0C0BFF992A49980",
-15247 => x"C0C0BFF992A499F8",
-15246 => x"C0C0BFF992A49982",
-15245 => x"C0C0BFF992A49992",
-15244 => x"C0C0BFF992A49999",
-15243 => x"C0C0BFF992A499B0",
-15242 => x"C0C0BFF992A499A4",
-15241 => x"C0C0BFF992A499F9",
-15240 => x"C0C0BFF992A499C0",
-15239 => x"C0C0BFF992A4B090",
-15238 => x"C0C0BFF992A4B080",
-15237 => x"C0C0BFF992A4B0F8",
-15236 => x"C0C0BFF992A4B082",
-15235 => x"C0C0BFF992A4B092",
-15234 => x"C0C0BFF992A4B099",
-15233 => x"C0C0BFF992A4B0B0",
-15232 => x"C0C0BFF992A4B0A4",
-15231 => x"C0C0BFF992A4B0F9",
-15230 => x"C0C0BFF992A4B0C0",
-15229 => x"C0C0BFF992A4A490",
-15228 => x"C0C0BFF992A4A480",
-15227 => x"C0C0BFF992A4A4F8",
-15226 => x"C0C0BFF992A4A482",
-15225 => x"C0C0BFF992A4A492",
-15224 => x"C0C0BFF992A4A499",
-15223 => x"C0C0BFF992A4A4B0",
-15222 => x"C0C0BFF992A4A4A4",
-15221 => x"C0C0BFF992A4A4F9",
-15220 => x"C0C0BFF992A4A4C0",
-15219 => x"C0C0BFF992A4F990",
-15218 => x"C0C0BFF992A4F980",
-15217 => x"C0C0BFF992A4F9F8",
-15216 => x"C0C0BFF992A4F982",
-15215 => x"C0C0BFF992A4F992",
-15214 => x"C0C0BFF992A4F999",
-15213 => x"C0C0BFF992A4F9B0",
-15212 => x"C0C0BFF992A4F9A4",
-15211 => x"C0C0BFF992A4F9F9",
-15210 => x"C0C0BFF992A4F9C0",
-15209 => x"C0C0BFF992A4C090",
-15208 => x"C0C0BFF992A4C080",
-15207 => x"C0C0BFF992A4C0F8",
-15206 => x"C0C0BFF992A4C082",
-15205 => x"C0C0BFF992A4C092",
-15204 => x"C0C0BFF992A4C099",
-15203 => x"C0C0BFF992A4C0B0",
-15202 => x"C0C0BFF992A4C0A4",
-15201 => x"C0C0BFF992A4C0F9",
-15200 => x"C0C0BFF992A4C0C0",
-15199 => x"C0C0BFF992F99090",
-15198 => x"C0C0BFF992F99080",
-15197 => x"C0C0BFF992F990F8",
-15196 => x"C0C0BFF992F99082",
-15195 => x"C0C0BFF992F99092",
-15194 => x"C0C0BFF992F99099",
-15193 => x"C0C0BFF992F990B0",
-15192 => x"C0C0BFF992F990A4",
-15191 => x"C0C0BFF992F990F9",
-15190 => x"C0C0BFF992F990C0",
-15189 => x"C0C0BFF992F98090",
-15188 => x"C0C0BFF992F98080",
-15187 => x"C0C0BFF992F980F8",
-15186 => x"C0C0BFF992F98082",
-15185 => x"C0C0BFF992F98092",
-15184 => x"C0C0BFF992F98099",
-15183 => x"C0C0BFF992F980B0",
-15182 => x"C0C0BFF992F980A4",
-15181 => x"C0C0BFF992F980F9",
-15180 => x"C0C0BFF992F980C0",
-15179 => x"C0C0BFF992F9F890",
-15178 => x"C0C0BFF992F9F880",
-15177 => x"C0C0BFF992F9F8F8",
-15176 => x"C0C0BFF992F9F882",
-15175 => x"C0C0BFF992F9F892",
-15174 => x"C0C0BFF992F9F899",
-15173 => x"C0C0BFF992F9F8B0",
-15172 => x"C0C0BFF992F9F8A4",
-15171 => x"C0C0BFF992F9F8F9",
-15170 => x"C0C0BFF992F9F8C0",
-15169 => x"C0C0BFF992F98290",
-15168 => x"C0C0BFF992F98280",
-15167 => x"C0C0BFF992F982F8",
-15166 => x"C0C0BFF992F98282",
-15165 => x"C0C0BFF992F98292",
-15164 => x"C0C0BFF992F98299",
-15163 => x"C0C0BFF992F982B0",
-15162 => x"C0C0BFF992F982A4",
-15161 => x"C0C0BFF992F982F9",
-15160 => x"C0C0BFF992F982C0",
-15159 => x"C0C0BFF992F99290",
-15158 => x"C0C0BFF992F99280",
-15157 => x"C0C0BFF992F992F8",
-15156 => x"C0C0BFF992F99282",
-15155 => x"C0C0BFF992F99292",
-15154 => x"C0C0BFF992F99299",
-15153 => x"C0C0BFF992F992B0",
-15152 => x"C0C0BFF992F992A4",
-15151 => x"C0C0BFF992F992F9",
-15150 => x"C0C0BFF992F992C0",
-15149 => x"C0C0BFF992F99990",
-15148 => x"C0C0BFF992F99980",
-15147 => x"C0C0BFF992F999F8",
-15146 => x"C0C0BFF992F99982",
-15145 => x"C0C0BFF992F99992",
-15144 => x"C0C0BFF992F99999",
-15143 => x"C0C0BFF992F999B0",
-15142 => x"C0C0BFF992F999A4",
-15141 => x"C0C0BFF992F999F9",
-15140 => x"C0C0BFF992F999C0",
-15139 => x"C0C0BFF992F9B090",
-15138 => x"C0C0BFF992F9B080",
-15137 => x"C0C0BFF992F9B0F8",
-15136 => x"C0C0BFF992F9B082",
-15135 => x"C0C0BFF992F9B092",
-15134 => x"C0C0BFF992F9B099",
-15133 => x"C0C0BFF992F9B0B0",
-15132 => x"C0C0BFF992F9B0A4",
-15131 => x"C0C0BFF992F9B0F9",
-15130 => x"C0C0BFF992F9B0C0",
-15129 => x"C0C0BFF992F9A490",
-15128 => x"C0C0BFF992F9A480",
-15127 => x"C0C0BFF992F9A4F8",
-15126 => x"C0C0BFF992F9A482",
-15125 => x"C0C0BFF992F9A492",
-15124 => x"C0C0BFF992F9A499",
-15123 => x"C0C0BFF992F9A4B0",
-15122 => x"C0C0BFF992F9A4A4",
-15121 => x"C0C0BFF992F9A4F9",
-15120 => x"C0C0BFF992F9A4C0",
-15119 => x"C0C0BFF992F9F990",
-15118 => x"C0C0BFF992F9F980",
-15117 => x"C0C0BFF992F9F9F8",
-15116 => x"C0C0BFF992F9F982",
-15115 => x"C0C0BFF992F9F992",
-15114 => x"C0C0BFF992F9F999",
-15113 => x"C0C0BFF992F9F9B0",
-15112 => x"C0C0BFF992F9F9A4",
-15111 => x"C0C0BFF992F9F9F9",
-15110 => x"C0C0BFF992F9F9C0",
-15109 => x"C0C0BFF992F9C090",
-15108 => x"C0C0BFF992F9C080",
-15107 => x"C0C0BFF992F9C0F8",
-15106 => x"C0C0BFF992F9C082",
-15105 => x"C0C0BFF992F9C092",
-15104 => x"C0C0BFF992F9C099",
-15103 => x"C0C0BFF992F9C0B0",
-15102 => x"C0C0BFF992F9C0A4",
-15101 => x"C0C0BFF992F9C0F9",
-15100 => x"C0C0BFF992F9C0C0",
-15099 => x"C0C0BFF992C09090",
-15098 => x"C0C0BFF992C09080",
-15097 => x"C0C0BFF992C090F8",
-15096 => x"C0C0BFF992C09082",
-15095 => x"C0C0BFF992C09092",
-15094 => x"C0C0BFF992C09099",
-15093 => x"C0C0BFF992C090B0",
-15092 => x"C0C0BFF992C090A4",
-15091 => x"C0C0BFF992C090F9",
-15090 => x"C0C0BFF992C090C0",
-15089 => x"C0C0BFF992C08090",
-15088 => x"C0C0BFF992C08080",
-15087 => x"C0C0BFF992C080F8",
-15086 => x"C0C0BFF992C08082",
-15085 => x"C0C0BFF992C08092",
-15084 => x"C0C0BFF992C08099",
-15083 => x"C0C0BFF992C080B0",
-15082 => x"C0C0BFF992C080A4",
-15081 => x"C0C0BFF992C080F9",
-15080 => x"C0C0BFF992C080C0",
-15079 => x"C0C0BFF992C0F890",
-15078 => x"C0C0BFF992C0F880",
-15077 => x"C0C0BFF992C0F8F8",
-15076 => x"C0C0BFF992C0F882",
-15075 => x"C0C0BFF992C0F892",
-15074 => x"C0C0BFF992C0F899",
-15073 => x"C0C0BFF992C0F8B0",
-15072 => x"C0C0BFF992C0F8A4",
-15071 => x"C0C0BFF992C0F8F9",
-15070 => x"C0C0BFF992C0F8C0",
-15069 => x"C0C0BFF992C08290",
-15068 => x"C0C0BFF992C08280",
-15067 => x"C0C0BFF992C082F8",
-15066 => x"C0C0BFF992C08282",
-15065 => x"C0C0BFF992C08292",
-15064 => x"C0C0BFF992C08299",
-15063 => x"C0C0BFF992C082B0",
-15062 => x"C0C0BFF992C082A4",
-15061 => x"C0C0BFF992C082F9",
-15060 => x"C0C0BFF992C082C0",
-15059 => x"C0C0BFF992C09290",
-15058 => x"C0C0BFF992C09280",
-15057 => x"C0C0BFF992C092F8",
-15056 => x"C0C0BFF992C09282",
-15055 => x"C0C0BFF992C09292",
-15054 => x"C0C0BFF992C09299",
-15053 => x"C0C0BFF992C092B0",
-15052 => x"C0C0BFF992C092A4",
-15051 => x"C0C0BFF992C092F9",
-15050 => x"C0C0BFF992C092C0",
-15049 => x"C0C0BFF992C09990",
-15048 => x"C0C0BFF992C09980",
-15047 => x"C0C0BFF992C099F8",
-15046 => x"C0C0BFF992C09982",
-15045 => x"C0C0BFF992C09992",
-15044 => x"C0C0BFF992C09999",
-15043 => x"C0C0BFF992C099B0",
-15042 => x"C0C0BFF992C099A4",
-15041 => x"C0C0BFF992C099F9",
-15040 => x"C0C0BFF992C099C0",
-15039 => x"C0C0BFF992C0B090",
-15038 => x"C0C0BFF992C0B080",
-15037 => x"C0C0BFF992C0B0F8",
-15036 => x"C0C0BFF992C0B082",
-15035 => x"C0C0BFF992C0B092",
-15034 => x"C0C0BFF992C0B099",
-15033 => x"C0C0BFF992C0B0B0",
-15032 => x"C0C0BFF992C0B0A4",
-15031 => x"C0C0BFF992C0B0F9",
-15030 => x"C0C0BFF992C0B0C0",
-15029 => x"C0C0BFF992C0A490",
-15028 => x"C0C0BFF992C0A480",
-15027 => x"C0C0BFF992C0A4F8",
-15026 => x"C0C0BFF992C0A482",
-15025 => x"C0C0BFF992C0A492",
-15024 => x"C0C0BFF992C0A499",
-15023 => x"C0C0BFF992C0A4B0",
-15022 => x"C0C0BFF992C0A4A4",
-15021 => x"C0C0BFF992C0A4F9",
-15020 => x"C0C0BFF992C0A4C0",
-15019 => x"C0C0BFF992C0F990",
-15018 => x"C0C0BFF992C0F980",
-15017 => x"C0C0BFF992C0F9F8",
-15016 => x"C0C0BFF992C0F982",
-15015 => x"C0C0BFF992C0F992",
-15014 => x"C0C0BFF992C0F999",
-15013 => x"C0C0BFF992C0F9B0",
-15012 => x"C0C0BFF992C0F9A4",
-15011 => x"C0C0BFF992C0F9F9",
-15010 => x"C0C0BFF992C0F9C0",
-15009 => x"C0C0BFF992C0C090",
-15008 => x"C0C0BFF992C0C080",
-15007 => x"C0C0BFF992C0C0F8",
-15006 => x"C0C0BFF992C0C082",
-15005 => x"C0C0BFF992C0C092",
-15004 => x"C0C0BFF992C0C099",
-15003 => x"C0C0BFF992C0C0B0",
-15002 => x"C0C0BFF992C0C0A4",
-15001 => x"C0C0BFF992C0C0F9",
-15000 => x"C0C0BFF992C0C0C0",
-14999 => x"C0C0BFF999909090",
-14998 => x"C0C0BFF999909080",
-14997 => x"C0C0BFF9999090F8",
-14996 => x"C0C0BFF999909082",
-14995 => x"C0C0BFF999909092",
-14994 => x"C0C0BFF999909099",
-14993 => x"C0C0BFF9999090B0",
-14992 => x"C0C0BFF9999090A4",
-14991 => x"C0C0BFF9999090F9",
-14990 => x"C0C0BFF9999090C0",
-14989 => x"C0C0BFF999908090",
-14988 => x"C0C0BFF999908080",
-14987 => x"C0C0BFF9999080F8",
-14986 => x"C0C0BFF999908082",
-14985 => x"C0C0BFF999908092",
-14984 => x"C0C0BFF999908099",
-14983 => x"C0C0BFF9999080B0",
-14982 => x"C0C0BFF9999080A4",
-14981 => x"C0C0BFF9999080F9",
-14980 => x"C0C0BFF9999080C0",
-14979 => x"C0C0BFF99990F890",
-14978 => x"C0C0BFF99990F880",
-14977 => x"C0C0BFF99990F8F8",
-14976 => x"C0C0BFF99990F882",
-14975 => x"C0C0BFF99990F892",
-14974 => x"C0C0BFF99990F899",
-14973 => x"C0C0BFF99990F8B0",
-14972 => x"C0C0BFF99990F8A4",
-14971 => x"C0C0BFF99990F8F9",
-14970 => x"C0C0BFF99990F8C0",
-14969 => x"C0C0BFF999908290",
-14968 => x"C0C0BFF999908280",
-14967 => x"C0C0BFF9999082F8",
-14966 => x"C0C0BFF999908282",
-14965 => x"C0C0BFF999908292",
-14964 => x"C0C0BFF999908299",
-14963 => x"C0C0BFF9999082B0",
-14962 => x"C0C0BFF9999082A4",
-14961 => x"C0C0BFF9999082F9",
-14960 => x"C0C0BFF9999082C0",
-14959 => x"C0C0BFF999909290",
-14958 => x"C0C0BFF999909280",
-14957 => x"C0C0BFF9999092F8",
-14956 => x"C0C0BFF999909282",
-14955 => x"C0C0BFF999909292",
-14954 => x"C0C0BFF999909299",
-14953 => x"C0C0BFF9999092B0",
-14952 => x"C0C0BFF9999092A4",
-14951 => x"C0C0BFF9999092F9",
-14950 => x"C0C0BFF9999092C0",
-14949 => x"C0C0BFF999909990",
-14948 => x"C0C0BFF999909980",
-14947 => x"C0C0BFF9999099F8",
-14946 => x"C0C0BFF999909982",
-14945 => x"C0C0BFF999909992",
-14944 => x"C0C0BFF999909999",
-14943 => x"C0C0BFF9999099B0",
-14942 => x"C0C0BFF9999099A4",
-14941 => x"C0C0BFF9999099F9",
-14940 => x"C0C0BFF9999099C0",
-14939 => x"C0C0BFF99990B090",
-14938 => x"C0C0BFF99990B080",
-14937 => x"C0C0BFF99990B0F8",
-14936 => x"C0C0BFF99990B082",
-14935 => x"C0C0BFF99990B092",
-14934 => x"C0C0BFF99990B099",
-14933 => x"C0C0BFF99990B0B0",
-14932 => x"C0C0BFF99990B0A4",
-14931 => x"C0C0BFF99990B0F9",
-14930 => x"C0C0BFF99990B0C0",
-14929 => x"C0C0BFF99990A490",
-14928 => x"C0C0BFF99990A480",
-14927 => x"C0C0BFF99990A4F8",
-14926 => x"C0C0BFF99990A482",
-14925 => x"C0C0BFF99990A492",
-14924 => x"C0C0BFF99990A499",
-14923 => x"C0C0BFF99990A4B0",
-14922 => x"C0C0BFF99990A4A4",
-14921 => x"C0C0BFF99990A4F9",
-14920 => x"C0C0BFF99990A4C0",
-14919 => x"C0C0BFF99990F990",
-14918 => x"C0C0BFF99990F980",
-14917 => x"C0C0BFF99990F9F8",
-14916 => x"C0C0BFF99990F982",
-14915 => x"C0C0BFF99990F992",
-14914 => x"C0C0BFF99990F999",
-14913 => x"C0C0BFF99990F9B0",
-14912 => x"C0C0BFF99990F9A4",
-14911 => x"C0C0BFF99990F9F9",
-14910 => x"C0C0BFF99990F9C0",
-14909 => x"C0C0BFF99990C090",
-14908 => x"C0C0BFF99990C080",
-14907 => x"C0C0BFF99990C0F8",
-14906 => x"C0C0BFF99990C082",
-14905 => x"C0C0BFF99990C092",
-14904 => x"C0C0BFF99990C099",
-14903 => x"C0C0BFF99990C0B0",
-14902 => x"C0C0BFF99990C0A4",
-14901 => x"C0C0BFF99990C0F9",
-14900 => x"C0C0BFF99990C0C0",
-14899 => x"C0C0BFF999809090",
-14898 => x"C0C0BFF999809080",
-14897 => x"C0C0BFF9998090F8",
-14896 => x"C0C0BFF999809082",
-14895 => x"C0C0BFF999809092",
-14894 => x"C0C0BFF999809099",
-14893 => x"C0C0BFF9998090B0",
-14892 => x"C0C0BFF9998090A4",
-14891 => x"C0C0BFF9998090F9",
-14890 => x"C0C0BFF9998090C0",
-14889 => x"C0C0BFF999808090",
-14888 => x"C0C0BFF999808080",
-14887 => x"C0C0BFF9998080F8",
-14886 => x"C0C0BFF999808082",
-14885 => x"C0C0BFF999808092",
-14884 => x"C0C0BFF999808099",
-14883 => x"C0C0BFF9998080B0",
-14882 => x"C0C0BFF9998080A4",
-14881 => x"C0C0BFF9998080F9",
-14880 => x"C0C0BFF9998080C0",
-14879 => x"C0C0BFF99980F890",
-14878 => x"C0C0BFF99980F880",
-14877 => x"C0C0BFF99980F8F8",
-14876 => x"C0C0BFF99980F882",
-14875 => x"C0C0BFF99980F892",
-14874 => x"C0C0BFF99980F899",
-14873 => x"C0C0BFF99980F8B0",
-14872 => x"C0C0BFF99980F8A4",
-14871 => x"C0C0BFF99980F8F9",
-14870 => x"C0C0BFF99980F8C0",
-14869 => x"C0C0BFF999808290",
-14868 => x"C0C0BFF999808280",
-14867 => x"C0C0BFF9998082F8",
-14866 => x"C0C0BFF999808282",
-14865 => x"C0C0BFF999808292",
-14864 => x"C0C0BFF999808299",
-14863 => x"C0C0BFF9998082B0",
-14862 => x"C0C0BFF9998082A4",
-14861 => x"C0C0BFF9998082F9",
-14860 => x"C0C0BFF9998082C0",
-14859 => x"C0C0BFF999809290",
-14858 => x"C0C0BFF999809280",
-14857 => x"C0C0BFF9998092F8",
-14856 => x"C0C0BFF999809282",
-14855 => x"C0C0BFF999809292",
-14854 => x"C0C0BFF999809299",
-14853 => x"C0C0BFF9998092B0",
-14852 => x"C0C0BFF9998092A4",
-14851 => x"C0C0BFF9998092F9",
-14850 => x"C0C0BFF9998092C0",
-14849 => x"C0C0BFF999809990",
-14848 => x"C0C0BFF999809980",
-14847 => x"C0C0BFF9998099F8",
-14846 => x"C0C0BFF999809982",
-14845 => x"C0C0BFF999809992",
-14844 => x"C0C0BFF999809999",
-14843 => x"C0C0BFF9998099B0",
-14842 => x"C0C0BFF9998099A4",
-14841 => x"C0C0BFF9998099F9",
-14840 => x"C0C0BFF9998099C0",
-14839 => x"C0C0BFF99980B090",
-14838 => x"C0C0BFF99980B080",
-14837 => x"C0C0BFF99980B0F8",
-14836 => x"C0C0BFF99980B082",
-14835 => x"C0C0BFF99980B092",
-14834 => x"C0C0BFF99980B099",
-14833 => x"C0C0BFF99980B0B0",
-14832 => x"C0C0BFF99980B0A4",
-14831 => x"C0C0BFF99980B0F9",
-14830 => x"C0C0BFF99980B0C0",
-14829 => x"C0C0BFF99980A490",
-14828 => x"C0C0BFF99980A480",
-14827 => x"C0C0BFF99980A4F8",
-14826 => x"C0C0BFF99980A482",
-14825 => x"C0C0BFF99980A492",
-14824 => x"C0C0BFF99980A499",
-14823 => x"C0C0BFF99980A4B0",
-14822 => x"C0C0BFF99980A4A4",
-14821 => x"C0C0BFF99980A4F9",
-14820 => x"C0C0BFF99980A4C0",
-14819 => x"C0C0BFF99980F990",
-14818 => x"C0C0BFF99980F980",
-14817 => x"C0C0BFF99980F9F8",
-14816 => x"C0C0BFF99980F982",
-14815 => x"C0C0BFF99980F992",
-14814 => x"C0C0BFF99980F999",
-14813 => x"C0C0BFF99980F9B0",
-14812 => x"C0C0BFF99980F9A4",
-14811 => x"C0C0BFF99980F9F9",
-14810 => x"C0C0BFF99980F9C0",
-14809 => x"C0C0BFF99980C090",
-14808 => x"C0C0BFF99980C080",
-14807 => x"C0C0BFF99980C0F8",
-14806 => x"C0C0BFF99980C082",
-14805 => x"C0C0BFF99980C092",
-14804 => x"C0C0BFF99980C099",
-14803 => x"C0C0BFF99980C0B0",
-14802 => x"C0C0BFF99980C0A4",
-14801 => x"C0C0BFF99980C0F9",
-14800 => x"C0C0BFF99980C0C0",
-14799 => x"C0C0BFF999F89090",
-14798 => x"C0C0BFF999F89080",
-14797 => x"C0C0BFF999F890F8",
-14796 => x"C0C0BFF999F89082",
-14795 => x"C0C0BFF999F89092",
-14794 => x"C0C0BFF999F89099",
-14793 => x"C0C0BFF999F890B0",
-14792 => x"C0C0BFF999F890A4",
-14791 => x"C0C0BFF999F890F9",
-14790 => x"C0C0BFF999F890C0",
-14789 => x"C0C0BFF999F88090",
-14788 => x"C0C0BFF999F88080",
-14787 => x"C0C0BFF999F880F8",
-14786 => x"C0C0BFF999F88082",
-14785 => x"C0C0BFF999F88092",
-14784 => x"C0C0BFF999F88099",
-14783 => x"C0C0BFF999F880B0",
-14782 => x"C0C0BFF999F880A4",
-14781 => x"C0C0BFF999F880F9",
-14780 => x"C0C0BFF999F880C0",
-14779 => x"C0C0BFF999F8F890",
-14778 => x"C0C0BFF999F8F880",
-14777 => x"C0C0BFF999F8F8F8",
-14776 => x"C0C0BFF999F8F882",
-14775 => x"C0C0BFF999F8F892",
-14774 => x"C0C0BFF999F8F899",
-14773 => x"C0C0BFF999F8F8B0",
-14772 => x"C0C0BFF999F8F8A4",
-14771 => x"C0C0BFF999F8F8F9",
-14770 => x"C0C0BFF999F8F8C0",
-14769 => x"C0C0BFF999F88290",
-14768 => x"C0C0BFF999F88280",
-14767 => x"C0C0BFF999F882F8",
-14766 => x"C0C0BFF999F88282",
-14765 => x"C0C0BFF999F88292",
-14764 => x"C0C0BFF999F88299",
-14763 => x"C0C0BFF999F882B0",
-14762 => x"C0C0BFF999F882A4",
-14761 => x"C0C0BFF999F882F9",
-14760 => x"C0C0BFF999F882C0",
-14759 => x"C0C0BFF999F89290",
-14758 => x"C0C0BFF999F89280",
-14757 => x"C0C0BFF999F892F8",
-14756 => x"C0C0BFF999F89282",
-14755 => x"C0C0BFF999F89292",
-14754 => x"C0C0BFF999F89299",
-14753 => x"C0C0BFF999F892B0",
-14752 => x"C0C0BFF999F892A4",
-14751 => x"C0C0BFF999F892F9",
-14750 => x"C0C0BFF999F892C0",
-14749 => x"C0C0BFF999F89990",
-14748 => x"C0C0BFF999F89980",
-14747 => x"C0C0BFF999F899F8",
-14746 => x"C0C0BFF999F89982",
-14745 => x"C0C0BFF999F89992",
-14744 => x"C0C0BFF999F89999",
-14743 => x"C0C0BFF999F899B0",
-14742 => x"C0C0BFF999F899A4",
-14741 => x"C0C0BFF999F899F9",
-14740 => x"C0C0BFF999F899C0",
-14739 => x"C0C0BFF999F8B090",
-14738 => x"C0C0BFF999F8B080",
-14737 => x"C0C0BFF999F8B0F8",
-14736 => x"C0C0BFF999F8B082",
-14735 => x"C0C0BFF999F8B092",
-14734 => x"C0C0BFF999F8B099",
-14733 => x"C0C0BFF999F8B0B0",
-14732 => x"C0C0BFF999F8B0A4",
-14731 => x"C0C0BFF999F8B0F9",
-14730 => x"C0C0BFF999F8B0C0",
-14729 => x"C0C0BFF999F8A490",
-14728 => x"C0C0BFF999F8A480",
-14727 => x"C0C0BFF999F8A4F8",
-14726 => x"C0C0BFF999F8A482",
-14725 => x"C0C0BFF999F8A492",
-14724 => x"C0C0BFF999F8A499",
-14723 => x"C0C0BFF999F8A4B0",
-14722 => x"C0C0BFF999F8A4A4",
-14721 => x"C0C0BFF999F8A4F9",
-14720 => x"C0C0BFF999F8A4C0",
-14719 => x"C0C0BFF999F8F990",
-14718 => x"C0C0BFF999F8F980",
-14717 => x"C0C0BFF999F8F9F8",
-14716 => x"C0C0BFF999F8F982",
-14715 => x"C0C0BFF999F8F992",
-14714 => x"C0C0BFF999F8F999",
-14713 => x"C0C0BFF999F8F9B0",
-14712 => x"C0C0BFF999F8F9A4",
-14711 => x"C0C0BFF999F8F9F9",
-14710 => x"C0C0BFF999F8F9C0",
-14709 => x"C0C0BFF999F8C090",
-14708 => x"C0C0BFF999F8C080",
-14707 => x"C0C0BFF999F8C0F8",
-14706 => x"C0C0BFF999F8C082",
-14705 => x"C0C0BFF999F8C092",
-14704 => x"C0C0BFF999F8C099",
-14703 => x"C0C0BFF999F8C0B0",
-14702 => x"C0C0BFF999F8C0A4",
-14701 => x"C0C0BFF999F8C0F9",
-14700 => x"C0C0BFF999F8C0C0",
-14699 => x"C0C0BFF999829090",
-14698 => x"C0C0BFF999829080",
-14697 => x"C0C0BFF9998290F8",
-14696 => x"C0C0BFF999829082",
-14695 => x"C0C0BFF999829092",
-14694 => x"C0C0BFF999829099",
-14693 => x"C0C0BFF9998290B0",
-14692 => x"C0C0BFF9998290A4",
-14691 => x"C0C0BFF9998290F9",
-14690 => x"C0C0BFF9998290C0",
-14689 => x"C0C0BFF999828090",
-14688 => x"C0C0BFF999828080",
-14687 => x"C0C0BFF9998280F8",
-14686 => x"C0C0BFF999828082",
-14685 => x"C0C0BFF999828092",
-14684 => x"C0C0BFF999828099",
-14683 => x"C0C0BFF9998280B0",
-14682 => x"C0C0BFF9998280A4",
-14681 => x"C0C0BFF9998280F9",
-14680 => x"C0C0BFF9998280C0",
-14679 => x"C0C0BFF99982F890",
-14678 => x"C0C0BFF99982F880",
-14677 => x"C0C0BFF99982F8F8",
-14676 => x"C0C0BFF99982F882",
-14675 => x"C0C0BFF99982F892",
-14674 => x"C0C0BFF99982F899",
-14673 => x"C0C0BFF99982F8B0",
-14672 => x"C0C0BFF99982F8A4",
-14671 => x"C0C0BFF99982F8F9",
-14670 => x"C0C0BFF99982F8C0",
-14669 => x"C0C0BFF999828290",
-14668 => x"C0C0BFF999828280",
-14667 => x"C0C0BFF9998282F8",
-14666 => x"C0C0BFF999828282",
-14665 => x"C0C0BFF999828292",
-14664 => x"C0C0BFF999828299",
-14663 => x"C0C0BFF9998282B0",
-14662 => x"C0C0BFF9998282A4",
-14661 => x"C0C0BFF9998282F9",
-14660 => x"C0C0BFF9998282C0",
-14659 => x"C0C0BFF999829290",
-14658 => x"C0C0BFF999829280",
-14657 => x"C0C0BFF9998292F8",
-14656 => x"C0C0BFF999829282",
-14655 => x"C0C0BFF999829292",
-14654 => x"C0C0BFF999829299",
-14653 => x"C0C0BFF9998292B0",
-14652 => x"C0C0BFF9998292A4",
-14651 => x"C0C0BFF9998292F9",
-14650 => x"C0C0BFF9998292C0",
-14649 => x"C0C0BFF999829990",
-14648 => x"C0C0BFF999829980",
-14647 => x"C0C0BFF9998299F8",
-14646 => x"C0C0BFF999829982",
-14645 => x"C0C0BFF999829992",
-14644 => x"C0C0BFF999829999",
-14643 => x"C0C0BFF9998299B0",
-14642 => x"C0C0BFF9998299A4",
-14641 => x"C0C0BFF9998299F9",
-14640 => x"C0C0BFF9998299C0",
-14639 => x"C0C0BFF99982B090",
-14638 => x"C0C0BFF99982B080",
-14637 => x"C0C0BFF99982B0F8",
-14636 => x"C0C0BFF99982B082",
-14635 => x"C0C0BFF99982B092",
-14634 => x"C0C0BFF99982B099",
-14633 => x"C0C0BFF99982B0B0",
-14632 => x"C0C0BFF99982B0A4",
-14631 => x"C0C0BFF99982B0F9",
-14630 => x"C0C0BFF99982B0C0",
-14629 => x"C0C0BFF99982A490",
-14628 => x"C0C0BFF99982A480",
-14627 => x"C0C0BFF99982A4F8",
-14626 => x"C0C0BFF99982A482",
-14625 => x"C0C0BFF99982A492",
-14624 => x"C0C0BFF99982A499",
-14623 => x"C0C0BFF99982A4B0",
-14622 => x"C0C0BFF99982A4A4",
-14621 => x"C0C0BFF99982A4F9",
-14620 => x"C0C0BFF99982A4C0",
-14619 => x"C0C0BFF99982F990",
-14618 => x"C0C0BFF99982F980",
-14617 => x"C0C0BFF99982F9F8",
-14616 => x"C0C0BFF99982F982",
-14615 => x"C0C0BFF99982F992",
-14614 => x"C0C0BFF99982F999",
-14613 => x"C0C0BFF99982F9B0",
-14612 => x"C0C0BFF99982F9A4",
-14611 => x"C0C0BFF99982F9F9",
-14610 => x"C0C0BFF99982F9C0",
-14609 => x"C0C0BFF99982C090",
-14608 => x"C0C0BFF99982C080",
-14607 => x"C0C0BFF99982C0F8",
-14606 => x"C0C0BFF99982C082",
-14605 => x"C0C0BFF99982C092",
-14604 => x"C0C0BFF99982C099",
-14603 => x"C0C0BFF99982C0B0",
-14602 => x"C0C0BFF99982C0A4",
-14601 => x"C0C0BFF99982C0F9",
-14600 => x"C0C0BFF99982C0C0",
-14599 => x"C0C0BFF999929090",
-14598 => x"C0C0BFF999929080",
-14597 => x"C0C0BFF9999290F8",
-14596 => x"C0C0BFF999929082",
-14595 => x"C0C0BFF999929092",
-14594 => x"C0C0BFF999929099",
-14593 => x"C0C0BFF9999290B0",
-14592 => x"C0C0BFF9999290A4",
-14591 => x"C0C0BFF9999290F9",
-14590 => x"C0C0BFF9999290C0",
-14589 => x"C0C0BFF999928090",
-14588 => x"C0C0BFF999928080",
-14587 => x"C0C0BFF9999280F8",
-14586 => x"C0C0BFF999928082",
-14585 => x"C0C0BFF999928092",
-14584 => x"C0C0BFF999928099",
-14583 => x"C0C0BFF9999280B0",
-14582 => x"C0C0BFF9999280A4",
-14581 => x"C0C0BFF9999280F9",
-14580 => x"C0C0BFF9999280C0",
-14579 => x"C0C0BFF99992F890",
-14578 => x"C0C0BFF99992F880",
-14577 => x"C0C0BFF99992F8F8",
-14576 => x"C0C0BFF99992F882",
-14575 => x"C0C0BFF99992F892",
-14574 => x"C0C0BFF99992F899",
-14573 => x"C0C0BFF99992F8B0",
-14572 => x"C0C0BFF99992F8A4",
-14571 => x"C0C0BFF99992F8F9",
-14570 => x"C0C0BFF99992F8C0",
-14569 => x"C0C0BFF999928290",
-14568 => x"C0C0BFF999928280",
-14567 => x"C0C0BFF9999282F8",
-14566 => x"C0C0BFF999928282",
-14565 => x"C0C0BFF999928292",
-14564 => x"C0C0BFF999928299",
-14563 => x"C0C0BFF9999282B0",
-14562 => x"C0C0BFF9999282A4",
-14561 => x"C0C0BFF9999282F9",
-14560 => x"C0C0BFF9999282C0",
-14559 => x"C0C0BFF999929290",
-14558 => x"C0C0BFF999929280",
-14557 => x"C0C0BFF9999292F8",
-14556 => x"C0C0BFF999929282",
-14555 => x"C0C0BFF999929292",
-14554 => x"C0C0BFF999929299",
-14553 => x"C0C0BFF9999292B0",
-14552 => x"C0C0BFF9999292A4",
-14551 => x"C0C0BFF9999292F9",
-14550 => x"C0C0BFF9999292C0",
-14549 => x"C0C0BFF999929990",
-14548 => x"C0C0BFF999929980",
-14547 => x"C0C0BFF9999299F8",
-14546 => x"C0C0BFF999929982",
-14545 => x"C0C0BFF999929992",
-14544 => x"C0C0BFF999929999",
-14543 => x"C0C0BFF9999299B0",
-14542 => x"C0C0BFF9999299A4",
-14541 => x"C0C0BFF9999299F9",
-14540 => x"C0C0BFF9999299C0",
-14539 => x"C0C0BFF99992B090",
-14538 => x"C0C0BFF99992B080",
-14537 => x"C0C0BFF99992B0F8",
-14536 => x"C0C0BFF99992B082",
-14535 => x"C0C0BFF99992B092",
-14534 => x"C0C0BFF99992B099",
-14533 => x"C0C0BFF99992B0B0",
-14532 => x"C0C0BFF99992B0A4",
-14531 => x"C0C0BFF99992B0F9",
-14530 => x"C0C0BFF99992B0C0",
-14529 => x"C0C0BFF99992A490",
-14528 => x"C0C0BFF99992A480",
-14527 => x"C0C0BFF99992A4F8",
-14526 => x"C0C0BFF99992A482",
-14525 => x"C0C0BFF99992A492",
-14524 => x"C0C0BFF99992A499",
-14523 => x"C0C0BFF99992A4B0",
-14522 => x"C0C0BFF99992A4A4",
-14521 => x"C0C0BFF99992A4F9",
-14520 => x"C0C0BFF99992A4C0",
-14519 => x"C0C0BFF99992F990",
-14518 => x"C0C0BFF99992F980",
-14517 => x"C0C0BFF99992F9F8",
-14516 => x"C0C0BFF99992F982",
-14515 => x"C0C0BFF99992F992",
-14514 => x"C0C0BFF99992F999",
-14513 => x"C0C0BFF99992F9B0",
-14512 => x"C0C0BFF99992F9A4",
-14511 => x"C0C0BFF99992F9F9",
-14510 => x"C0C0BFF99992F9C0",
-14509 => x"C0C0BFF99992C090",
-14508 => x"C0C0BFF99992C080",
-14507 => x"C0C0BFF99992C0F8",
-14506 => x"C0C0BFF99992C082",
-14505 => x"C0C0BFF99992C092",
-14504 => x"C0C0BFF99992C099",
-14503 => x"C0C0BFF99992C0B0",
-14502 => x"C0C0BFF99992C0A4",
-14501 => x"C0C0BFF99992C0F9",
-14500 => x"C0C0BFF99992C0C0",
-14499 => x"C0C0BFF999999090",
-14498 => x"C0C0BFF999999080",
-14497 => x"C0C0BFF9999990F8",
-14496 => x"C0C0BFF999999082",
-14495 => x"C0C0BFF999999092",
-14494 => x"C0C0BFF999999099",
-14493 => x"C0C0BFF9999990B0",
-14492 => x"C0C0BFF9999990A4",
-14491 => x"C0C0BFF9999990F9",
-14490 => x"C0C0BFF9999990C0",
-14489 => x"C0C0BFF999998090",
-14488 => x"C0C0BFF999998080",
-14487 => x"C0C0BFF9999980F8",
-14486 => x"C0C0BFF999998082",
-14485 => x"C0C0BFF999998092",
-14484 => x"C0C0BFF999998099",
-14483 => x"C0C0BFF9999980B0",
-14482 => x"C0C0BFF9999980A4",
-14481 => x"C0C0BFF9999980F9",
-14480 => x"C0C0BFF9999980C0",
-14479 => x"C0C0BFF99999F890",
-14478 => x"C0C0BFF99999F880",
-14477 => x"C0C0BFF99999F8F8",
-14476 => x"C0C0BFF99999F882",
-14475 => x"C0C0BFF99999F892",
-14474 => x"C0C0BFF99999F899",
-14473 => x"C0C0BFF99999F8B0",
-14472 => x"C0C0BFF99999F8A4",
-14471 => x"C0C0BFF99999F8F9",
-14470 => x"C0C0BFF99999F8C0",
-14469 => x"C0C0BFF999998290",
-14468 => x"C0C0BFF999998280",
-14467 => x"C0C0BFF9999982F8",
-14466 => x"C0C0BFF999998282",
-14465 => x"C0C0BFF999998292",
-14464 => x"C0C0BFF999998299",
-14463 => x"C0C0BFF9999982B0",
-14462 => x"C0C0BFF9999982A4",
-14461 => x"C0C0BFF9999982F9",
-14460 => x"C0C0BFF9999982C0",
-14459 => x"C0C0BFF999999290",
-14458 => x"C0C0BFF999999280",
-14457 => x"C0C0BFF9999992F8",
-14456 => x"C0C0BFF999999282",
-14455 => x"C0C0BFF999999292",
-14454 => x"C0C0BFF999999299",
-14453 => x"C0C0BFF9999992B0",
-14452 => x"C0C0BFF9999992A4",
-14451 => x"C0C0BFF9999992F9",
-14450 => x"C0C0BFF9999992C0",
-14449 => x"C0C0BFF999999990",
-14448 => x"C0C0BFF999999980",
-14447 => x"C0C0BFF9999999F8",
-14446 => x"C0C0BFF999999982",
-14445 => x"C0C0BFF999999992",
-14444 => x"C0C0BFF999999999",
-14443 => x"C0C0BFF9999999B0",
-14442 => x"C0C0BFF9999999A4",
-14441 => x"C0C0BFF9999999F9",
-14440 => x"C0C0BFF9999999C0",
-14439 => x"C0C0BFF99999B090",
-14438 => x"C0C0BFF99999B080",
-14437 => x"C0C0BFF99999B0F8",
-14436 => x"C0C0BFF99999B082",
-14435 => x"C0C0BFF99999B092",
-14434 => x"C0C0BFF99999B099",
-14433 => x"C0C0BFF99999B0B0",
-14432 => x"C0C0BFF99999B0A4",
-14431 => x"C0C0BFF99999B0F9",
-14430 => x"C0C0BFF99999B0C0",
-14429 => x"C0C0BFF99999A490",
-14428 => x"C0C0BFF99999A480",
-14427 => x"C0C0BFF99999A4F8",
-14426 => x"C0C0BFF99999A482",
-14425 => x"C0C0BFF99999A492",
-14424 => x"C0C0BFF99999A499",
-14423 => x"C0C0BFF99999A4B0",
-14422 => x"C0C0BFF99999A4A4",
-14421 => x"C0C0BFF99999A4F9",
-14420 => x"C0C0BFF99999A4C0",
-14419 => x"C0C0BFF99999F990",
-14418 => x"C0C0BFF99999F980",
-14417 => x"C0C0BFF99999F9F8",
-14416 => x"C0C0BFF99999F982",
-14415 => x"C0C0BFF99999F992",
-14414 => x"C0C0BFF99999F999",
-14413 => x"C0C0BFF99999F9B0",
-14412 => x"C0C0BFF99999F9A4",
-14411 => x"C0C0BFF99999F9F9",
-14410 => x"C0C0BFF99999F9C0",
-14409 => x"C0C0BFF99999C090",
-14408 => x"C0C0BFF99999C080",
-14407 => x"C0C0BFF99999C0F8",
-14406 => x"C0C0BFF99999C082",
-14405 => x"C0C0BFF99999C092",
-14404 => x"C0C0BFF99999C099",
-14403 => x"C0C0BFF99999C0B0",
-14402 => x"C0C0BFF99999C0A4",
-14401 => x"C0C0BFF99999C0F9",
-14400 => x"C0C0BFF99999C0C0",
-14399 => x"C0C0BFF999B09090",
-14398 => x"C0C0BFF999B09080",
-14397 => x"C0C0BFF999B090F8",
-14396 => x"C0C0BFF999B09082",
-14395 => x"C0C0BFF999B09092",
-14394 => x"C0C0BFF999B09099",
-14393 => x"C0C0BFF999B090B0",
-14392 => x"C0C0BFF999B090A4",
-14391 => x"C0C0BFF999B090F9",
-14390 => x"C0C0BFF999B090C0",
-14389 => x"C0C0BFF999B08090",
-14388 => x"C0C0BFF999B08080",
-14387 => x"C0C0BFF999B080F8",
-14386 => x"C0C0BFF999B08082",
-14385 => x"C0C0BFF999B08092",
-14384 => x"C0C0BFF999B08099",
-14383 => x"C0C0BFF999B080B0",
-14382 => x"C0C0BFF999B080A4",
-14381 => x"C0C0BFF999B080F9",
-14380 => x"C0C0BFF999B080C0",
-14379 => x"C0C0BFF999B0F890",
-14378 => x"C0C0BFF999B0F880",
-14377 => x"C0C0BFF999B0F8F8",
-14376 => x"C0C0BFF999B0F882",
-14375 => x"C0C0BFF999B0F892",
-14374 => x"C0C0BFF999B0F899",
-14373 => x"C0C0BFF999B0F8B0",
-14372 => x"C0C0BFF999B0F8A4",
-14371 => x"C0C0BFF999B0F8F9",
-14370 => x"C0C0BFF999B0F8C0",
-14369 => x"C0C0BFF999B08290",
-14368 => x"C0C0BFF999B08280",
-14367 => x"C0C0BFF999B082F8",
-14366 => x"C0C0BFF999B08282",
-14365 => x"C0C0BFF999B08292",
-14364 => x"C0C0BFF999B08299",
-14363 => x"C0C0BFF999B082B0",
-14362 => x"C0C0BFF999B082A4",
-14361 => x"C0C0BFF999B082F9",
-14360 => x"C0C0BFF999B082C0",
-14359 => x"C0C0BFF999B09290",
-14358 => x"C0C0BFF999B09280",
-14357 => x"C0C0BFF999B092F8",
-14356 => x"C0C0BFF999B09282",
-14355 => x"C0C0BFF999B09292",
-14354 => x"C0C0BFF999B09299",
-14353 => x"C0C0BFF999B092B0",
-14352 => x"C0C0BFF999B092A4",
-14351 => x"C0C0BFF999B092F9",
-14350 => x"C0C0BFF999B092C0",
-14349 => x"C0C0BFF999B09990",
-14348 => x"C0C0BFF999B09980",
-14347 => x"C0C0BFF999B099F8",
-14346 => x"C0C0BFF999B09982",
-14345 => x"C0C0BFF999B09992",
-14344 => x"C0C0BFF999B09999",
-14343 => x"C0C0BFF999B099B0",
-14342 => x"C0C0BFF999B099A4",
-14341 => x"C0C0BFF999B099F9",
-14340 => x"C0C0BFF999B099C0",
-14339 => x"C0C0BFF999B0B090",
-14338 => x"C0C0BFF999B0B080",
-14337 => x"C0C0BFF999B0B0F8",
-14336 => x"C0C0BFF999B0B082",
-14335 => x"C0C0BFF999B0B092",
-14334 => x"C0C0BFF999B0B099",
-14333 => x"C0C0BFF999B0B0B0",
-14332 => x"C0C0BFF999B0B0A4",
-14331 => x"C0C0BFF999B0B0F9",
-14330 => x"C0C0BFF999B0B0C0",
-14329 => x"C0C0BFF999B0A490",
-14328 => x"C0C0BFF999B0A480",
-14327 => x"C0C0BFF999B0A4F8",
-14326 => x"C0C0BFF999B0A482",
-14325 => x"C0C0BFF999B0A492",
-14324 => x"C0C0BFF999B0A499",
-14323 => x"C0C0BFF999B0A4B0",
-14322 => x"C0C0BFF999B0A4A4",
-14321 => x"C0C0BFF999B0A4F9",
-14320 => x"C0C0BFF999B0A4C0",
-14319 => x"C0C0BFF999B0F990",
-14318 => x"C0C0BFF999B0F980",
-14317 => x"C0C0BFF999B0F9F8",
-14316 => x"C0C0BFF999B0F982",
-14315 => x"C0C0BFF999B0F992",
-14314 => x"C0C0BFF999B0F999",
-14313 => x"C0C0BFF999B0F9B0",
-14312 => x"C0C0BFF999B0F9A4",
-14311 => x"C0C0BFF999B0F9F9",
-14310 => x"C0C0BFF999B0F9C0",
-14309 => x"C0C0BFF999B0C090",
-14308 => x"C0C0BFF999B0C080",
-14307 => x"C0C0BFF999B0C0F8",
-14306 => x"C0C0BFF999B0C082",
-14305 => x"C0C0BFF999B0C092",
-14304 => x"C0C0BFF999B0C099",
-14303 => x"C0C0BFF999B0C0B0",
-14302 => x"C0C0BFF999B0C0A4",
-14301 => x"C0C0BFF999B0C0F9",
-14300 => x"C0C0BFF999B0C0C0",
-14299 => x"C0C0BFF999A49090",
-14298 => x"C0C0BFF999A49080",
-14297 => x"C0C0BFF999A490F8",
-14296 => x"C0C0BFF999A49082",
-14295 => x"C0C0BFF999A49092",
-14294 => x"C0C0BFF999A49099",
-14293 => x"C0C0BFF999A490B0",
-14292 => x"C0C0BFF999A490A4",
-14291 => x"C0C0BFF999A490F9",
-14290 => x"C0C0BFF999A490C0",
-14289 => x"C0C0BFF999A48090",
-14288 => x"C0C0BFF999A48080",
-14287 => x"C0C0BFF999A480F8",
-14286 => x"C0C0BFF999A48082",
-14285 => x"C0C0BFF999A48092",
-14284 => x"C0C0BFF999A48099",
-14283 => x"C0C0BFF999A480B0",
-14282 => x"C0C0BFF999A480A4",
-14281 => x"C0C0BFF999A480F9",
-14280 => x"C0C0BFF999A480C0",
-14279 => x"C0C0BFF999A4F890",
-14278 => x"C0C0BFF999A4F880",
-14277 => x"C0C0BFF999A4F8F8",
-14276 => x"C0C0BFF999A4F882",
-14275 => x"C0C0BFF999A4F892",
-14274 => x"C0C0BFF999A4F899",
-14273 => x"C0C0BFF999A4F8B0",
-14272 => x"C0C0BFF999A4F8A4",
-14271 => x"C0C0BFF999A4F8F9",
-14270 => x"C0C0BFF999A4F8C0",
-14269 => x"C0C0BFF999A48290",
-14268 => x"C0C0BFF999A48280",
-14267 => x"C0C0BFF999A482F8",
-14266 => x"C0C0BFF999A48282",
-14265 => x"C0C0BFF999A48292",
-14264 => x"C0C0BFF999A48299",
-14263 => x"C0C0BFF999A482B0",
-14262 => x"C0C0BFF999A482A4",
-14261 => x"C0C0BFF999A482F9",
-14260 => x"C0C0BFF999A482C0",
-14259 => x"C0C0BFF999A49290",
-14258 => x"C0C0BFF999A49280",
-14257 => x"C0C0BFF999A492F8",
-14256 => x"C0C0BFF999A49282",
-14255 => x"C0C0BFF999A49292",
-14254 => x"C0C0BFF999A49299",
-14253 => x"C0C0BFF999A492B0",
-14252 => x"C0C0BFF999A492A4",
-14251 => x"C0C0BFF999A492F9",
-14250 => x"C0C0BFF999A492C0",
-14249 => x"C0C0BFF999A49990",
-14248 => x"C0C0BFF999A49980",
-14247 => x"C0C0BFF999A499F8",
-14246 => x"C0C0BFF999A49982",
-14245 => x"C0C0BFF999A49992",
-14244 => x"C0C0BFF999A49999",
-14243 => x"C0C0BFF999A499B0",
-14242 => x"C0C0BFF999A499A4",
-14241 => x"C0C0BFF999A499F9",
-14240 => x"C0C0BFF999A499C0",
-14239 => x"C0C0BFF999A4B090",
-14238 => x"C0C0BFF999A4B080",
-14237 => x"C0C0BFF999A4B0F8",
-14236 => x"C0C0BFF999A4B082",
-14235 => x"C0C0BFF999A4B092",
-14234 => x"C0C0BFF999A4B099",
-14233 => x"C0C0BFF999A4B0B0",
-14232 => x"C0C0BFF999A4B0A4",
-14231 => x"C0C0BFF999A4B0F9",
-14230 => x"C0C0BFF999A4B0C0",
-14229 => x"C0C0BFF999A4A490",
-14228 => x"C0C0BFF999A4A480",
-14227 => x"C0C0BFF999A4A4F8",
-14226 => x"C0C0BFF999A4A482",
-14225 => x"C0C0BFF999A4A492",
-14224 => x"C0C0BFF999A4A499",
-14223 => x"C0C0BFF999A4A4B0",
-14222 => x"C0C0BFF999A4A4A4",
-14221 => x"C0C0BFF999A4A4F9",
-14220 => x"C0C0BFF999A4A4C0",
-14219 => x"C0C0BFF999A4F990",
-14218 => x"C0C0BFF999A4F980",
-14217 => x"C0C0BFF999A4F9F8",
-14216 => x"C0C0BFF999A4F982",
-14215 => x"C0C0BFF999A4F992",
-14214 => x"C0C0BFF999A4F999",
-14213 => x"C0C0BFF999A4F9B0",
-14212 => x"C0C0BFF999A4F9A4",
-14211 => x"C0C0BFF999A4F9F9",
-14210 => x"C0C0BFF999A4F9C0",
-14209 => x"C0C0BFF999A4C090",
-14208 => x"C0C0BFF999A4C080",
-14207 => x"C0C0BFF999A4C0F8",
-14206 => x"C0C0BFF999A4C082",
-14205 => x"C0C0BFF999A4C092",
-14204 => x"C0C0BFF999A4C099",
-14203 => x"C0C0BFF999A4C0B0",
-14202 => x"C0C0BFF999A4C0A4",
-14201 => x"C0C0BFF999A4C0F9",
-14200 => x"C0C0BFF999A4C0C0",
-14199 => x"C0C0BFF999F99090",
-14198 => x"C0C0BFF999F99080",
-14197 => x"C0C0BFF999F990F8",
-14196 => x"C0C0BFF999F99082",
-14195 => x"C0C0BFF999F99092",
-14194 => x"C0C0BFF999F99099",
-14193 => x"C0C0BFF999F990B0",
-14192 => x"C0C0BFF999F990A4",
-14191 => x"C0C0BFF999F990F9",
-14190 => x"C0C0BFF999F990C0",
-14189 => x"C0C0BFF999F98090",
-14188 => x"C0C0BFF999F98080",
-14187 => x"C0C0BFF999F980F8",
-14186 => x"C0C0BFF999F98082",
-14185 => x"C0C0BFF999F98092",
-14184 => x"C0C0BFF999F98099",
-14183 => x"C0C0BFF999F980B0",
-14182 => x"C0C0BFF999F980A4",
-14181 => x"C0C0BFF999F980F9",
-14180 => x"C0C0BFF999F980C0",
-14179 => x"C0C0BFF999F9F890",
-14178 => x"C0C0BFF999F9F880",
-14177 => x"C0C0BFF999F9F8F8",
-14176 => x"C0C0BFF999F9F882",
-14175 => x"C0C0BFF999F9F892",
-14174 => x"C0C0BFF999F9F899",
-14173 => x"C0C0BFF999F9F8B0",
-14172 => x"C0C0BFF999F9F8A4",
-14171 => x"C0C0BFF999F9F8F9",
-14170 => x"C0C0BFF999F9F8C0",
-14169 => x"C0C0BFF999F98290",
-14168 => x"C0C0BFF999F98280",
-14167 => x"C0C0BFF999F982F8",
-14166 => x"C0C0BFF999F98282",
-14165 => x"C0C0BFF999F98292",
-14164 => x"C0C0BFF999F98299",
-14163 => x"C0C0BFF999F982B0",
-14162 => x"C0C0BFF999F982A4",
-14161 => x"C0C0BFF999F982F9",
-14160 => x"C0C0BFF999F982C0",
-14159 => x"C0C0BFF999F99290",
-14158 => x"C0C0BFF999F99280",
-14157 => x"C0C0BFF999F992F8",
-14156 => x"C0C0BFF999F99282",
-14155 => x"C0C0BFF999F99292",
-14154 => x"C0C0BFF999F99299",
-14153 => x"C0C0BFF999F992B0",
-14152 => x"C0C0BFF999F992A4",
-14151 => x"C0C0BFF999F992F9",
-14150 => x"C0C0BFF999F992C0",
-14149 => x"C0C0BFF999F99990",
-14148 => x"C0C0BFF999F99980",
-14147 => x"C0C0BFF999F999F8",
-14146 => x"C0C0BFF999F99982",
-14145 => x"C0C0BFF999F99992",
-14144 => x"C0C0BFF999F99999",
-14143 => x"C0C0BFF999F999B0",
-14142 => x"C0C0BFF999F999A4",
-14141 => x"C0C0BFF999F999F9",
-14140 => x"C0C0BFF999F999C0",
-14139 => x"C0C0BFF999F9B090",
-14138 => x"C0C0BFF999F9B080",
-14137 => x"C0C0BFF999F9B0F8",
-14136 => x"C0C0BFF999F9B082",
-14135 => x"C0C0BFF999F9B092",
-14134 => x"C0C0BFF999F9B099",
-14133 => x"C0C0BFF999F9B0B0",
-14132 => x"C0C0BFF999F9B0A4",
-14131 => x"C0C0BFF999F9B0F9",
-14130 => x"C0C0BFF999F9B0C0",
-14129 => x"C0C0BFF999F9A490",
-14128 => x"C0C0BFF999F9A480",
-14127 => x"C0C0BFF999F9A4F8",
-14126 => x"C0C0BFF999F9A482",
-14125 => x"C0C0BFF999F9A492",
-14124 => x"C0C0BFF999F9A499",
-14123 => x"C0C0BFF999F9A4B0",
-14122 => x"C0C0BFF999F9A4A4",
-14121 => x"C0C0BFF999F9A4F9",
-14120 => x"C0C0BFF999F9A4C0",
-14119 => x"C0C0BFF999F9F990",
-14118 => x"C0C0BFF999F9F980",
-14117 => x"C0C0BFF999F9F9F8",
-14116 => x"C0C0BFF999F9F982",
-14115 => x"C0C0BFF999F9F992",
-14114 => x"C0C0BFF999F9F999",
-14113 => x"C0C0BFF999F9F9B0",
-14112 => x"C0C0BFF999F9F9A4",
-14111 => x"C0C0BFF999F9F9F9",
-14110 => x"C0C0BFF999F9F9C0",
-14109 => x"C0C0BFF999F9C090",
-14108 => x"C0C0BFF999F9C080",
-14107 => x"C0C0BFF999F9C0F8",
-14106 => x"C0C0BFF999F9C082",
-14105 => x"C0C0BFF999F9C092",
-14104 => x"C0C0BFF999F9C099",
-14103 => x"C0C0BFF999F9C0B0",
-14102 => x"C0C0BFF999F9C0A4",
-14101 => x"C0C0BFF999F9C0F9",
-14100 => x"C0C0BFF999F9C0C0",
-14099 => x"C0C0BFF999C09090",
-14098 => x"C0C0BFF999C09080",
-14097 => x"C0C0BFF999C090F8",
-14096 => x"C0C0BFF999C09082",
-14095 => x"C0C0BFF999C09092",
-14094 => x"C0C0BFF999C09099",
-14093 => x"C0C0BFF999C090B0",
-14092 => x"C0C0BFF999C090A4",
-14091 => x"C0C0BFF999C090F9",
-14090 => x"C0C0BFF999C090C0",
-14089 => x"C0C0BFF999C08090",
-14088 => x"C0C0BFF999C08080",
-14087 => x"C0C0BFF999C080F8",
-14086 => x"C0C0BFF999C08082",
-14085 => x"C0C0BFF999C08092",
-14084 => x"C0C0BFF999C08099",
-14083 => x"C0C0BFF999C080B0",
-14082 => x"C0C0BFF999C080A4",
-14081 => x"C0C0BFF999C080F9",
-14080 => x"C0C0BFF999C080C0",
-14079 => x"C0C0BFF999C0F890",
-14078 => x"C0C0BFF999C0F880",
-14077 => x"C0C0BFF999C0F8F8",
-14076 => x"C0C0BFF999C0F882",
-14075 => x"C0C0BFF999C0F892",
-14074 => x"C0C0BFF999C0F899",
-14073 => x"C0C0BFF999C0F8B0",
-14072 => x"C0C0BFF999C0F8A4",
-14071 => x"C0C0BFF999C0F8F9",
-14070 => x"C0C0BFF999C0F8C0",
-14069 => x"C0C0BFF999C08290",
-14068 => x"C0C0BFF999C08280",
-14067 => x"C0C0BFF999C082F8",
-14066 => x"C0C0BFF999C08282",
-14065 => x"C0C0BFF999C08292",
-14064 => x"C0C0BFF999C08299",
-14063 => x"C0C0BFF999C082B0",
-14062 => x"C0C0BFF999C082A4",
-14061 => x"C0C0BFF999C082F9",
-14060 => x"C0C0BFF999C082C0",
-14059 => x"C0C0BFF999C09290",
-14058 => x"C0C0BFF999C09280",
-14057 => x"C0C0BFF999C092F8",
-14056 => x"C0C0BFF999C09282",
-14055 => x"C0C0BFF999C09292",
-14054 => x"C0C0BFF999C09299",
-14053 => x"C0C0BFF999C092B0",
-14052 => x"C0C0BFF999C092A4",
-14051 => x"C0C0BFF999C092F9",
-14050 => x"C0C0BFF999C092C0",
-14049 => x"C0C0BFF999C09990",
-14048 => x"C0C0BFF999C09980",
-14047 => x"C0C0BFF999C099F8",
-14046 => x"C0C0BFF999C09982",
-14045 => x"C0C0BFF999C09992",
-14044 => x"C0C0BFF999C09999",
-14043 => x"C0C0BFF999C099B0",
-14042 => x"C0C0BFF999C099A4",
-14041 => x"C0C0BFF999C099F9",
-14040 => x"C0C0BFF999C099C0",
-14039 => x"C0C0BFF999C0B090",
-14038 => x"C0C0BFF999C0B080",
-14037 => x"C0C0BFF999C0B0F8",
-14036 => x"C0C0BFF999C0B082",
-14035 => x"C0C0BFF999C0B092",
-14034 => x"C0C0BFF999C0B099",
-14033 => x"C0C0BFF999C0B0B0",
-14032 => x"C0C0BFF999C0B0A4",
-14031 => x"C0C0BFF999C0B0F9",
-14030 => x"C0C0BFF999C0B0C0",
-14029 => x"C0C0BFF999C0A490",
-14028 => x"C0C0BFF999C0A480",
-14027 => x"C0C0BFF999C0A4F8",
-14026 => x"C0C0BFF999C0A482",
-14025 => x"C0C0BFF999C0A492",
-14024 => x"C0C0BFF999C0A499",
-14023 => x"C0C0BFF999C0A4B0",
-14022 => x"C0C0BFF999C0A4A4",
-14021 => x"C0C0BFF999C0A4F9",
-14020 => x"C0C0BFF999C0A4C0",
-14019 => x"C0C0BFF999C0F990",
-14018 => x"C0C0BFF999C0F980",
-14017 => x"C0C0BFF999C0F9F8",
-14016 => x"C0C0BFF999C0F982",
-14015 => x"C0C0BFF999C0F992",
-14014 => x"C0C0BFF999C0F999",
-14013 => x"C0C0BFF999C0F9B0",
-14012 => x"C0C0BFF999C0F9A4",
-14011 => x"C0C0BFF999C0F9F9",
-14010 => x"C0C0BFF999C0F9C0",
-14009 => x"C0C0BFF999C0C090",
-14008 => x"C0C0BFF999C0C080",
-14007 => x"C0C0BFF999C0C0F8",
-14006 => x"C0C0BFF999C0C082",
-14005 => x"C0C0BFF999C0C092",
-14004 => x"C0C0BFF999C0C099",
-14003 => x"C0C0BFF999C0C0B0",
-14002 => x"C0C0BFF999C0C0A4",
-14001 => x"C0C0BFF999C0C0F9",
-14000 => x"C0C0BFF999C0C0C0",
-13999 => x"C0C0BFF9B0909090",
-13998 => x"C0C0BFF9B0909080",
-13997 => x"C0C0BFF9B09090F8",
-13996 => x"C0C0BFF9B0909082",
-13995 => x"C0C0BFF9B0909092",
-13994 => x"C0C0BFF9B0909099",
-13993 => x"C0C0BFF9B09090B0",
-13992 => x"C0C0BFF9B09090A4",
-13991 => x"C0C0BFF9B09090F9",
-13990 => x"C0C0BFF9B09090C0",
-13989 => x"C0C0BFF9B0908090",
-13988 => x"C0C0BFF9B0908080",
-13987 => x"C0C0BFF9B09080F8",
-13986 => x"C0C0BFF9B0908082",
-13985 => x"C0C0BFF9B0908092",
-13984 => x"C0C0BFF9B0908099",
-13983 => x"C0C0BFF9B09080B0",
-13982 => x"C0C0BFF9B09080A4",
-13981 => x"C0C0BFF9B09080F9",
-13980 => x"C0C0BFF9B09080C0",
-13979 => x"C0C0BFF9B090F890",
-13978 => x"C0C0BFF9B090F880",
-13977 => x"C0C0BFF9B090F8F8",
-13976 => x"C0C0BFF9B090F882",
-13975 => x"C0C0BFF9B090F892",
-13974 => x"C0C0BFF9B090F899",
-13973 => x"C0C0BFF9B090F8B0",
-13972 => x"C0C0BFF9B090F8A4",
-13971 => x"C0C0BFF9B090F8F9",
-13970 => x"C0C0BFF9B090F8C0",
-13969 => x"C0C0BFF9B0908290",
-13968 => x"C0C0BFF9B0908280",
-13967 => x"C0C0BFF9B09082F8",
-13966 => x"C0C0BFF9B0908282",
-13965 => x"C0C0BFF9B0908292",
-13964 => x"C0C0BFF9B0908299",
-13963 => x"C0C0BFF9B09082B0",
-13962 => x"C0C0BFF9B09082A4",
-13961 => x"C0C0BFF9B09082F9",
-13960 => x"C0C0BFF9B09082C0",
-13959 => x"C0C0BFF9B0909290",
-13958 => x"C0C0BFF9B0909280",
-13957 => x"C0C0BFF9B09092F8",
-13956 => x"C0C0BFF9B0909282",
-13955 => x"C0C0BFF9B0909292",
-13954 => x"C0C0BFF9B0909299",
-13953 => x"C0C0BFF9B09092B0",
-13952 => x"C0C0BFF9B09092A4",
-13951 => x"C0C0BFF9B09092F9",
-13950 => x"C0C0BFF9B09092C0",
-13949 => x"C0C0BFF9B0909990",
-13948 => x"C0C0BFF9B0909980",
-13947 => x"C0C0BFF9B09099F8",
-13946 => x"C0C0BFF9B0909982",
-13945 => x"C0C0BFF9B0909992",
-13944 => x"C0C0BFF9B0909999",
-13943 => x"C0C0BFF9B09099B0",
-13942 => x"C0C0BFF9B09099A4",
-13941 => x"C0C0BFF9B09099F9",
-13940 => x"C0C0BFF9B09099C0",
-13939 => x"C0C0BFF9B090B090",
-13938 => x"C0C0BFF9B090B080",
-13937 => x"C0C0BFF9B090B0F8",
-13936 => x"C0C0BFF9B090B082",
-13935 => x"C0C0BFF9B090B092",
-13934 => x"C0C0BFF9B090B099",
-13933 => x"C0C0BFF9B090B0B0",
-13932 => x"C0C0BFF9B090B0A4",
-13931 => x"C0C0BFF9B090B0F9",
-13930 => x"C0C0BFF9B090B0C0",
-13929 => x"C0C0BFF9B090A490",
-13928 => x"C0C0BFF9B090A480",
-13927 => x"C0C0BFF9B090A4F8",
-13926 => x"C0C0BFF9B090A482",
-13925 => x"C0C0BFF9B090A492",
-13924 => x"C0C0BFF9B090A499",
-13923 => x"C0C0BFF9B090A4B0",
-13922 => x"C0C0BFF9B090A4A4",
-13921 => x"C0C0BFF9B090A4F9",
-13920 => x"C0C0BFF9B090A4C0",
-13919 => x"C0C0BFF9B090F990",
-13918 => x"C0C0BFF9B090F980",
-13917 => x"C0C0BFF9B090F9F8",
-13916 => x"C0C0BFF9B090F982",
-13915 => x"C0C0BFF9B090F992",
-13914 => x"C0C0BFF9B090F999",
-13913 => x"C0C0BFF9B090F9B0",
-13912 => x"C0C0BFF9B090F9A4",
-13911 => x"C0C0BFF9B090F9F9",
-13910 => x"C0C0BFF9B090F9C0",
-13909 => x"C0C0BFF9B090C090",
-13908 => x"C0C0BFF9B090C080",
-13907 => x"C0C0BFF9B090C0F8",
-13906 => x"C0C0BFF9B090C082",
-13905 => x"C0C0BFF9B090C092",
-13904 => x"C0C0BFF9B090C099",
-13903 => x"C0C0BFF9B090C0B0",
-13902 => x"C0C0BFF9B090C0A4",
-13901 => x"C0C0BFF9B090C0F9",
-13900 => x"C0C0BFF9B090C0C0",
-13899 => x"C0C0BFF9B0809090",
-13898 => x"C0C0BFF9B0809080",
-13897 => x"C0C0BFF9B08090F8",
-13896 => x"C0C0BFF9B0809082",
-13895 => x"C0C0BFF9B0809092",
-13894 => x"C0C0BFF9B0809099",
-13893 => x"C0C0BFF9B08090B0",
-13892 => x"C0C0BFF9B08090A4",
-13891 => x"C0C0BFF9B08090F9",
-13890 => x"C0C0BFF9B08090C0",
-13889 => x"C0C0BFF9B0808090",
-13888 => x"C0C0BFF9B0808080",
-13887 => x"C0C0BFF9B08080F8",
-13886 => x"C0C0BFF9B0808082",
-13885 => x"C0C0BFF9B0808092",
-13884 => x"C0C0BFF9B0808099",
-13883 => x"C0C0BFF9B08080B0",
-13882 => x"C0C0BFF9B08080A4",
-13881 => x"C0C0BFF9B08080F9",
-13880 => x"C0C0BFF9B08080C0",
-13879 => x"C0C0BFF9B080F890",
-13878 => x"C0C0BFF9B080F880",
-13877 => x"C0C0BFF9B080F8F8",
-13876 => x"C0C0BFF9B080F882",
-13875 => x"C0C0BFF9B080F892",
-13874 => x"C0C0BFF9B080F899",
-13873 => x"C0C0BFF9B080F8B0",
-13872 => x"C0C0BFF9B080F8A4",
-13871 => x"C0C0BFF9B080F8F9",
-13870 => x"C0C0BFF9B080F8C0",
-13869 => x"C0C0BFF9B0808290",
-13868 => x"C0C0BFF9B0808280",
-13867 => x"C0C0BFF9B08082F8",
-13866 => x"C0C0BFF9B0808282",
-13865 => x"C0C0BFF9B0808292",
-13864 => x"C0C0BFF9B0808299",
-13863 => x"C0C0BFF9B08082B0",
-13862 => x"C0C0BFF9B08082A4",
-13861 => x"C0C0BFF9B08082F9",
-13860 => x"C0C0BFF9B08082C0",
-13859 => x"C0C0BFF9B0809290",
-13858 => x"C0C0BFF9B0809280",
-13857 => x"C0C0BFF9B08092F8",
-13856 => x"C0C0BFF9B0809282",
-13855 => x"C0C0BFF9B0809292",
-13854 => x"C0C0BFF9B0809299",
-13853 => x"C0C0BFF9B08092B0",
-13852 => x"C0C0BFF9B08092A4",
-13851 => x"C0C0BFF9B08092F9",
-13850 => x"C0C0BFF9B08092C0",
-13849 => x"C0C0BFF9B0809990",
-13848 => x"C0C0BFF9B0809980",
-13847 => x"C0C0BFF9B08099F8",
-13846 => x"C0C0BFF9B0809982",
-13845 => x"C0C0BFF9B0809992",
-13844 => x"C0C0BFF9B0809999",
-13843 => x"C0C0BFF9B08099B0",
-13842 => x"C0C0BFF9B08099A4",
-13841 => x"C0C0BFF9B08099F9",
-13840 => x"C0C0BFF9B08099C0",
-13839 => x"C0C0BFF9B080B090",
-13838 => x"C0C0BFF9B080B080",
-13837 => x"C0C0BFF9B080B0F8",
-13836 => x"C0C0BFF9B080B082",
-13835 => x"C0C0BFF9B080B092",
-13834 => x"C0C0BFF9B080B099",
-13833 => x"C0C0BFF9B080B0B0",
-13832 => x"C0C0BFF9B080B0A4",
-13831 => x"C0C0BFF9B080B0F9",
-13830 => x"C0C0BFF9B080B0C0",
-13829 => x"C0C0BFF9B080A490",
-13828 => x"C0C0BFF9B080A480",
-13827 => x"C0C0BFF9B080A4F8",
-13826 => x"C0C0BFF9B080A482",
-13825 => x"C0C0BFF9B080A492",
-13824 => x"C0C0BFF9B080A499",
-13823 => x"C0C0BFF9B080A4B0",
-13822 => x"C0C0BFF9B080A4A4",
-13821 => x"C0C0BFF9B080A4F9",
-13820 => x"C0C0BFF9B080A4C0",
-13819 => x"C0C0BFF9B080F990",
-13818 => x"C0C0BFF9B080F980",
-13817 => x"C0C0BFF9B080F9F8",
-13816 => x"C0C0BFF9B080F982",
-13815 => x"C0C0BFF9B080F992",
-13814 => x"C0C0BFF9B080F999",
-13813 => x"C0C0BFF9B080F9B0",
-13812 => x"C0C0BFF9B080F9A4",
-13811 => x"C0C0BFF9B080F9F9",
-13810 => x"C0C0BFF9B080F9C0",
-13809 => x"C0C0BFF9B080C090",
-13808 => x"C0C0BFF9B080C080",
-13807 => x"C0C0BFF9B080C0F8",
-13806 => x"C0C0BFF9B080C082",
-13805 => x"C0C0BFF9B080C092",
-13804 => x"C0C0BFF9B080C099",
-13803 => x"C0C0BFF9B080C0B0",
-13802 => x"C0C0BFF9B080C0A4",
-13801 => x"C0C0BFF9B080C0F9",
-13800 => x"C0C0BFF9B080C0C0",
-13799 => x"C0C0BFF9B0F89090",
-13798 => x"C0C0BFF9B0F89080",
-13797 => x"C0C0BFF9B0F890F8",
-13796 => x"C0C0BFF9B0F89082",
-13795 => x"C0C0BFF9B0F89092",
-13794 => x"C0C0BFF9B0F89099",
-13793 => x"C0C0BFF9B0F890B0",
-13792 => x"C0C0BFF9B0F890A4",
-13791 => x"C0C0BFF9B0F890F9",
-13790 => x"C0C0BFF9B0F890C0",
-13789 => x"C0C0BFF9B0F88090",
-13788 => x"C0C0BFF9B0F88080",
-13787 => x"C0C0BFF9B0F880F8",
-13786 => x"C0C0BFF9B0F88082",
-13785 => x"C0C0BFF9B0F88092",
-13784 => x"C0C0BFF9B0F88099",
-13783 => x"C0C0BFF9B0F880B0",
-13782 => x"C0C0BFF9B0F880A4",
-13781 => x"C0C0BFF9B0F880F9",
-13780 => x"C0C0BFF9B0F880C0",
-13779 => x"C0C0BFF9B0F8F890",
-13778 => x"C0C0BFF9B0F8F880",
-13777 => x"C0C0BFF9B0F8F8F8",
-13776 => x"C0C0BFF9B0F8F882",
-13775 => x"C0C0BFF9B0F8F892",
-13774 => x"C0C0BFF9B0F8F899",
-13773 => x"C0C0BFF9B0F8F8B0",
-13772 => x"C0C0BFF9B0F8F8A4",
-13771 => x"C0C0BFF9B0F8F8F9",
-13770 => x"C0C0BFF9B0F8F8C0",
-13769 => x"C0C0BFF9B0F88290",
-13768 => x"C0C0BFF9B0F88280",
-13767 => x"C0C0BFF9B0F882F8",
-13766 => x"C0C0BFF9B0F88282",
-13765 => x"C0C0BFF9B0F88292",
-13764 => x"C0C0BFF9B0F88299",
-13763 => x"C0C0BFF9B0F882B0",
-13762 => x"C0C0BFF9B0F882A4",
-13761 => x"C0C0BFF9B0F882F9",
-13760 => x"C0C0BFF9B0F882C0",
-13759 => x"C0C0BFF9B0F89290",
-13758 => x"C0C0BFF9B0F89280",
-13757 => x"C0C0BFF9B0F892F8",
-13756 => x"C0C0BFF9B0F89282",
-13755 => x"C0C0BFF9B0F89292",
-13754 => x"C0C0BFF9B0F89299",
-13753 => x"C0C0BFF9B0F892B0",
-13752 => x"C0C0BFF9B0F892A4",
-13751 => x"C0C0BFF9B0F892F9",
-13750 => x"C0C0BFF9B0F892C0",
-13749 => x"C0C0BFF9B0F89990",
-13748 => x"C0C0BFF9B0F89980",
-13747 => x"C0C0BFF9B0F899F8",
-13746 => x"C0C0BFF9B0F89982",
-13745 => x"C0C0BFF9B0F89992",
-13744 => x"C0C0BFF9B0F89999",
-13743 => x"C0C0BFF9B0F899B0",
-13742 => x"C0C0BFF9B0F899A4",
-13741 => x"C0C0BFF9B0F899F9",
-13740 => x"C0C0BFF9B0F899C0",
-13739 => x"C0C0BFF9B0F8B090",
-13738 => x"C0C0BFF9B0F8B080",
-13737 => x"C0C0BFF9B0F8B0F8",
-13736 => x"C0C0BFF9B0F8B082",
-13735 => x"C0C0BFF9B0F8B092",
-13734 => x"C0C0BFF9B0F8B099",
-13733 => x"C0C0BFF9B0F8B0B0",
-13732 => x"C0C0BFF9B0F8B0A4",
-13731 => x"C0C0BFF9B0F8B0F9",
-13730 => x"C0C0BFF9B0F8B0C0",
-13729 => x"C0C0BFF9B0F8A490",
-13728 => x"C0C0BFF9B0F8A480",
-13727 => x"C0C0BFF9B0F8A4F8",
-13726 => x"C0C0BFF9B0F8A482",
-13725 => x"C0C0BFF9B0F8A492",
-13724 => x"C0C0BFF9B0F8A499",
-13723 => x"C0C0BFF9B0F8A4B0",
-13722 => x"C0C0BFF9B0F8A4A4",
-13721 => x"C0C0BFF9B0F8A4F9",
-13720 => x"C0C0BFF9B0F8A4C0",
-13719 => x"C0C0BFF9B0F8F990",
-13718 => x"C0C0BFF9B0F8F980",
-13717 => x"C0C0BFF9B0F8F9F8",
-13716 => x"C0C0BFF9B0F8F982",
-13715 => x"C0C0BFF9B0F8F992",
-13714 => x"C0C0BFF9B0F8F999",
-13713 => x"C0C0BFF9B0F8F9B0",
-13712 => x"C0C0BFF9B0F8F9A4",
-13711 => x"C0C0BFF9B0F8F9F9",
-13710 => x"C0C0BFF9B0F8F9C0",
-13709 => x"C0C0BFF9B0F8C090",
-13708 => x"C0C0BFF9B0F8C080",
-13707 => x"C0C0BFF9B0F8C0F8",
-13706 => x"C0C0BFF9B0F8C082",
-13705 => x"C0C0BFF9B0F8C092",
-13704 => x"C0C0BFF9B0F8C099",
-13703 => x"C0C0BFF9B0F8C0B0",
-13702 => x"C0C0BFF9B0F8C0A4",
-13701 => x"C0C0BFF9B0F8C0F9",
-13700 => x"C0C0BFF9B0F8C0C0",
-13699 => x"C0C0BFF9B0829090",
-13698 => x"C0C0BFF9B0829080",
-13697 => x"C0C0BFF9B08290F8",
-13696 => x"C0C0BFF9B0829082",
-13695 => x"C0C0BFF9B0829092",
-13694 => x"C0C0BFF9B0829099",
-13693 => x"C0C0BFF9B08290B0",
-13692 => x"C0C0BFF9B08290A4",
-13691 => x"C0C0BFF9B08290F9",
-13690 => x"C0C0BFF9B08290C0",
-13689 => x"C0C0BFF9B0828090",
-13688 => x"C0C0BFF9B0828080",
-13687 => x"C0C0BFF9B08280F8",
-13686 => x"C0C0BFF9B0828082",
-13685 => x"C0C0BFF9B0828092",
-13684 => x"C0C0BFF9B0828099",
-13683 => x"C0C0BFF9B08280B0",
-13682 => x"C0C0BFF9B08280A4",
-13681 => x"C0C0BFF9B08280F9",
-13680 => x"C0C0BFF9B08280C0",
-13679 => x"C0C0BFF9B082F890",
-13678 => x"C0C0BFF9B082F880",
-13677 => x"C0C0BFF9B082F8F8",
-13676 => x"C0C0BFF9B082F882",
-13675 => x"C0C0BFF9B082F892",
-13674 => x"C0C0BFF9B082F899",
-13673 => x"C0C0BFF9B082F8B0",
-13672 => x"C0C0BFF9B082F8A4",
-13671 => x"C0C0BFF9B082F8F9",
-13670 => x"C0C0BFF9B082F8C0",
-13669 => x"C0C0BFF9B0828290",
-13668 => x"C0C0BFF9B0828280",
-13667 => x"C0C0BFF9B08282F8",
-13666 => x"C0C0BFF9B0828282",
-13665 => x"C0C0BFF9B0828292",
-13664 => x"C0C0BFF9B0828299",
-13663 => x"C0C0BFF9B08282B0",
-13662 => x"C0C0BFF9B08282A4",
-13661 => x"C0C0BFF9B08282F9",
-13660 => x"C0C0BFF9B08282C0",
-13659 => x"C0C0BFF9B0829290",
-13658 => x"C0C0BFF9B0829280",
-13657 => x"C0C0BFF9B08292F8",
-13656 => x"C0C0BFF9B0829282",
-13655 => x"C0C0BFF9B0829292",
-13654 => x"C0C0BFF9B0829299",
-13653 => x"C0C0BFF9B08292B0",
-13652 => x"C0C0BFF9B08292A4",
-13651 => x"C0C0BFF9B08292F9",
-13650 => x"C0C0BFF9B08292C0",
-13649 => x"C0C0BFF9B0829990",
-13648 => x"C0C0BFF9B0829980",
-13647 => x"C0C0BFF9B08299F8",
-13646 => x"C0C0BFF9B0829982",
-13645 => x"C0C0BFF9B0829992",
-13644 => x"C0C0BFF9B0829999",
-13643 => x"C0C0BFF9B08299B0",
-13642 => x"C0C0BFF9B08299A4",
-13641 => x"C0C0BFF9B08299F9",
-13640 => x"C0C0BFF9B08299C0",
-13639 => x"C0C0BFF9B082B090",
-13638 => x"C0C0BFF9B082B080",
-13637 => x"C0C0BFF9B082B0F8",
-13636 => x"C0C0BFF9B082B082",
-13635 => x"C0C0BFF9B082B092",
-13634 => x"C0C0BFF9B082B099",
-13633 => x"C0C0BFF9B082B0B0",
-13632 => x"C0C0BFF9B082B0A4",
-13631 => x"C0C0BFF9B082B0F9",
-13630 => x"C0C0BFF9B082B0C0",
-13629 => x"C0C0BFF9B082A490",
-13628 => x"C0C0BFF9B082A480",
-13627 => x"C0C0BFF9B082A4F8",
-13626 => x"C0C0BFF9B082A482",
-13625 => x"C0C0BFF9B082A492",
-13624 => x"C0C0BFF9B082A499",
-13623 => x"C0C0BFF9B082A4B0",
-13622 => x"C0C0BFF9B082A4A4",
-13621 => x"C0C0BFF9B082A4F9",
-13620 => x"C0C0BFF9B082A4C0",
-13619 => x"C0C0BFF9B082F990",
-13618 => x"C0C0BFF9B082F980",
-13617 => x"C0C0BFF9B082F9F8",
-13616 => x"C0C0BFF9B082F982",
-13615 => x"C0C0BFF9B082F992",
-13614 => x"C0C0BFF9B082F999",
-13613 => x"C0C0BFF9B082F9B0",
-13612 => x"C0C0BFF9B082F9A4",
-13611 => x"C0C0BFF9B082F9F9",
-13610 => x"C0C0BFF9B082F9C0",
-13609 => x"C0C0BFF9B082C090",
-13608 => x"C0C0BFF9B082C080",
-13607 => x"C0C0BFF9B082C0F8",
-13606 => x"C0C0BFF9B082C082",
-13605 => x"C0C0BFF9B082C092",
-13604 => x"C0C0BFF9B082C099",
-13603 => x"C0C0BFF9B082C0B0",
-13602 => x"C0C0BFF9B082C0A4",
-13601 => x"C0C0BFF9B082C0F9",
-13600 => x"C0C0BFF9B082C0C0",
-13599 => x"C0C0BFF9B0929090",
-13598 => x"C0C0BFF9B0929080",
-13597 => x"C0C0BFF9B09290F8",
-13596 => x"C0C0BFF9B0929082",
-13595 => x"C0C0BFF9B0929092",
-13594 => x"C0C0BFF9B0929099",
-13593 => x"C0C0BFF9B09290B0",
-13592 => x"C0C0BFF9B09290A4",
-13591 => x"C0C0BFF9B09290F9",
-13590 => x"C0C0BFF9B09290C0",
-13589 => x"C0C0BFF9B0928090",
-13588 => x"C0C0BFF9B0928080",
-13587 => x"C0C0BFF9B09280F8",
-13586 => x"C0C0BFF9B0928082",
-13585 => x"C0C0BFF9B0928092",
-13584 => x"C0C0BFF9B0928099",
-13583 => x"C0C0BFF9B09280B0",
-13582 => x"C0C0BFF9B09280A4",
-13581 => x"C0C0BFF9B09280F9",
-13580 => x"C0C0BFF9B09280C0",
-13579 => x"C0C0BFF9B092F890",
-13578 => x"C0C0BFF9B092F880",
-13577 => x"C0C0BFF9B092F8F8",
-13576 => x"C0C0BFF9B092F882",
-13575 => x"C0C0BFF9B092F892",
-13574 => x"C0C0BFF9B092F899",
-13573 => x"C0C0BFF9B092F8B0",
-13572 => x"C0C0BFF9B092F8A4",
-13571 => x"C0C0BFF9B092F8F9",
-13570 => x"C0C0BFF9B092F8C0",
-13569 => x"C0C0BFF9B0928290",
-13568 => x"C0C0BFF9B0928280",
-13567 => x"C0C0BFF9B09282F8",
-13566 => x"C0C0BFF9B0928282",
-13565 => x"C0C0BFF9B0928292",
-13564 => x"C0C0BFF9B0928299",
-13563 => x"C0C0BFF9B09282B0",
-13562 => x"C0C0BFF9B09282A4",
-13561 => x"C0C0BFF9B09282F9",
-13560 => x"C0C0BFF9B09282C0",
-13559 => x"C0C0BFF9B0929290",
-13558 => x"C0C0BFF9B0929280",
-13557 => x"C0C0BFF9B09292F8",
-13556 => x"C0C0BFF9B0929282",
-13555 => x"C0C0BFF9B0929292",
-13554 => x"C0C0BFF9B0929299",
-13553 => x"C0C0BFF9B09292B0",
-13552 => x"C0C0BFF9B09292A4",
-13551 => x"C0C0BFF9B09292F9",
-13550 => x"C0C0BFF9B09292C0",
-13549 => x"C0C0BFF9B0929990",
-13548 => x"C0C0BFF9B0929980",
-13547 => x"C0C0BFF9B09299F8",
-13546 => x"C0C0BFF9B0929982",
-13545 => x"C0C0BFF9B0929992",
-13544 => x"C0C0BFF9B0929999",
-13543 => x"C0C0BFF9B09299B0",
-13542 => x"C0C0BFF9B09299A4",
-13541 => x"C0C0BFF9B09299F9",
-13540 => x"C0C0BFF9B09299C0",
-13539 => x"C0C0BFF9B092B090",
-13538 => x"C0C0BFF9B092B080",
-13537 => x"C0C0BFF9B092B0F8",
-13536 => x"C0C0BFF9B092B082",
-13535 => x"C0C0BFF9B092B092",
-13534 => x"C0C0BFF9B092B099",
-13533 => x"C0C0BFF9B092B0B0",
-13532 => x"C0C0BFF9B092B0A4",
-13531 => x"C0C0BFF9B092B0F9",
-13530 => x"C0C0BFF9B092B0C0",
-13529 => x"C0C0BFF9B092A490",
-13528 => x"C0C0BFF9B092A480",
-13527 => x"C0C0BFF9B092A4F8",
-13526 => x"C0C0BFF9B092A482",
-13525 => x"C0C0BFF9B092A492",
-13524 => x"C0C0BFF9B092A499",
-13523 => x"C0C0BFF9B092A4B0",
-13522 => x"C0C0BFF9B092A4A4",
-13521 => x"C0C0BFF9B092A4F9",
-13520 => x"C0C0BFF9B092A4C0",
-13519 => x"C0C0BFF9B092F990",
-13518 => x"C0C0BFF9B092F980",
-13517 => x"C0C0BFF9B092F9F8",
-13516 => x"C0C0BFF9B092F982",
-13515 => x"C0C0BFF9B092F992",
-13514 => x"C0C0BFF9B092F999",
-13513 => x"C0C0BFF9B092F9B0",
-13512 => x"C0C0BFF9B092F9A4",
-13511 => x"C0C0BFF9B092F9F9",
-13510 => x"C0C0BFF9B092F9C0",
-13509 => x"C0C0BFF9B092C090",
-13508 => x"C0C0BFF9B092C080",
-13507 => x"C0C0BFF9B092C0F8",
-13506 => x"C0C0BFF9B092C082",
-13505 => x"C0C0BFF9B092C092",
-13504 => x"C0C0BFF9B092C099",
-13503 => x"C0C0BFF9B092C0B0",
-13502 => x"C0C0BFF9B092C0A4",
-13501 => x"C0C0BFF9B092C0F9",
-13500 => x"C0C0BFF9B092C0C0",
-13499 => x"C0C0BFF9B0999090",
-13498 => x"C0C0BFF9B0999080",
-13497 => x"C0C0BFF9B09990F8",
-13496 => x"C0C0BFF9B0999082",
-13495 => x"C0C0BFF9B0999092",
-13494 => x"C0C0BFF9B0999099",
-13493 => x"C0C0BFF9B09990B0",
-13492 => x"C0C0BFF9B09990A4",
-13491 => x"C0C0BFF9B09990F9",
-13490 => x"C0C0BFF9B09990C0",
-13489 => x"C0C0BFF9B0998090",
-13488 => x"C0C0BFF9B0998080",
-13487 => x"C0C0BFF9B09980F8",
-13486 => x"C0C0BFF9B0998082",
-13485 => x"C0C0BFF9B0998092",
-13484 => x"C0C0BFF9B0998099",
-13483 => x"C0C0BFF9B09980B0",
-13482 => x"C0C0BFF9B09980A4",
-13481 => x"C0C0BFF9B09980F9",
-13480 => x"C0C0BFF9B09980C0",
-13479 => x"C0C0BFF9B099F890",
-13478 => x"C0C0BFF9B099F880",
-13477 => x"C0C0BFF9B099F8F8",
-13476 => x"C0C0BFF9B099F882",
-13475 => x"C0C0BFF9B099F892",
-13474 => x"C0C0BFF9B099F899",
-13473 => x"C0C0BFF9B099F8B0",
-13472 => x"C0C0BFF9B099F8A4",
-13471 => x"C0C0BFF9B099F8F9",
-13470 => x"C0C0BFF9B099F8C0",
-13469 => x"C0C0BFF9B0998290",
-13468 => x"C0C0BFF9B0998280",
-13467 => x"C0C0BFF9B09982F8",
-13466 => x"C0C0BFF9B0998282",
-13465 => x"C0C0BFF9B0998292",
-13464 => x"C0C0BFF9B0998299",
-13463 => x"C0C0BFF9B09982B0",
-13462 => x"C0C0BFF9B09982A4",
-13461 => x"C0C0BFF9B09982F9",
-13460 => x"C0C0BFF9B09982C0",
-13459 => x"C0C0BFF9B0999290",
-13458 => x"C0C0BFF9B0999280",
-13457 => x"C0C0BFF9B09992F8",
-13456 => x"C0C0BFF9B0999282",
-13455 => x"C0C0BFF9B0999292",
-13454 => x"C0C0BFF9B0999299",
-13453 => x"C0C0BFF9B09992B0",
-13452 => x"C0C0BFF9B09992A4",
-13451 => x"C0C0BFF9B09992F9",
-13450 => x"C0C0BFF9B09992C0",
-13449 => x"C0C0BFF9B0999990",
-13448 => x"C0C0BFF9B0999980",
-13447 => x"C0C0BFF9B09999F8",
-13446 => x"C0C0BFF9B0999982",
-13445 => x"C0C0BFF9B0999992",
-13444 => x"C0C0BFF9B0999999",
-13443 => x"C0C0BFF9B09999B0",
-13442 => x"C0C0BFF9B09999A4",
-13441 => x"C0C0BFF9B09999F9",
-13440 => x"C0C0BFF9B09999C0",
-13439 => x"C0C0BFF9B099B090",
-13438 => x"C0C0BFF9B099B080",
-13437 => x"C0C0BFF9B099B0F8",
-13436 => x"C0C0BFF9B099B082",
-13435 => x"C0C0BFF9B099B092",
-13434 => x"C0C0BFF9B099B099",
-13433 => x"C0C0BFF9B099B0B0",
-13432 => x"C0C0BFF9B099B0A4",
-13431 => x"C0C0BFF9B099B0F9",
-13430 => x"C0C0BFF9B099B0C0",
-13429 => x"C0C0BFF9B099A490",
-13428 => x"C0C0BFF9B099A480",
-13427 => x"C0C0BFF9B099A4F8",
-13426 => x"C0C0BFF9B099A482",
-13425 => x"C0C0BFF9B099A492",
-13424 => x"C0C0BFF9B099A499",
-13423 => x"C0C0BFF9B099A4B0",
-13422 => x"C0C0BFF9B099A4A4",
-13421 => x"C0C0BFF9B099A4F9",
-13420 => x"C0C0BFF9B099A4C0",
-13419 => x"C0C0BFF9B099F990",
-13418 => x"C0C0BFF9B099F980",
-13417 => x"C0C0BFF9B099F9F8",
-13416 => x"C0C0BFF9B099F982",
-13415 => x"C0C0BFF9B099F992",
-13414 => x"C0C0BFF9B099F999",
-13413 => x"C0C0BFF9B099F9B0",
-13412 => x"C0C0BFF9B099F9A4",
-13411 => x"C0C0BFF9B099F9F9",
-13410 => x"C0C0BFF9B099F9C0",
-13409 => x"C0C0BFF9B099C090",
-13408 => x"C0C0BFF9B099C080",
-13407 => x"C0C0BFF9B099C0F8",
-13406 => x"C0C0BFF9B099C082",
-13405 => x"C0C0BFF9B099C092",
-13404 => x"C0C0BFF9B099C099",
-13403 => x"C0C0BFF9B099C0B0",
-13402 => x"C0C0BFF9B099C0A4",
-13401 => x"C0C0BFF9B099C0F9",
-13400 => x"C0C0BFF9B099C0C0",
-13399 => x"C0C0BFF9B0B09090",
-13398 => x"C0C0BFF9B0B09080",
-13397 => x"C0C0BFF9B0B090F8",
-13396 => x"C0C0BFF9B0B09082",
-13395 => x"C0C0BFF9B0B09092",
-13394 => x"C0C0BFF9B0B09099",
-13393 => x"C0C0BFF9B0B090B0",
-13392 => x"C0C0BFF9B0B090A4",
-13391 => x"C0C0BFF9B0B090F9",
-13390 => x"C0C0BFF9B0B090C0",
-13389 => x"C0C0BFF9B0B08090",
-13388 => x"C0C0BFF9B0B08080",
-13387 => x"C0C0BFF9B0B080F8",
-13386 => x"C0C0BFF9B0B08082",
-13385 => x"C0C0BFF9B0B08092",
-13384 => x"C0C0BFF9B0B08099",
-13383 => x"C0C0BFF9B0B080B0",
-13382 => x"C0C0BFF9B0B080A4",
-13381 => x"C0C0BFF9B0B080F9",
-13380 => x"C0C0BFF9B0B080C0",
-13379 => x"C0C0BFF9B0B0F890",
-13378 => x"C0C0BFF9B0B0F880",
-13377 => x"C0C0BFF9B0B0F8F8",
-13376 => x"C0C0BFF9B0B0F882",
-13375 => x"C0C0BFF9B0B0F892",
-13374 => x"C0C0BFF9B0B0F899",
-13373 => x"C0C0BFF9B0B0F8B0",
-13372 => x"C0C0BFF9B0B0F8A4",
-13371 => x"C0C0BFF9B0B0F8F9",
-13370 => x"C0C0BFF9B0B0F8C0",
-13369 => x"C0C0BFF9B0B08290",
-13368 => x"C0C0BFF9B0B08280",
-13367 => x"C0C0BFF9B0B082F8",
-13366 => x"C0C0BFF9B0B08282",
-13365 => x"C0C0BFF9B0B08292",
-13364 => x"C0C0BFF9B0B08299",
-13363 => x"C0C0BFF9B0B082B0",
-13362 => x"C0C0BFF9B0B082A4",
-13361 => x"C0C0BFF9B0B082F9",
-13360 => x"C0C0BFF9B0B082C0",
-13359 => x"C0C0BFF9B0B09290",
-13358 => x"C0C0BFF9B0B09280",
-13357 => x"C0C0BFF9B0B092F8",
-13356 => x"C0C0BFF9B0B09282",
-13355 => x"C0C0BFF9B0B09292",
-13354 => x"C0C0BFF9B0B09299",
-13353 => x"C0C0BFF9B0B092B0",
-13352 => x"C0C0BFF9B0B092A4",
-13351 => x"C0C0BFF9B0B092F9",
-13350 => x"C0C0BFF9B0B092C0",
-13349 => x"C0C0BFF9B0B09990",
-13348 => x"C0C0BFF9B0B09980",
-13347 => x"C0C0BFF9B0B099F8",
-13346 => x"C0C0BFF9B0B09982",
-13345 => x"C0C0BFF9B0B09992",
-13344 => x"C0C0BFF9B0B09999",
-13343 => x"C0C0BFF9B0B099B0",
-13342 => x"C0C0BFF9B0B099A4",
-13341 => x"C0C0BFF9B0B099F9",
-13340 => x"C0C0BFF9B0B099C0",
-13339 => x"C0C0BFF9B0B0B090",
-13338 => x"C0C0BFF9B0B0B080",
-13337 => x"C0C0BFF9B0B0B0F8",
-13336 => x"C0C0BFF9B0B0B082",
-13335 => x"C0C0BFF9B0B0B092",
-13334 => x"C0C0BFF9B0B0B099",
-13333 => x"C0C0BFF9B0B0B0B0",
-13332 => x"C0C0BFF9B0B0B0A4",
-13331 => x"C0C0BFF9B0B0B0F9",
-13330 => x"C0C0BFF9B0B0B0C0",
-13329 => x"C0C0BFF9B0B0A490",
-13328 => x"C0C0BFF9B0B0A480",
-13327 => x"C0C0BFF9B0B0A4F8",
-13326 => x"C0C0BFF9B0B0A482",
-13325 => x"C0C0BFF9B0B0A492",
-13324 => x"C0C0BFF9B0B0A499",
-13323 => x"C0C0BFF9B0B0A4B0",
-13322 => x"C0C0BFF9B0B0A4A4",
-13321 => x"C0C0BFF9B0B0A4F9",
-13320 => x"C0C0BFF9B0B0A4C0",
-13319 => x"C0C0BFF9B0B0F990",
-13318 => x"C0C0BFF9B0B0F980",
-13317 => x"C0C0BFF9B0B0F9F8",
-13316 => x"C0C0BFF9B0B0F982",
-13315 => x"C0C0BFF9B0B0F992",
-13314 => x"C0C0BFF9B0B0F999",
-13313 => x"C0C0BFF9B0B0F9B0",
-13312 => x"C0C0BFF9B0B0F9A4",
-13311 => x"C0C0BFF9B0B0F9F9",
-13310 => x"C0C0BFF9B0B0F9C0",
-13309 => x"C0C0BFF9B0B0C090",
-13308 => x"C0C0BFF9B0B0C080",
-13307 => x"C0C0BFF9B0B0C0F8",
-13306 => x"C0C0BFF9B0B0C082",
-13305 => x"C0C0BFF9B0B0C092",
-13304 => x"C0C0BFF9B0B0C099",
-13303 => x"C0C0BFF9B0B0C0B0",
-13302 => x"C0C0BFF9B0B0C0A4",
-13301 => x"C0C0BFF9B0B0C0F9",
-13300 => x"C0C0BFF9B0B0C0C0",
-13299 => x"C0C0BFF9B0A49090",
-13298 => x"C0C0BFF9B0A49080",
-13297 => x"C0C0BFF9B0A490F8",
-13296 => x"C0C0BFF9B0A49082",
-13295 => x"C0C0BFF9B0A49092",
-13294 => x"C0C0BFF9B0A49099",
-13293 => x"C0C0BFF9B0A490B0",
-13292 => x"C0C0BFF9B0A490A4",
-13291 => x"C0C0BFF9B0A490F9",
-13290 => x"C0C0BFF9B0A490C0",
-13289 => x"C0C0BFF9B0A48090",
-13288 => x"C0C0BFF9B0A48080",
-13287 => x"C0C0BFF9B0A480F8",
-13286 => x"C0C0BFF9B0A48082",
-13285 => x"C0C0BFF9B0A48092",
-13284 => x"C0C0BFF9B0A48099",
-13283 => x"C0C0BFF9B0A480B0",
-13282 => x"C0C0BFF9B0A480A4",
-13281 => x"C0C0BFF9B0A480F9",
-13280 => x"C0C0BFF9B0A480C0",
-13279 => x"C0C0BFF9B0A4F890",
-13278 => x"C0C0BFF9B0A4F880",
-13277 => x"C0C0BFF9B0A4F8F8",
-13276 => x"C0C0BFF9B0A4F882",
-13275 => x"C0C0BFF9B0A4F892",
-13274 => x"C0C0BFF9B0A4F899",
-13273 => x"C0C0BFF9B0A4F8B0",
-13272 => x"C0C0BFF9B0A4F8A4",
-13271 => x"C0C0BFF9B0A4F8F9",
-13270 => x"C0C0BFF9B0A4F8C0",
-13269 => x"C0C0BFF9B0A48290",
-13268 => x"C0C0BFF9B0A48280",
-13267 => x"C0C0BFF9B0A482F8",
-13266 => x"C0C0BFF9B0A48282",
-13265 => x"C0C0BFF9B0A48292",
-13264 => x"C0C0BFF9B0A48299",
-13263 => x"C0C0BFF9B0A482B0",
-13262 => x"C0C0BFF9B0A482A4",
-13261 => x"C0C0BFF9B0A482F9",
-13260 => x"C0C0BFF9B0A482C0",
-13259 => x"C0C0BFF9B0A49290",
-13258 => x"C0C0BFF9B0A49280",
-13257 => x"C0C0BFF9B0A492F8",
-13256 => x"C0C0BFF9B0A49282",
-13255 => x"C0C0BFF9B0A49292",
-13254 => x"C0C0BFF9B0A49299",
-13253 => x"C0C0BFF9B0A492B0",
-13252 => x"C0C0BFF9B0A492A4",
-13251 => x"C0C0BFF9B0A492F9",
-13250 => x"C0C0BFF9B0A492C0",
-13249 => x"C0C0BFF9B0A49990",
-13248 => x"C0C0BFF9B0A49980",
-13247 => x"C0C0BFF9B0A499F8",
-13246 => x"C0C0BFF9B0A49982",
-13245 => x"C0C0BFF9B0A49992",
-13244 => x"C0C0BFF9B0A49999",
-13243 => x"C0C0BFF9B0A499B0",
-13242 => x"C0C0BFF9B0A499A4",
-13241 => x"C0C0BFF9B0A499F9",
-13240 => x"C0C0BFF9B0A499C0",
-13239 => x"C0C0BFF9B0A4B090",
-13238 => x"C0C0BFF9B0A4B080",
-13237 => x"C0C0BFF9B0A4B0F8",
-13236 => x"C0C0BFF9B0A4B082",
-13235 => x"C0C0BFF9B0A4B092",
-13234 => x"C0C0BFF9B0A4B099",
-13233 => x"C0C0BFF9B0A4B0B0",
-13232 => x"C0C0BFF9B0A4B0A4",
-13231 => x"C0C0BFF9B0A4B0F9",
-13230 => x"C0C0BFF9B0A4B0C0",
-13229 => x"C0C0BFF9B0A4A490",
-13228 => x"C0C0BFF9B0A4A480",
-13227 => x"C0C0BFF9B0A4A4F8",
-13226 => x"C0C0BFF9B0A4A482",
-13225 => x"C0C0BFF9B0A4A492",
-13224 => x"C0C0BFF9B0A4A499",
-13223 => x"C0C0BFF9B0A4A4B0",
-13222 => x"C0C0BFF9B0A4A4A4",
-13221 => x"C0C0BFF9B0A4A4F9",
-13220 => x"C0C0BFF9B0A4A4C0",
-13219 => x"C0C0BFF9B0A4F990",
-13218 => x"C0C0BFF9B0A4F980",
-13217 => x"C0C0BFF9B0A4F9F8",
-13216 => x"C0C0BFF9B0A4F982",
-13215 => x"C0C0BFF9B0A4F992",
-13214 => x"C0C0BFF9B0A4F999",
-13213 => x"C0C0BFF9B0A4F9B0",
-13212 => x"C0C0BFF9B0A4F9A4",
-13211 => x"C0C0BFF9B0A4F9F9",
-13210 => x"C0C0BFF9B0A4F9C0",
-13209 => x"C0C0BFF9B0A4C090",
-13208 => x"C0C0BFF9B0A4C080",
-13207 => x"C0C0BFF9B0A4C0F8",
-13206 => x"C0C0BFF9B0A4C082",
-13205 => x"C0C0BFF9B0A4C092",
-13204 => x"C0C0BFF9B0A4C099",
-13203 => x"C0C0BFF9B0A4C0B0",
-13202 => x"C0C0BFF9B0A4C0A4",
-13201 => x"C0C0BFF9B0A4C0F9",
-13200 => x"C0C0BFF9B0A4C0C0",
-13199 => x"C0C0BFF9B0F99090",
-13198 => x"C0C0BFF9B0F99080",
-13197 => x"C0C0BFF9B0F990F8",
-13196 => x"C0C0BFF9B0F99082",
-13195 => x"C0C0BFF9B0F99092",
-13194 => x"C0C0BFF9B0F99099",
-13193 => x"C0C0BFF9B0F990B0",
-13192 => x"C0C0BFF9B0F990A4",
-13191 => x"C0C0BFF9B0F990F9",
-13190 => x"C0C0BFF9B0F990C0",
-13189 => x"C0C0BFF9B0F98090",
-13188 => x"C0C0BFF9B0F98080",
-13187 => x"C0C0BFF9B0F980F8",
-13186 => x"C0C0BFF9B0F98082",
-13185 => x"C0C0BFF9B0F98092",
-13184 => x"C0C0BFF9B0F98099",
-13183 => x"C0C0BFF9B0F980B0",
-13182 => x"C0C0BFF9B0F980A4",
-13181 => x"C0C0BFF9B0F980F9",
-13180 => x"C0C0BFF9B0F980C0",
-13179 => x"C0C0BFF9B0F9F890",
-13178 => x"C0C0BFF9B0F9F880",
-13177 => x"C0C0BFF9B0F9F8F8",
-13176 => x"C0C0BFF9B0F9F882",
-13175 => x"C0C0BFF9B0F9F892",
-13174 => x"C0C0BFF9B0F9F899",
-13173 => x"C0C0BFF9B0F9F8B0",
-13172 => x"C0C0BFF9B0F9F8A4",
-13171 => x"C0C0BFF9B0F9F8F9",
-13170 => x"C0C0BFF9B0F9F8C0",
-13169 => x"C0C0BFF9B0F98290",
-13168 => x"C0C0BFF9B0F98280",
-13167 => x"C0C0BFF9B0F982F8",
-13166 => x"C0C0BFF9B0F98282",
-13165 => x"C0C0BFF9B0F98292",
-13164 => x"C0C0BFF9B0F98299",
-13163 => x"C0C0BFF9B0F982B0",
-13162 => x"C0C0BFF9B0F982A4",
-13161 => x"C0C0BFF9B0F982F9",
-13160 => x"C0C0BFF9B0F982C0",
-13159 => x"C0C0BFF9B0F99290",
-13158 => x"C0C0BFF9B0F99280",
-13157 => x"C0C0BFF9B0F992F8",
-13156 => x"C0C0BFF9B0F99282",
-13155 => x"C0C0BFF9B0F99292",
-13154 => x"C0C0BFF9B0F99299",
-13153 => x"C0C0BFF9B0F992B0",
-13152 => x"C0C0BFF9B0F992A4",
-13151 => x"C0C0BFF9B0F992F9",
-13150 => x"C0C0BFF9B0F992C0",
-13149 => x"C0C0BFF9B0F99990",
-13148 => x"C0C0BFF9B0F99980",
-13147 => x"C0C0BFF9B0F999F8",
-13146 => x"C0C0BFF9B0F99982",
-13145 => x"C0C0BFF9B0F99992",
-13144 => x"C0C0BFF9B0F99999",
-13143 => x"C0C0BFF9B0F999B0",
-13142 => x"C0C0BFF9B0F999A4",
-13141 => x"C0C0BFF9B0F999F9",
-13140 => x"C0C0BFF9B0F999C0",
-13139 => x"C0C0BFF9B0F9B090",
-13138 => x"C0C0BFF9B0F9B080",
-13137 => x"C0C0BFF9B0F9B0F8",
-13136 => x"C0C0BFF9B0F9B082",
-13135 => x"C0C0BFF9B0F9B092",
-13134 => x"C0C0BFF9B0F9B099",
-13133 => x"C0C0BFF9B0F9B0B0",
-13132 => x"C0C0BFF9B0F9B0A4",
-13131 => x"C0C0BFF9B0F9B0F9",
-13130 => x"C0C0BFF9B0F9B0C0",
-13129 => x"C0C0BFF9B0F9A490",
-13128 => x"C0C0BFF9B0F9A480",
-13127 => x"C0C0BFF9B0F9A4F8",
-13126 => x"C0C0BFF9B0F9A482",
-13125 => x"C0C0BFF9B0F9A492",
-13124 => x"C0C0BFF9B0F9A499",
-13123 => x"C0C0BFF9B0F9A4B0",
-13122 => x"C0C0BFF9B0F9A4A4",
-13121 => x"C0C0BFF9B0F9A4F9",
-13120 => x"C0C0BFF9B0F9A4C0",
-13119 => x"C0C0BFF9B0F9F990",
-13118 => x"C0C0BFF9B0F9F980",
-13117 => x"C0C0BFF9B0F9F9F8",
-13116 => x"C0C0BFF9B0F9F982",
-13115 => x"C0C0BFF9B0F9F992",
-13114 => x"C0C0BFF9B0F9F999",
-13113 => x"C0C0BFF9B0F9F9B0",
-13112 => x"C0C0BFF9B0F9F9A4",
-13111 => x"C0C0BFF9B0F9F9F9",
-13110 => x"C0C0BFF9B0F9F9C0",
-13109 => x"C0C0BFF9B0F9C090",
-13108 => x"C0C0BFF9B0F9C080",
-13107 => x"C0C0BFF9B0F9C0F8",
-13106 => x"C0C0BFF9B0F9C082",
-13105 => x"C0C0BFF9B0F9C092",
-13104 => x"C0C0BFF9B0F9C099",
-13103 => x"C0C0BFF9B0F9C0B0",
-13102 => x"C0C0BFF9B0F9C0A4",
-13101 => x"C0C0BFF9B0F9C0F9",
-13100 => x"C0C0BFF9B0F9C0C0",
-13099 => x"C0C0BFF9B0C09090",
-13098 => x"C0C0BFF9B0C09080",
-13097 => x"C0C0BFF9B0C090F8",
-13096 => x"C0C0BFF9B0C09082",
-13095 => x"C0C0BFF9B0C09092",
-13094 => x"C0C0BFF9B0C09099",
-13093 => x"C0C0BFF9B0C090B0",
-13092 => x"C0C0BFF9B0C090A4",
-13091 => x"C0C0BFF9B0C090F9",
-13090 => x"C0C0BFF9B0C090C0",
-13089 => x"C0C0BFF9B0C08090",
-13088 => x"C0C0BFF9B0C08080",
-13087 => x"C0C0BFF9B0C080F8",
-13086 => x"C0C0BFF9B0C08082",
-13085 => x"C0C0BFF9B0C08092",
-13084 => x"C0C0BFF9B0C08099",
-13083 => x"C0C0BFF9B0C080B0",
-13082 => x"C0C0BFF9B0C080A4",
-13081 => x"C0C0BFF9B0C080F9",
-13080 => x"C0C0BFF9B0C080C0",
-13079 => x"C0C0BFF9B0C0F890",
-13078 => x"C0C0BFF9B0C0F880",
-13077 => x"C0C0BFF9B0C0F8F8",
-13076 => x"C0C0BFF9B0C0F882",
-13075 => x"C0C0BFF9B0C0F892",
-13074 => x"C0C0BFF9B0C0F899",
-13073 => x"C0C0BFF9B0C0F8B0",
-13072 => x"C0C0BFF9B0C0F8A4",
-13071 => x"C0C0BFF9B0C0F8F9",
-13070 => x"C0C0BFF9B0C0F8C0",
-13069 => x"C0C0BFF9B0C08290",
-13068 => x"C0C0BFF9B0C08280",
-13067 => x"C0C0BFF9B0C082F8",
-13066 => x"C0C0BFF9B0C08282",
-13065 => x"C0C0BFF9B0C08292",
-13064 => x"C0C0BFF9B0C08299",
-13063 => x"C0C0BFF9B0C082B0",
-13062 => x"C0C0BFF9B0C082A4",
-13061 => x"C0C0BFF9B0C082F9",
-13060 => x"C0C0BFF9B0C082C0",
-13059 => x"C0C0BFF9B0C09290",
-13058 => x"C0C0BFF9B0C09280",
-13057 => x"C0C0BFF9B0C092F8",
-13056 => x"C0C0BFF9B0C09282",
-13055 => x"C0C0BFF9B0C09292",
-13054 => x"C0C0BFF9B0C09299",
-13053 => x"C0C0BFF9B0C092B0",
-13052 => x"C0C0BFF9B0C092A4",
-13051 => x"C0C0BFF9B0C092F9",
-13050 => x"C0C0BFF9B0C092C0",
-13049 => x"C0C0BFF9B0C09990",
-13048 => x"C0C0BFF9B0C09980",
-13047 => x"C0C0BFF9B0C099F8",
-13046 => x"C0C0BFF9B0C09982",
-13045 => x"C0C0BFF9B0C09992",
-13044 => x"C0C0BFF9B0C09999",
-13043 => x"C0C0BFF9B0C099B0",
-13042 => x"C0C0BFF9B0C099A4",
-13041 => x"C0C0BFF9B0C099F9",
-13040 => x"C0C0BFF9B0C099C0",
-13039 => x"C0C0BFF9B0C0B090",
-13038 => x"C0C0BFF9B0C0B080",
-13037 => x"C0C0BFF9B0C0B0F8",
-13036 => x"C0C0BFF9B0C0B082",
-13035 => x"C0C0BFF9B0C0B092",
-13034 => x"C0C0BFF9B0C0B099",
-13033 => x"C0C0BFF9B0C0B0B0",
-13032 => x"C0C0BFF9B0C0B0A4",
-13031 => x"C0C0BFF9B0C0B0F9",
-13030 => x"C0C0BFF9B0C0B0C0",
-13029 => x"C0C0BFF9B0C0A490",
-13028 => x"C0C0BFF9B0C0A480",
-13027 => x"C0C0BFF9B0C0A4F8",
-13026 => x"C0C0BFF9B0C0A482",
-13025 => x"C0C0BFF9B0C0A492",
-13024 => x"C0C0BFF9B0C0A499",
-13023 => x"C0C0BFF9B0C0A4B0",
-13022 => x"C0C0BFF9B0C0A4A4",
-13021 => x"C0C0BFF9B0C0A4F9",
-13020 => x"C0C0BFF9B0C0A4C0",
-13019 => x"C0C0BFF9B0C0F990",
-13018 => x"C0C0BFF9B0C0F980",
-13017 => x"C0C0BFF9B0C0F9F8",
-13016 => x"C0C0BFF9B0C0F982",
-13015 => x"C0C0BFF9B0C0F992",
-13014 => x"C0C0BFF9B0C0F999",
-13013 => x"C0C0BFF9B0C0F9B0",
-13012 => x"C0C0BFF9B0C0F9A4",
-13011 => x"C0C0BFF9B0C0F9F9",
-13010 => x"C0C0BFF9B0C0F9C0",
-13009 => x"C0C0BFF9B0C0C090",
-13008 => x"C0C0BFF9B0C0C080",
-13007 => x"C0C0BFF9B0C0C0F8",
-13006 => x"C0C0BFF9B0C0C082",
-13005 => x"C0C0BFF9B0C0C092",
-13004 => x"C0C0BFF9B0C0C099",
-13003 => x"C0C0BFF9B0C0C0B0",
-13002 => x"C0C0BFF9B0C0C0A4",
-13001 => x"C0C0BFF9B0C0C0F9",
-13000 => x"C0C0BFF9B0C0C0C0",
-12999 => x"C0C0BFF9A4909090",
-12998 => x"C0C0BFF9A4909080",
-12997 => x"C0C0BFF9A49090F8",
-12996 => x"C0C0BFF9A4909082",
-12995 => x"C0C0BFF9A4909092",
-12994 => x"C0C0BFF9A4909099",
-12993 => x"C0C0BFF9A49090B0",
-12992 => x"C0C0BFF9A49090A4",
-12991 => x"C0C0BFF9A49090F9",
-12990 => x"C0C0BFF9A49090C0",
-12989 => x"C0C0BFF9A4908090",
-12988 => x"C0C0BFF9A4908080",
-12987 => x"C0C0BFF9A49080F8",
-12986 => x"C0C0BFF9A4908082",
-12985 => x"C0C0BFF9A4908092",
-12984 => x"C0C0BFF9A4908099",
-12983 => x"C0C0BFF9A49080B0",
-12982 => x"C0C0BFF9A49080A4",
-12981 => x"C0C0BFF9A49080F9",
-12980 => x"C0C0BFF9A49080C0",
-12979 => x"C0C0BFF9A490F890",
-12978 => x"C0C0BFF9A490F880",
-12977 => x"C0C0BFF9A490F8F8",
-12976 => x"C0C0BFF9A490F882",
-12975 => x"C0C0BFF9A490F892",
-12974 => x"C0C0BFF9A490F899",
-12973 => x"C0C0BFF9A490F8B0",
-12972 => x"C0C0BFF9A490F8A4",
-12971 => x"C0C0BFF9A490F8F9",
-12970 => x"C0C0BFF9A490F8C0",
-12969 => x"C0C0BFF9A4908290",
-12968 => x"C0C0BFF9A4908280",
-12967 => x"C0C0BFF9A49082F8",
-12966 => x"C0C0BFF9A4908282",
-12965 => x"C0C0BFF9A4908292",
-12964 => x"C0C0BFF9A4908299",
-12963 => x"C0C0BFF9A49082B0",
-12962 => x"C0C0BFF9A49082A4",
-12961 => x"C0C0BFF9A49082F9",
-12960 => x"C0C0BFF9A49082C0",
-12959 => x"C0C0BFF9A4909290",
-12958 => x"C0C0BFF9A4909280",
-12957 => x"C0C0BFF9A49092F8",
-12956 => x"C0C0BFF9A4909282",
-12955 => x"C0C0BFF9A4909292",
-12954 => x"C0C0BFF9A4909299",
-12953 => x"C0C0BFF9A49092B0",
-12952 => x"C0C0BFF9A49092A4",
-12951 => x"C0C0BFF9A49092F9",
-12950 => x"C0C0BFF9A49092C0",
-12949 => x"C0C0BFF9A4909990",
-12948 => x"C0C0BFF9A4909980",
-12947 => x"C0C0BFF9A49099F8",
-12946 => x"C0C0BFF9A4909982",
-12945 => x"C0C0BFF9A4909992",
-12944 => x"C0C0BFF9A4909999",
-12943 => x"C0C0BFF9A49099B0",
-12942 => x"C0C0BFF9A49099A4",
-12941 => x"C0C0BFF9A49099F9",
-12940 => x"C0C0BFF9A49099C0",
-12939 => x"C0C0BFF9A490B090",
-12938 => x"C0C0BFF9A490B080",
-12937 => x"C0C0BFF9A490B0F8",
-12936 => x"C0C0BFF9A490B082",
-12935 => x"C0C0BFF9A490B092",
-12934 => x"C0C0BFF9A490B099",
-12933 => x"C0C0BFF9A490B0B0",
-12932 => x"C0C0BFF9A490B0A4",
-12931 => x"C0C0BFF9A490B0F9",
-12930 => x"C0C0BFF9A490B0C0",
-12929 => x"C0C0BFF9A490A490",
-12928 => x"C0C0BFF9A490A480",
-12927 => x"C0C0BFF9A490A4F8",
-12926 => x"C0C0BFF9A490A482",
-12925 => x"C0C0BFF9A490A492",
-12924 => x"C0C0BFF9A490A499",
-12923 => x"C0C0BFF9A490A4B0",
-12922 => x"C0C0BFF9A490A4A4",
-12921 => x"C0C0BFF9A490A4F9",
-12920 => x"C0C0BFF9A490A4C0",
-12919 => x"C0C0BFF9A490F990",
-12918 => x"C0C0BFF9A490F980",
-12917 => x"C0C0BFF9A490F9F8",
-12916 => x"C0C0BFF9A490F982",
-12915 => x"C0C0BFF9A490F992",
-12914 => x"C0C0BFF9A490F999",
-12913 => x"C0C0BFF9A490F9B0",
-12912 => x"C0C0BFF9A490F9A4",
-12911 => x"C0C0BFF9A490F9F9",
-12910 => x"C0C0BFF9A490F9C0",
-12909 => x"C0C0BFF9A490C090",
-12908 => x"C0C0BFF9A490C080",
-12907 => x"C0C0BFF9A490C0F8",
-12906 => x"C0C0BFF9A490C082",
-12905 => x"C0C0BFF9A490C092",
-12904 => x"C0C0BFF9A490C099",
-12903 => x"C0C0BFF9A490C0B0",
-12902 => x"C0C0BFF9A490C0A4",
-12901 => x"C0C0BFF9A490C0F9",
-12900 => x"C0C0BFF9A490C0C0",
-12899 => x"C0C0BFF9A4809090",
-12898 => x"C0C0BFF9A4809080",
-12897 => x"C0C0BFF9A48090F8",
-12896 => x"C0C0BFF9A4809082",
-12895 => x"C0C0BFF9A4809092",
-12894 => x"C0C0BFF9A4809099",
-12893 => x"C0C0BFF9A48090B0",
-12892 => x"C0C0BFF9A48090A4",
-12891 => x"C0C0BFF9A48090F9",
-12890 => x"C0C0BFF9A48090C0",
-12889 => x"C0C0BFF9A4808090",
-12888 => x"C0C0BFF9A4808080",
-12887 => x"C0C0BFF9A48080F8",
-12886 => x"C0C0BFF9A4808082",
-12885 => x"C0C0BFF9A4808092",
-12884 => x"C0C0BFF9A4808099",
-12883 => x"C0C0BFF9A48080B0",
-12882 => x"C0C0BFF9A48080A4",
-12881 => x"C0C0BFF9A48080F9",
-12880 => x"C0C0BFF9A48080C0",
-12879 => x"C0C0BFF9A480F890",
-12878 => x"C0C0BFF9A480F880",
-12877 => x"C0C0BFF9A480F8F8",
-12876 => x"C0C0BFF9A480F882",
-12875 => x"C0C0BFF9A480F892",
-12874 => x"C0C0BFF9A480F899",
-12873 => x"C0C0BFF9A480F8B0",
-12872 => x"C0C0BFF9A480F8A4",
-12871 => x"C0C0BFF9A480F8F9",
-12870 => x"C0C0BFF9A480F8C0",
-12869 => x"C0C0BFF9A4808290",
-12868 => x"C0C0BFF9A4808280",
-12867 => x"C0C0BFF9A48082F8",
-12866 => x"C0C0BFF9A4808282",
-12865 => x"C0C0BFF9A4808292",
-12864 => x"C0C0BFF9A4808299",
-12863 => x"C0C0BFF9A48082B0",
-12862 => x"C0C0BFF9A48082A4",
-12861 => x"C0C0BFF9A48082F9",
-12860 => x"C0C0BFF9A48082C0",
-12859 => x"C0C0BFF9A4809290",
-12858 => x"C0C0BFF9A4809280",
-12857 => x"C0C0BFF9A48092F8",
-12856 => x"C0C0BFF9A4809282",
-12855 => x"C0C0BFF9A4809292",
-12854 => x"C0C0BFF9A4809299",
-12853 => x"C0C0BFF9A48092B0",
-12852 => x"C0C0BFF9A48092A4",
-12851 => x"C0C0BFF9A48092F9",
-12850 => x"C0C0BFF9A48092C0",
-12849 => x"C0C0BFF9A4809990",
-12848 => x"C0C0BFF9A4809980",
-12847 => x"C0C0BFF9A48099F8",
-12846 => x"C0C0BFF9A4809982",
-12845 => x"C0C0BFF9A4809992",
-12844 => x"C0C0BFF9A4809999",
-12843 => x"C0C0BFF9A48099B0",
-12842 => x"C0C0BFF9A48099A4",
-12841 => x"C0C0BFF9A48099F9",
-12840 => x"C0C0BFF9A48099C0",
-12839 => x"C0C0BFF9A480B090",
-12838 => x"C0C0BFF9A480B080",
-12837 => x"C0C0BFF9A480B0F8",
-12836 => x"C0C0BFF9A480B082",
-12835 => x"C0C0BFF9A480B092",
-12834 => x"C0C0BFF9A480B099",
-12833 => x"C0C0BFF9A480B0B0",
-12832 => x"C0C0BFF9A480B0A4",
-12831 => x"C0C0BFF9A480B0F9",
-12830 => x"C0C0BFF9A480B0C0",
-12829 => x"C0C0BFF9A480A490",
-12828 => x"C0C0BFF9A480A480",
-12827 => x"C0C0BFF9A480A4F8",
-12826 => x"C0C0BFF9A480A482",
-12825 => x"C0C0BFF9A480A492",
-12824 => x"C0C0BFF9A480A499",
-12823 => x"C0C0BFF9A480A4B0",
-12822 => x"C0C0BFF9A480A4A4",
-12821 => x"C0C0BFF9A480A4F9",
-12820 => x"C0C0BFF9A480A4C0",
-12819 => x"C0C0BFF9A480F990",
-12818 => x"C0C0BFF9A480F980",
-12817 => x"C0C0BFF9A480F9F8",
-12816 => x"C0C0BFF9A480F982",
-12815 => x"C0C0BFF9A480F992",
-12814 => x"C0C0BFF9A480F999",
-12813 => x"C0C0BFF9A480F9B0",
-12812 => x"C0C0BFF9A480F9A4",
-12811 => x"C0C0BFF9A480F9F9",
-12810 => x"C0C0BFF9A480F9C0",
-12809 => x"C0C0BFF9A480C090",
-12808 => x"C0C0BFF9A480C080",
-12807 => x"C0C0BFF9A480C0F8",
-12806 => x"C0C0BFF9A480C082",
-12805 => x"C0C0BFF9A480C092",
-12804 => x"C0C0BFF9A480C099",
-12803 => x"C0C0BFF9A480C0B0",
-12802 => x"C0C0BFF9A480C0A4",
-12801 => x"C0C0BFF9A480C0F9",
-12800 => x"C0C0BFF9A480C0C0",
-12799 => x"C0C0BFF9A4F89090",
-12798 => x"C0C0BFF9A4F89080",
-12797 => x"C0C0BFF9A4F890F8",
-12796 => x"C0C0BFF9A4F89082",
-12795 => x"C0C0BFF9A4F89092",
-12794 => x"C0C0BFF9A4F89099",
-12793 => x"C0C0BFF9A4F890B0",
-12792 => x"C0C0BFF9A4F890A4",
-12791 => x"C0C0BFF9A4F890F9",
-12790 => x"C0C0BFF9A4F890C0",
-12789 => x"C0C0BFF9A4F88090",
-12788 => x"C0C0BFF9A4F88080",
-12787 => x"C0C0BFF9A4F880F8",
-12786 => x"C0C0BFF9A4F88082",
-12785 => x"C0C0BFF9A4F88092",
-12784 => x"C0C0BFF9A4F88099",
-12783 => x"C0C0BFF9A4F880B0",
-12782 => x"C0C0BFF9A4F880A4",
-12781 => x"C0C0BFF9A4F880F9",
-12780 => x"C0C0BFF9A4F880C0",
-12779 => x"C0C0BFF9A4F8F890",
-12778 => x"C0C0BFF9A4F8F880",
-12777 => x"C0C0BFF9A4F8F8F8",
-12776 => x"C0C0BFF9A4F8F882",
-12775 => x"C0C0BFF9A4F8F892",
-12774 => x"C0C0BFF9A4F8F899",
-12773 => x"C0C0BFF9A4F8F8B0",
-12772 => x"C0C0BFF9A4F8F8A4",
-12771 => x"C0C0BFF9A4F8F8F9",
-12770 => x"C0C0BFF9A4F8F8C0",
-12769 => x"C0C0BFF9A4F88290",
-12768 => x"C0C0BFF9A4F88280",
-12767 => x"C0C0BFF9A4F882F8",
-12766 => x"C0C0BFF9A4F88282",
-12765 => x"C0C0BFF9A4F88292",
-12764 => x"C0C0BFF9A4F88299",
-12763 => x"C0C0BFF9A4F882B0",
-12762 => x"C0C0BFF9A4F882A4",
-12761 => x"C0C0BFF9A4F882F9",
-12760 => x"C0C0BFF9A4F882C0",
-12759 => x"C0C0BFF9A4F89290",
-12758 => x"C0C0BFF9A4F89280",
-12757 => x"C0C0BFF9A4F892F8",
-12756 => x"C0C0BFF9A4F89282",
-12755 => x"C0C0BFF9A4F89292",
-12754 => x"C0C0BFF9A4F89299",
-12753 => x"C0C0BFF9A4F892B0",
-12752 => x"C0C0BFF9A4F892A4",
-12751 => x"C0C0BFF9A4F892F9",
-12750 => x"C0C0BFF9A4F892C0",
-12749 => x"C0C0BFF9A4F89990",
-12748 => x"C0C0BFF9A4F89980",
-12747 => x"C0C0BFF9A4F899F8",
-12746 => x"C0C0BFF9A4F89982",
-12745 => x"C0C0BFF9A4F89992",
-12744 => x"C0C0BFF9A4F89999",
-12743 => x"C0C0BFF9A4F899B0",
-12742 => x"C0C0BFF9A4F899A4",
-12741 => x"C0C0BFF9A4F899F9",
-12740 => x"C0C0BFF9A4F899C0",
-12739 => x"C0C0BFF9A4F8B090",
-12738 => x"C0C0BFF9A4F8B080",
-12737 => x"C0C0BFF9A4F8B0F8",
-12736 => x"C0C0BFF9A4F8B082",
-12735 => x"C0C0BFF9A4F8B092",
-12734 => x"C0C0BFF9A4F8B099",
-12733 => x"C0C0BFF9A4F8B0B0",
-12732 => x"C0C0BFF9A4F8B0A4",
-12731 => x"C0C0BFF9A4F8B0F9",
-12730 => x"C0C0BFF9A4F8B0C0",
-12729 => x"C0C0BFF9A4F8A490",
-12728 => x"C0C0BFF9A4F8A480",
-12727 => x"C0C0BFF9A4F8A4F8",
-12726 => x"C0C0BFF9A4F8A482",
-12725 => x"C0C0BFF9A4F8A492",
-12724 => x"C0C0BFF9A4F8A499",
-12723 => x"C0C0BFF9A4F8A4B0",
-12722 => x"C0C0BFF9A4F8A4A4",
-12721 => x"C0C0BFF9A4F8A4F9",
-12720 => x"C0C0BFF9A4F8A4C0",
-12719 => x"C0C0BFF9A4F8F990",
-12718 => x"C0C0BFF9A4F8F980",
-12717 => x"C0C0BFF9A4F8F9F8",
-12716 => x"C0C0BFF9A4F8F982",
-12715 => x"C0C0BFF9A4F8F992",
-12714 => x"C0C0BFF9A4F8F999",
-12713 => x"C0C0BFF9A4F8F9B0",
-12712 => x"C0C0BFF9A4F8F9A4",
-12711 => x"C0C0BFF9A4F8F9F9",
-12710 => x"C0C0BFF9A4F8F9C0",
-12709 => x"C0C0BFF9A4F8C090",
-12708 => x"C0C0BFF9A4F8C080",
-12707 => x"C0C0BFF9A4F8C0F8",
-12706 => x"C0C0BFF9A4F8C082",
-12705 => x"C0C0BFF9A4F8C092",
-12704 => x"C0C0BFF9A4F8C099",
-12703 => x"C0C0BFF9A4F8C0B0",
-12702 => x"C0C0BFF9A4F8C0A4",
-12701 => x"C0C0BFF9A4F8C0F9",
-12700 => x"C0C0BFF9A4F8C0C0",
-12699 => x"C0C0BFF9A4829090",
-12698 => x"C0C0BFF9A4829080",
-12697 => x"C0C0BFF9A48290F8",
-12696 => x"C0C0BFF9A4829082",
-12695 => x"C0C0BFF9A4829092",
-12694 => x"C0C0BFF9A4829099",
-12693 => x"C0C0BFF9A48290B0",
-12692 => x"C0C0BFF9A48290A4",
-12691 => x"C0C0BFF9A48290F9",
-12690 => x"C0C0BFF9A48290C0",
-12689 => x"C0C0BFF9A4828090",
-12688 => x"C0C0BFF9A4828080",
-12687 => x"C0C0BFF9A48280F8",
-12686 => x"C0C0BFF9A4828082",
-12685 => x"C0C0BFF9A4828092",
-12684 => x"C0C0BFF9A4828099",
-12683 => x"C0C0BFF9A48280B0",
-12682 => x"C0C0BFF9A48280A4",
-12681 => x"C0C0BFF9A48280F9",
-12680 => x"C0C0BFF9A48280C0",
-12679 => x"C0C0BFF9A482F890",
-12678 => x"C0C0BFF9A482F880",
-12677 => x"C0C0BFF9A482F8F8",
-12676 => x"C0C0BFF9A482F882",
-12675 => x"C0C0BFF9A482F892",
-12674 => x"C0C0BFF9A482F899",
-12673 => x"C0C0BFF9A482F8B0",
-12672 => x"C0C0BFF9A482F8A4",
-12671 => x"C0C0BFF9A482F8F9",
-12670 => x"C0C0BFF9A482F8C0",
-12669 => x"C0C0BFF9A4828290",
-12668 => x"C0C0BFF9A4828280",
-12667 => x"C0C0BFF9A48282F8",
-12666 => x"C0C0BFF9A4828282",
-12665 => x"C0C0BFF9A4828292",
-12664 => x"C0C0BFF9A4828299",
-12663 => x"C0C0BFF9A48282B0",
-12662 => x"C0C0BFF9A48282A4",
-12661 => x"C0C0BFF9A48282F9",
-12660 => x"C0C0BFF9A48282C0",
-12659 => x"C0C0BFF9A4829290",
-12658 => x"C0C0BFF9A4829280",
-12657 => x"C0C0BFF9A48292F8",
-12656 => x"C0C0BFF9A4829282",
-12655 => x"C0C0BFF9A4829292",
-12654 => x"C0C0BFF9A4829299",
-12653 => x"C0C0BFF9A48292B0",
-12652 => x"C0C0BFF9A48292A4",
-12651 => x"C0C0BFF9A48292F9",
-12650 => x"C0C0BFF9A48292C0",
-12649 => x"C0C0BFF9A4829990",
-12648 => x"C0C0BFF9A4829980",
-12647 => x"C0C0BFF9A48299F8",
-12646 => x"C0C0BFF9A4829982",
-12645 => x"C0C0BFF9A4829992",
-12644 => x"C0C0BFF9A4829999",
-12643 => x"C0C0BFF9A48299B0",
-12642 => x"C0C0BFF9A48299A4",
-12641 => x"C0C0BFF9A48299F9",
-12640 => x"C0C0BFF9A48299C0",
-12639 => x"C0C0BFF9A482B090",
-12638 => x"C0C0BFF9A482B080",
-12637 => x"C0C0BFF9A482B0F8",
-12636 => x"C0C0BFF9A482B082",
-12635 => x"C0C0BFF9A482B092",
-12634 => x"C0C0BFF9A482B099",
-12633 => x"C0C0BFF9A482B0B0",
-12632 => x"C0C0BFF9A482B0A4",
-12631 => x"C0C0BFF9A482B0F9",
-12630 => x"C0C0BFF9A482B0C0",
-12629 => x"C0C0BFF9A482A490",
-12628 => x"C0C0BFF9A482A480",
-12627 => x"C0C0BFF9A482A4F8",
-12626 => x"C0C0BFF9A482A482",
-12625 => x"C0C0BFF9A482A492",
-12624 => x"C0C0BFF9A482A499",
-12623 => x"C0C0BFF9A482A4B0",
-12622 => x"C0C0BFF9A482A4A4",
-12621 => x"C0C0BFF9A482A4F9",
-12620 => x"C0C0BFF9A482A4C0",
-12619 => x"C0C0BFF9A482F990",
-12618 => x"C0C0BFF9A482F980",
-12617 => x"C0C0BFF9A482F9F8",
-12616 => x"C0C0BFF9A482F982",
-12615 => x"C0C0BFF9A482F992",
-12614 => x"C0C0BFF9A482F999",
-12613 => x"C0C0BFF9A482F9B0",
-12612 => x"C0C0BFF9A482F9A4",
-12611 => x"C0C0BFF9A482F9F9",
-12610 => x"C0C0BFF9A482F9C0",
-12609 => x"C0C0BFF9A482C090",
-12608 => x"C0C0BFF9A482C080",
-12607 => x"C0C0BFF9A482C0F8",
-12606 => x"C0C0BFF9A482C082",
-12605 => x"C0C0BFF9A482C092",
-12604 => x"C0C0BFF9A482C099",
-12603 => x"C0C0BFF9A482C0B0",
-12602 => x"C0C0BFF9A482C0A4",
-12601 => x"C0C0BFF9A482C0F9",
-12600 => x"C0C0BFF9A482C0C0",
-12599 => x"C0C0BFF9A4929090",
-12598 => x"C0C0BFF9A4929080",
-12597 => x"C0C0BFF9A49290F8",
-12596 => x"C0C0BFF9A4929082",
-12595 => x"C0C0BFF9A4929092",
-12594 => x"C0C0BFF9A4929099",
-12593 => x"C0C0BFF9A49290B0",
-12592 => x"C0C0BFF9A49290A4",
-12591 => x"C0C0BFF9A49290F9",
-12590 => x"C0C0BFF9A49290C0",
-12589 => x"C0C0BFF9A4928090",
-12588 => x"C0C0BFF9A4928080",
-12587 => x"C0C0BFF9A49280F8",
-12586 => x"C0C0BFF9A4928082",
-12585 => x"C0C0BFF9A4928092",
-12584 => x"C0C0BFF9A4928099",
-12583 => x"C0C0BFF9A49280B0",
-12582 => x"C0C0BFF9A49280A4",
-12581 => x"C0C0BFF9A49280F9",
-12580 => x"C0C0BFF9A49280C0",
-12579 => x"C0C0BFF9A492F890",
-12578 => x"C0C0BFF9A492F880",
-12577 => x"C0C0BFF9A492F8F8",
-12576 => x"C0C0BFF9A492F882",
-12575 => x"C0C0BFF9A492F892",
-12574 => x"C0C0BFF9A492F899",
-12573 => x"C0C0BFF9A492F8B0",
-12572 => x"C0C0BFF9A492F8A4",
-12571 => x"C0C0BFF9A492F8F9",
-12570 => x"C0C0BFF9A492F8C0",
-12569 => x"C0C0BFF9A4928290",
-12568 => x"C0C0BFF9A4928280",
-12567 => x"C0C0BFF9A49282F8",
-12566 => x"C0C0BFF9A4928282",
-12565 => x"C0C0BFF9A4928292",
-12564 => x"C0C0BFF9A4928299",
-12563 => x"C0C0BFF9A49282B0",
-12562 => x"C0C0BFF9A49282A4",
-12561 => x"C0C0BFF9A49282F9",
-12560 => x"C0C0BFF9A49282C0",
-12559 => x"C0C0BFF9A4929290",
-12558 => x"C0C0BFF9A4929280",
-12557 => x"C0C0BFF9A49292F8",
-12556 => x"C0C0BFF9A4929282",
-12555 => x"C0C0BFF9A4929292",
-12554 => x"C0C0BFF9A4929299",
-12553 => x"C0C0BFF9A49292B0",
-12552 => x"C0C0BFF9A49292A4",
-12551 => x"C0C0BFF9A49292F9",
-12550 => x"C0C0BFF9A49292C0",
-12549 => x"C0C0BFF9A4929990",
-12548 => x"C0C0BFF9A4929980",
-12547 => x"C0C0BFF9A49299F8",
-12546 => x"C0C0BFF9A4929982",
-12545 => x"C0C0BFF9A4929992",
-12544 => x"C0C0BFF9A4929999",
-12543 => x"C0C0BFF9A49299B0",
-12542 => x"C0C0BFF9A49299A4",
-12541 => x"C0C0BFF9A49299F9",
-12540 => x"C0C0BFF9A49299C0",
-12539 => x"C0C0BFF9A492B090",
-12538 => x"C0C0BFF9A492B080",
-12537 => x"C0C0BFF9A492B0F8",
-12536 => x"C0C0BFF9A492B082",
-12535 => x"C0C0BFF9A492B092",
-12534 => x"C0C0BFF9A492B099",
-12533 => x"C0C0BFF9A492B0B0",
-12532 => x"C0C0BFF9A492B0A4",
-12531 => x"C0C0BFF9A492B0F9",
-12530 => x"C0C0BFF9A492B0C0",
-12529 => x"C0C0BFF9A492A490",
-12528 => x"C0C0BFF9A492A480",
-12527 => x"C0C0BFF9A492A4F8",
-12526 => x"C0C0BFF9A492A482",
-12525 => x"C0C0BFF9A492A492",
-12524 => x"C0C0BFF9A492A499",
-12523 => x"C0C0BFF9A492A4B0",
-12522 => x"C0C0BFF9A492A4A4",
-12521 => x"C0C0BFF9A492A4F9",
-12520 => x"C0C0BFF9A492A4C0",
-12519 => x"C0C0BFF9A492F990",
-12518 => x"C0C0BFF9A492F980",
-12517 => x"C0C0BFF9A492F9F8",
-12516 => x"C0C0BFF9A492F982",
-12515 => x"C0C0BFF9A492F992",
-12514 => x"C0C0BFF9A492F999",
-12513 => x"C0C0BFF9A492F9B0",
-12512 => x"C0C0BFF9A492F9A4",
-12511 => x"C0C0BFF9A492F9F9",
-12510 => x"C0C0BFF9A492F9C0",
-12509 => x"C0C0BFF9A492C090",
-12508 => x"C0C0BFF9A492C080",
-12507 => x"C0C0BFF9A492C0F8",
-12506 => x"C0C0BFF9A492C082",
-12505 => x"C0C0BFF9A492C092",
-12504 => x"C0C0BFF9A492C099",
-12503 => x"C0C0BFF9A492C0B0",
-12502 => x"C0C0BFF9A492C0A4",
-12501 => x"C0C0BFF9A492C0F9",
-12500 => x"C0C0BFF9A492C0C0",
-12499 => x"C0C0BFF9A4999090",
-12498 => x"C0C0BFF9A4999080",
-12497 => x"C0C0BFF9A49990F8",
-12496 => x"C0C0BFF9A4999082",
-12495 => x"C0C0BFF9A4999092",
-12494 => x"C0C0BFF9A4999099",
-12493 => x"C0C0BFF9A49990B0",
-12492 => x"C0C0BFF9A49990A4",
-12491 => x"C0C0BFF9A49990F9",
-12490 => x"C0C0BFF9A49990C0",
-12489 => x"C0C0BFF9A4998090",
-12488 => x"C0C0BFF9A4998080",
-12487 => x"C0C0BFF9A49980F8",
-12486 => x"C0C0BFF9A4998082",
-12485 => x"C0C0BFF9A4998092",
-12484 => x"C0C0BFF9A4998099",
-12483 => x"C0C0BFF9A49980B0",
-12482 => x"C0C0BFF9A49980A4",
-12481 => x"C0C0BFF9A49980F9",
-12480 => x"C0C0BFF9A49980C0",
-12479 => x"C0C0BFF9A499F890",
-12478 => x"C0C0BFF9A499F880",
-12477 => x"C0C0BFF9A499F8F8",
-12476 => x"C0C0BFF9A499F882",
-12475 => x"C0C0BFF9A499F892",
-12474 => x"C0C0BFF9A499F899",
-12473 => x"C0C0BFF9A499F8B0",
-12472 => x"C0C0BFF9A499F8A4",
-12471 => x"C0C0BFF9A499F8F9",
-12470 => x"C0C0BFF9A499F8C0",
-12469 => x"C0C0BFF9A4998290",
-12468 => x"C0C0BFF9A4998280",
-12467 => x"C0C0BFF9A49982F8",
-12466 => x"C0C0BFF9A4998282",
-12465 => x"C0C0BFF9A4998292",
-12464 => x"C0C0BFF9A4998299",
-12463 => x"C0C0BFF9A49982B0",
-12462 => x"C0C0BFF9A49982A4",
-12461 => x"C0C0BFF9A49982F9",
-12460 => x"C0C0BFF9A49982C0",
-12459 => x"C0C0BFF9A4999290",
-12458 => x"C0C0BFF9A4999280",
-12457 => x"C0C0BFF9A49992F8",
-12456 => x"C0C0BFF9A4999282",
-12455 => x"C0C0BFF9A4999292",
-12454 => x"C0C0BFF9A4999299",
-12453 => x"C0C0BFF9A49992B0",
-12452 => x"C0C0BFF9A49992A4",
-12451 => x"C0C0BFF9A49992F9",
-12450 => x"C0C0BFF9A49992C0",
-12449 => x"C0C0BFF9A4999990",
-12448 => x"C0C0BFF9A4999980",
-12447 => x"C0C0BFF9A49999F8",
-12446 => x"C0C0BFF9A4999982",
-12445 => x"C0C0BFF9A4999992",
-12444 => x"C0C0BFF9A4999999",
-12443 => x"C0C0BFF9A49999B0",
-12442 => x"C0C0BFF9A49999A4",
-12441 => x"C0C0BFF9A49999F9",
-12440 => x"C0C0BFF9A49999C0",
-12439 => x"C0C0BFF9A499B090",
-12438 => x"C0C0BFF9A499B080",
-12437 => x"C0C0BFF9A499B0F8",
-12436 => x"C0C0BFF9A499B082",
-12435 => x"C0C0BFF9A499B092",
-12434 => x"C0C0BFF9A499B099",
-12433 => x"C0C0BFF9A499B0B0",
-12432 => x"C0C0BFF9A499B0A4",
-12431 => x"C0C0BFF9A499B0F9",
-12430 => x"C0C0BFF9A499B0C0",
-12429 => x"C0C0BFF9A499A490",
-12428 => x"C0C0BFF9A499A480",
-12427 => x"C0C0BFF9A499A4F8",
-12426 => x"C0C0BFF9A499A482",
-12425 => x"C0C0BFF9A499A492",
-12424 => x"C0C0BFF9A499A499",
-12423 => x"C0C0BFF9A499A4B0",
-12422 => x"C0C0BFF9A499A4A4",
-12421 => x"C0C0BFF9A499A4F9",
-12420 => x"C0C0BFF9A499A4C0",
-12419 => x"C0C0BFF9A499F990",
-12418 => x"C0C0BFF9A499F980",
-12417 => x"C0C0BFF9A499F9F8",
-12416 => x"C0C0BFF9A499F982",
-12415 => x"C0C0BFF9A499F992",
-12414 => x"C0C0BFF9A499F999",
-12413 => x"C0C0BFF9A499F9B0",
-12412 => x"C0C0BFF9A499F9A4",
-12411 => x"C0C0BFF9A499F9F9",
-12410 => x"C0C0BFF9A499F9C0",
-12409 => x"C0C0BFF9A499C090",
-12408 => x"C0C0BFF9A499C080",
-12407 => x"C0C0BFF9A499C0F8",
-12406 => x"C0C0BFF9A499C082",
-12405 => x"C0C0BFF9A499C092",
-12404 => x"C0C0BFF9A499C099",
-12403 => x"C0C0BFF9A499C0B0",
-12402 => x"C0C0BFF9A499C0A4",
-12401 => x"C0C0BFF9A499C0F9",
-12400 => x"C0C0BFF9A499C0C0",
-12399 => x"C0C0BFF9A4B09090",
-12398 => x"C0C0BFF9A4B09080",
-12397 => x"C0C0BFF9A4B090F8",
-12396 => x"C0C0BFF9A4B09082",
-12395 => x"C0C0BFF9A4B09092",
-12394 => x"C0C0BFF9A4B09099",
-12393 => x"C0C0BFF9A4B090B0",
-12392 => x"C0C0BFF9A4B090A4",
-12391 => x"C0C0BFF9A4B090F9",
-12390 => x"C0C0BFF9A4B090C0",
-12389 => x"C0C0BFF9A4B08090",
-12388 => x"C0C0BFF9A4B08080",
-12387 => x"C0C0BFF9A4B080F8",
-12386 => x"C0C0BFF9A4B08082",
-12385 => x"C0C0BFF9A4B08092",
-12384 => x"C0C0BFF9A4B08099",
-12383 => x"C0C0BFF9A4B080B0",
-12382 => x"C0C0BFF9A4B080A4",
-12381 => x"C0C0BFF9A4B080F9",
-12380 => x"C0C0BFF9A4B080C0",
-12379 => x"C0C0BFF9A4B0F890",
-12378 => x"C0C0BFF9A4B0F880",
-12377 => x"C0C0BFF9A4B0F8F8",
-12376 => x"C0C0BFF9A4B0F882",
-12375 => x"C0C0BFF9A4B0F892",
-12374 => x"C0C0BFF9A4B0F899",
-12373 => x"C0C0BFF9A4B0F8B0",
-12372 => x"C0C0BFF9A4B0F8A4",
-12371 => x"C0C0BFF9A4B0F8F9",
-12370 => x"C0C0BFF9A4B0F8C0",
-12369 => x"C0C0BFF9A4B08290",
-12368 => x"C0C0BFF9A4B08280",
-12367 => x"C0C0BFF9A4B082F8",
-12366 => x"C0C0BFF9A4B08282",
-12365 => x"C0C0BFF9A4B08292",
-12364 => x"C0C0BFF9A4B08299",
-12363 => x"C0C0BFF9A4B082B0",
-12362 => x"C0C0BFF9A4B082A4",
-12361 => x"C0C0BFF9A4B082F9",
-12360 => x"C0C0BFF9A4B082C0",
-12359 => x"C0C0BFF9A4B09290",
-12358 => x"C0C0BFF9A4B09280",
-12357 => x"C0C0BFF9A4B092F8",
-12356 => x"C0C0BFF9A4B09282",
-12355 => x"C0C0BFF9A4B09292",
-12354 => x"C0C0BFF9A4B09299",
-12353 => x"C0C0BFF9A4B092B0",
-12352 => x"C0C0BFF9A4B092A4",
-12351 => x"C0C0BFF9A4B092F9",
-12350 => x"C0C0BFF9A4B092C0",
-12349 => x"C0C0BFF9A4B09990",
-12348 => x"C0C0BFF9A4B09980",
-12347 => x"C0C0BFF9A4B099F8",
-12346 => x"C0C0BFF9A4B09982",
-12345 => x"C0C0BFF9A4B09992",
-12344 => x"C0C0BFF9A4B09999",
-12343 => x"C0C0BFF9A4B099B0",
-12342 => x"C0C0BFF9A4B099A4",
-12341 => x"C0C0BFF9A4B099F9",
-12340 => x"C0C0BFF9A4B099C0",
-12339 => x"C0C0BFF9A4B0B090",
-12338 => x"C0C0BFF9A4B0B080",
-12337 => x"C0C0BFF9A4B0B0F8",
-12336 => x"C0C0BFF9A4B0B082",
-12335 => x"C0C0BFF9A4B0B092",
-12334 => x"C0C0BFF9A4B0B099",
-12333 => x"C0C0BFF9A4B0B0B0",
-12332 => x"C0C0BFF9A4B0B0A4",
-12331 => x"C0C0BFF9A4B0B0F9",
-12330 => x"C0C0BFF9A4B0B0C0",
-12329 => x"C0C0BFF9A4B0A490",
-12328 => x"C0C0BFF9A4B0A480",
-12327 => x"C0C0BFF9A4B0A4F8",
-12326 => x"C0C0BFF9A4B0A482",
-12325 => x"C0C0BFF9A4B0A492",
-12324 => x"C0C0BFF9A4B0A499",
-12323 => x"C0C0BFF9A4B0A4B0",
-12322 => x"C0C0BFF9A4B0A4A4",
-12321 => x"C0C0BFF9A4B0A4F9",
-12320 => x"C0C0BFF9A4B0A4C0",
-12319 => x"C0C0BFF9A4B0F990",
-12318 => x"C0C0BFF9A4B0F980",
-12317 => x"C0C0BFF9A4B0F9F8",
-12316 => x"C0C0BFF9A4B0F982",
-12315 => x"C0C0BFF9A4B0F992",
-12314 => x"C0C0BFF9A4B0F999",
-12313 => x"C0C0BFF9A4B0F9B0",
-12312 => x"C0C0BFF9A4B0F9A4",
-12311 => x"C0C0BFF9A4B0F9F9",
-12310 => x"C0C0BFF9A4B0F9C0",
-12309 => x"C0C0BFF9A4B0C090",
-12308 => x"C0C0BFF9A4B0C080",
-12307 => x"C0C0BFF9A4B0C0F8",
-12306 => x"C0C0BFF9A4B0C082",
-12305 => x"C0C0BFF9A4B0C092",
-12304 => x"C0C0BFF9A4B0C099",
-12303 => x"C0C0BFF9A4B0C0B0",
-12302 => x"C0C0BFF9A4B0C0A4",
-12301 => x"C0C0BFF9A4B0C0F9",
-12300 => x"C0C0BFF9A4B0C0C0",
-12299 => x"C0C0BFF9A4A49090",
-12298 => x"C0C0BFF9A4A49080",
-12297 => x"C0C0BFF9A4A490F8",
-12296 => x"C0C0BFF9A4A49082",
-12295 => x"C0C0BFF9A4A49092",
-12294 => x"C0C0BFF9A4A49099",
-12293 => x"C0C0BFF9A4A490B0",
-12292 => x"C0C0BFF9A4A490A4",
-12291 => x"C0C0BFF9A4A490F9",
-12290 => x"C0C0BFF9A4A490C0",
-12289 => x"C0C0BFF9A4A48090",
-12288 => x"C0C0BFF9A4A48080",
-12287 => x"C0C0BFF9A4A480F8",
-12286 => x"C0C0BFF9A4A48082",
-12285 => x"C0C0BFF9A4A48092",
-12284 => x"C0C0BFF9A4A48099",
-12283 => x"C0C0BFF9A4A480B0",
-12282 => x"C0C0BFF9A4A480A4",
-12281 => x"C0C0BFF9A4A480F9",
-12280 => x"C0C0BFF9A4A480C0",
-12279 => x"C0C0BFF9A4A4F890",
-12278 => x"C0C0BFF9A4A4F880",
-12277 => x"C0C0BFF9A4A4F8F8",
-12276 => x"C0C0BFF9A4A4F882",
-12275 => x"C0C0BFF9A4A4F892",
-12274 => x"C0C0BFF9A4A4F899",
-12273 => x"C0C0BFF9A4A4F8B0",
-12272 => x"C0C0BFF9A4A4F8A4",
-12271 => x"C0C0BFF9A4A4F8F9",
-12270 => x"C0C0BFF9A4A4F8C0",
-12269 => x"C0C0BFF9A4A48290",
-12268 => x"C0C0BFF9A4A48280",
-12267 => x"C0C0BFF9A4A482F8",
-12266 => x"C0C0BFF9A4A48282",
-12265 => x"C0C0BFF9A4A48292",
-12264 => x"C0C0BFF9A4A48299",
-12263 => x"C0C0BFF9A4A482B0",
-12262 => x"C0C0BFF9A4A482A4",
-12261 => x"C0C0BFF9A4A482F9",
-12260 => x"C0C0BFF9A4A482C0",
-12259 => x"C0C0BFF9A4A49290",
-12258 => x"C0C0BFF9A4A49280",
-12257 => x"C0C0BFF9A4A492F8",
-12256 => x"C0C0BFF9A4A49282",
-12255 => x"C0C0BFF9A4A49292",
-12254 => x"C0C0BFF9A4A49299",
-12253 => x"C0C0BFF9A4A492B0",
-12252 => x"C0C0BFF9A4A492A4",
-12251 => x"C0C0BFF9A4A492F9",
-12250 => x"C0C0BFF9A4A492C0",
-12249 => x"C0C0BFF9A4A49990",
-12248 => x"C0C0BFF9A4A49980",
-12247 => x"C0C0BFF9A4A499F8",
-12246 => x"C0C0BFF9A4A49982",
-12245 => x"C0C0BFF9A4A49992",
-12244 => x"C0C0BFF9A4A49999",
-12243 => x"C0C0BFF9A4A499B0",
-12242 => x"C0C0BFF9A4A499A4",
-12241 => x"C0C0BFF9A4A499F9",
-12240 => x"C0C0BFF9A4A499C0",
-12239 => x"C0C0BFF9A4A4B090",
-12238 => x"C0C0BFF9A4A4B080",
-12237 => x"C0C0BFF9A4A4B0F8",
-12236 => x"C0C0BFF9A4A4B082",
-12235 => x"C0C0BFF9A4A4B092",
-12234 => x"C0C0BFF9A4A4B099",
-12233 => x"C0C0BFF9A4A4B0B0",
-12232 => x"C0C0BFF9A4A4B0A4",
-12231 => x"C0C0BFF9A4A4B0F9",
-12230 => x"C0C0BFF9A4A4B0C0",
-12229 => x"C0C0BFF9A4A4A490",
-12228 => x"C0C0BFF9A4A4A480",
-12227 => x"C0C0BFF9A4A4A4F8",
-12226 => x"C0C0BFF9A4A4A482",
-12225 => x"C0C0BFF9A4A4A492",
-12224 => x"C0C0BFF9A4A4A499",
-12223 => x"C0C0BFF9A4A4A4B0",
-12222 => x"C0C0BFF9A4A4A4A4",
-12221 => x"C0C0BFF9A4A4A4F9",
-12220 => x"C0C0BFF9A4A4A4C0",
-12219 => x"C0C0BFF9A4A4F990",
-12218 => x"C0C0BFF9A4A4F980",
-12217 => x"C0C0BFF9A4A4F9F8",
-12216 => x"C0C0BFF9A4A4F982",
-12215 => x"C0C0BFF9A4A4F992",
-12214 => x"C0C0BFF9A4A4F999",
-12213 => x"C0C0BFF9A4A4F9B0",
-12212 => x"C0C0BFF9A4A4F9A4",
-12211 => x"C0C0BFF9A4A4F9F9",
-12210 => x"C0C0BFF9A4A4F9C0",
-12209 => x"C0C0BFF9A4A4C090",
-12208 => x"C0C0BFF9A4A4C080",
-12207 => x"C0C0BFF9A4A4C0F8",
-12206 => x"C0C0BFF9A4A4C082",
-12205 => x"C0C0BFF9A4A4C092",
-12204 => x"C0C0BFF9A4A4C099",
-12203 => x"C0C0BFF9A4A4C0B0",
-12202 => x"C0C0BFF9A4A4C0A4",
-12201 => x"C0C0BFF9A4A4C0F9",
-12200 => x"C0C0BFF9A4A4C0C0",
-12199 => x"C0C0BFF9A4F99090",
-12198 => x"C0C0BFF9A4F99080",
-12197 => x"C0C0BFF9A4F990F8",
-12196 => x"C0C0BFF9A4F99082",
-12195 => x"C0C0BFF9A4F99092",
-12194 => x"C0C0BFF9A4F99099",
-12193 => x"C0C0BFF9A4F990B0",
-12192 => x"C0C0BFF9A4F990A4",
-12191 => x"C0C0BFF9A4F990F9",
-12190 => x"C0C0BFF9A4F990C0",
-12189 => x"C0C0BFF9A4F98090",
-12188 => x"C0C0BFF9A4F98080",
-12187 => x"C0C0BFF9A4F980F8",
-12186 => x"C0C0BFF9A4F98082",
-12185 => x"C0C0BFF9A4F98092",
-12184 => x"C0C0BFF9A4F98099",
-12183 => x"C0C0BFF9A4F980B0",
-12182 => x"C0C0BFF9A4F980A4",
-12181 => x"C0C0BFF9A4F980F9",
-12180 => x"C0C0BFF9A4F980C0",
-12179 => x"C0C0BFF9A4F9F890",
-12178 => x"C0C0BFF9A4F9F880",
-12177 => x"C0C0BFF9A4F9F8F8",
-12176 => x"C0C0BFF9A4F9F882",
-12175 => x"C0C0BFF9A4F9F892",
-12174 => x"C0C0BFF9A4F9F899",
-12173 => x"C0C0BFF9A4F9F8B0",
-12172 => x"C0C0BFF9A4F9F8A4",
-12171 => x"C0C0BFF9A4F9F8F9",
-12170 => x"C0C0BFF9A4F9F8C0",
-12169 => x"C0C0BFF9A4F98290",
-12168 => x"C0C0BFF9A4F98280",
-12167 => x"C0C0BFF9A4F982F8",
-12166 => x"C0C0BFF9A4F98282",
-12165 => x"C0C0BFF9A4F98292",
-12164 => x"C0C0BFF9A4F98299",
-12163 => x"C0C0BFF9A4F982B0",
-12162 => x"C0C0BFF9A4F982A4",
-12161 => x"C0C0BFF9A4F982F9",
-12160 => x"C0C0BFF9A4F982C0",
-12159 => x"C0C0BFF9A4F99290",
-12158 => x"C0C0BFF9A4F99280",
-12157 => x"C0C0BFF9A4F992F8",
-12156 => x"C0C0BFF9A4F99282",
-12155 => x"C0C0BFF9A4F99292",
-12154 => x"C0C0BFF9A4F99299",
-12153 => x"C0C0BFF9A4F992B0",
-12152 => x"C0C0BFF9A4F992A4",
-12151 => x"C0C0BFF9A4F992F9",
-12150 => x"C0C0BFF9A4F992C0",
-12149 => x"C0C0BFF9A4F99990",
-12148 => x"C0C0BFF9A4F99980",
-12147 => x"C0C0BFF9A4F999F8",
-12146 => x"C0C0BFF9A4F99982",
-12145 => x"C0C0BFF9A4F99992",
-12144 => x"C0C0BFF9A4F99999",
-12143 => x"C0C0BFF9A4F999B0",
-12142 => x"C0C0BFF9A4F999A4",
-12141 => x"C0C0BFF9A4F999F9",
-12140 => x"C0C0BFF9A4F999C0",
-12139 => x"C0C0BFF9A4F9B090",
-12138 => x"C0C0BFF9A4F9B080",
-12137 => x"C0C0BFF9A4F9B0F8",
-12136 => x"C0C0BFF9A4F9B082",
-12135 => x"C0C0BFF9A4F9B092",
-12134 => x"C0C0BFF9A4F9B099",
-12133 => x"C0C0BFF9A4F9B0B0",
-12132 => x"C0C0BFF9A4F9B0A4",
-12131 => x"C0C0BFF9A4F9B0F9",
-12130 => x"C0C0BFF9A4F9B0C0",
-12129 => x"C0C0BFF9A4F9A490",
-12128 => x"C0C0BFF9A4F9A480",
-12127 => x"C0C0BFF9A4F9A4F8",
-12126 => x"C0C0BFF9A4F9A482",
-12125 => x"C0C0BFF9A4F9A492",
-12124 => x"C0C0BFF9A4F9A499",
-12123 => x"C0C0BFF9A4F9A4B0",
-12122 => x"C0C0BFF9A4F9A4A4",
-12121 => x"C0C0BFF9A4F9A4F9",
-12120 => x"C0C0BFF9A4F9A4C0",
-12119 => x"C0C0BFF9A4F9F990",
-12118 => x"C0C0BFF9A4F9F980",
-12117 => x"C0C0BFF9A4F9F9F8",
-12116 => x"C0C0BFF9A4F9F982",
-12115 => x"C0C0BFF9A4F9F992",
-12114 => x"C0C0BFF9A4F9F999",
-12113 => x"C0C0BFF9A4F9F9B0",
-12112 => x"C0C0BFF9A4F9F9A4",
-12111 => x"C0C0BFF9A4F9F9F9",
-12110 => x"C0C0BFF9A4F9F9C0",
-12109 => x"C0C0BFF9A4F9C090",
-12108 => x"C0C0BFF9A4F9C080",
-12107 => x"C0C0BFF9A4F9C0F8",
-12106 => x"C0C0BFF9A4F9C082",
-12105 => x"C0C0BFF9A4F9C092",
-12104 => x"C0C0BFF9A4F9C099",
-12103 => x"C0C0BFF9A4F9C0B0",
-12102 => x"C0C0BFF9A4F9C0A4",
-12101 => x"C0C0BFF9A4F9C0F9",
-12100 => x"C0C0BFF9A4F9C0C0",
-12099 => x"C0C0BFF9A4C09090",
-12098 => x"C0C0BFF9A4C09080",
-12097 => x"C0C0BFF9A4C090F8",
-12096 => x"C0C0BFF9A4C09082",
-12095 => x"C0C0BFF9A4C09092",
-12094 => x"C0C0BFF9A4C09099",
-12093 => x"C0C0BFF9A4C090B0",
-12092 => x"C0C0BFF9A4C090A4",
-12091 => x"C0C0BFF9A4C090F9",
-12090 => x"C0C0BFF9A4C090C0",
-12089 => x"C0C0BFF9A4C08090",
-12088 => x"C0C0BFF9A4C08080",
-12087 => x"C0C0BFF9A4C080F8",
-12086 => x"C0C0BFF9A4C08082",
-12085 => x"C0C0BFF9A4C08092",
-12084 => x"C0C0BFF9A4C08099",
-12083 => x"C0C0BFF9A4C080B0",
-12082 => x"C0C0BFF9A4C080A4",
-12081 => x"C0C0BFF9A4C080F9",
-12080 => x"C0C0BFF9A4C080C0",
-12079 => x"C0C0BFF9A4C0F890",
-12078 => x"C0C0BFF9A4C0F880",
-12077 => x"C0C0BFF9A4C0F8F8",
-12076 => x"C0C0BFF9A4C0F882",
-12075 => x"C0C0BFF9A4C0F892",
-12074 => x"C0C0BFF9A4C0F899",
-12073 => x"C0C0BFF9A4C0F8B0",
-12072 => x"C0C0BFF9A4C0F8A4",
-12071 => x"C0C0BFF9A4C0F8F9",
-12070 => x"C0C0BFF9A4C0F8C0",
-12069 => x"C0C0BFF9A4C08290",
-12068 => x"C0C0BFF9A4C08280",
-12067 => x"C0C0BFF9A4C082F8",
-12066 => x"C0C0BFF9A4C08282",
-12065 => x"C0C0BFF9A4C08292",
-12064 => x"C0C0BFF9A4C08299",
-12063 => x"C0C0BFF9A4C082B0",
-12062 => x"C0C0BFF9A4C082A4",
-12061 => x"C0C0BFF9A4C082F9",
-12060 => x"C0C0BFF9A4C082C0",
-12059 => x"C0C0BFF9A4C09290",
-12058 => x"C0C0BFF9A4C09280",
-12057 => x"C0C0BFF9A4C092F8",
-12056 => x"C0C0BFF9A4C09282",
-12055 => x"C0C0BFF9A4C09292",
-12054 => x"C0C0BFF9A4C09299",
-12053 => x"C0C0BFF9A4C092B0",
-12052 => x"C0C0BFF9A4C092A4",
-12051 => x"C0C0BFF9A4C092F9",
-12050 => x"C0C0BFF9A4C092C0",
-12049 => x"C0C0BFF9A4C09990",
-12048 => x"C0C0BFF9A4C09980",
-12047 => x"C0C0BFF9A4C099F8",
-12046 => x"C0C0BFF9A4C09982",
-12045 => x"C0C0BFF9A4C09992",
-12044 => x"C0C0BFF9A4C09999",
-12043 => x"C0C0BFF9A4C099B0",
-12042 => x"C0C0BFF9A4C099A4",
-12041 => x"C0C0BFF9A4C099F9",
-12040 => x"C0C0BFF9A4C099C0",
-12039 => x"C0C0BFF9A4C0B090",
-12038 => x"C0C0BFF9A4C0B080",
-12037 => x"C0C0BFF9A4C0B0F8",
-12036 => x"C0C0BFF9A4C0B082",
-12035 => x"C0C0BFF9A4C0B092",
-12034 => x"C0C0BFF9A4C0B099",
-12033 => x"C0C0BFF9A4C0B0B0",
-12032 => x"C0C0BFF9A4C0B0A4",
-12031 => x"C0C0BFF9A4C0B0F9",
-12030 => x"C0C0BFF9A4C0B0C0",
-12029 => x"C0C0BFF9A4C0A490",
-12028 => x"C0C0BFF9A4C0A480",
-12027 => x"C0C0BFF9A4C0A4F8",
-12026 => x"C0C0BFF9A4C0A482",
-12025 => x"C0C0BFF9A4C0A492",
-12024 => x"C0C0BFF9A4C0A499",
-12023 => x"C0C0BFF9A4C0A4B0",
-12022 => x"C0C0BFF9A4C0A4A4",
-12021 => x"C0C0BFF9A4C0A4F9",
-12020 => x"C0C0BFF9A4C0A4C0",
-12019 => x"C0C0BFF9A4C0F990",
-12018 => x"C0C0BFF9A4C0F980",
-12017 => x"C0C0BFF9A4C0F9F8",
-12016 => x"C0C0BFF9A4C0F982",
-12015 => x"C0C0BFF9A4C0F992",
-12014 => x"C0C0BFF9A4C0F999",
-12013 => x"C0C0BFF9A4C0F9B0",
-12012 => x"C0C0BFF9A4C0F9A4",
-12011 => x"C0C0BFF9A4C0F9F9",
-12010 => x"C0C0BFF9A4C0F9C0",
-12009 => x"C0C0BFF9A4C0C090",
-12008 => x"C0C0BFF9A4C0C080",
-12007 => x"C0C0BFF9A4C0C0F8",
-12006 => x"C0C0BFF9A4C0C082",
-12005 => x"C0C0BFF9A4C0C092",
-12004 => x"C0C0BFF9A4C0C099",
-12003 => x"C0C0BFF9A4C0C0B0",
-12002 => x"C0C0BFF9A4C0C0A4",
-12001 => x"C0C0BFF9A4C0C0F9",
-12000 => x"C0C0BFF9A4C0C0C0",
-11999 => x"C0C0BFF9F9909090",
-11998 => x"C0C0BFF9F9909080",
-11997 => x"C0C0BFF9F99090F8",
-11996 => x"C0C0BFF9F9909082",
-11995 => x"C0C0BFF9F9909092",
-11994 => x"C0C0BFF9F9909099",
-11993 => x"C0C0BFF9F99090B0",
-11992 => x"C0C0BFF9F99090A4",
-11991 => x"C0C0BFF9F99090F9",
-11990 => x"C0C0BFF9F99090C0",
-11989 => x"C0C0BFF9F9908090",
-11988 => x"C0C0BFF9F9908080",
-11987 => x"C0C0BFF9F99080F8",
-11986 => x"C0C0BFF9F9908082",
-11985 => x"C0C0BFF9F9908092",
-11984 => x"C0C0BFF9F9908099",
-11983 => x"C0C0BFF9F99080B0",
-11982 => x"C0C0BFF9F99080A4",
-11981 => x"C0C0BFF9F99080F9",
-11980 => x"C0C0BFF9F99080C0",
-11979 => x"C0C0BFF9F990F890",
-11978 => x"C0C0BFF9F990F880",
-11977 => x"C0C0BFF9F990F8F8",
-11976 => x"C0C0BFF9F990F882",
-11975 => x"C0C0BFF9F990F892",
-11974 => x"C0C0BFF9F990F899",
-11973 => x"C0C0BFF9F990F8B0",
-11972 => x"C0C0BFF9F990F8A4",
-11971 => x"C0C0BFF9F990F8F9",
-11970 => x"C0C0BFF9F990F8C0",
-11969 => x"C0C0BFF9F9908290",
-11968 => x"C0C0BFF9F9908280",
-11967 => x"C0C0BFF9F99082F8",
-11966 => x"C0C0BFF9F9908282",
-11965 => x"C0C0BFF9F9908292",
-11964 => x"C0C0BFF9F9908299",
-11963 => x"C0C0BFF9F99082B0",
-11962 => x"C0C0BFF9F99082A4",
-11961 => x"C0C0BFF9F99082F9",
-11960 => x"C0C0BFF9F99082C0",
-11959 => x"C0C0BFF9F9909290",
-11958 => x"C0C0BFF9F9909280",
-11957 => x"C0C0BFF9F99092F8",
-11956 => x"C0C0BFF9F9909282",
-11955 => x"C0C0BFF9F9909292",
-11954 => x"C0C0BFF9F9909299",
-11953 => x"C0C0BFF9F99092B0",
-11952 => x"C0C0BFF9F99092A4",
-11951 => x"C0C0BFF9F99092F9",
-11950 => x"C0C0BFF9F99092C0",
-11949 => x"C0C0BFF9F9909990",
-11948 => x"C0C0BFF9F9909980",
-11947 => x"C0C0BFF9F99099F8",
-11946 => x"C0C0BFF9F9909982",
-11945 => x"C0C0BFF9F9909992",
-11944 => x"C0C0BFF9F9909999",
-11943 => x"C0C0BFF9F99099B0",
-11942 => x"C0C0BFF9F99099A4",
-11941 => x"C0C0BFF9F99099F9",
-11940 => x"C0C0BFF9F99099C0",
-11939 => x"C0C0BFF9F990B090",
-11938 => x"C0C0BFF9F990B080",
-11937 => x"C0C0BFF9F990B0F8",
-11936 => x"C0C0BFF9F990B082",
-11935 => x"C0C0BFF9F990B092",
-11934 => x"C0C0BFF9F990B099",
-11933 => x"C0C0BFF9F990B0B0",
-11932 => x"C0C0BFF9F990B0A4",
-11931 => x"C0C0BFF9F990B0F9",
-11930 => x"C0C0BFF9F990B0C0",
-11929 => x"C0C0BFF9F990A490",
-11928 => x"C0C0BFF9F990A480",
-11927 => x"C0C0BFF9F990A4F8",
-11926 => x"C0C0BFF9F990A482",
-11925 => x"C0C0BFF9F990A492",
-11924 => x"C0C0BFF9F990A499",
-11923 => x"C0C0BFF9F990A4B0",
-11922 => x"C0C0BFF9F990A4A4",
-11921 => x"C0C0BFF9F990A4F9",
-11920 => x"C0C0BFF9F990A4C0",
-11919 => x"C0C0BFF9F990F990",
-11918 => x"C0C0BFF9F990F980",
-11917 => x"C0C0BFF9F990F9F8",
-11916 => x"C0C0BFF9F990F982",
-11915 => x"C0C0BFF9F990F992",
-11914 => x"C0C0BFF9F990F999",
-11913 => x"C0C0BFF9F990F9B0",
-11912 => x"C0C0BFF9F990F9A4",
-11911 => x"C0C0BFF9F990F9F9",
-11910 => x"C0C0BFF9F990F9C0",
-11909 => x"C0C0BFF9F990C090",
-11908 => x"C0C0BFF9F990C080",
-11907 => x"C0C0BFF9F990C0F8",
-11906 => x"C0C0BFF9F990C082",
-11905 => x"C0C0BFF9F990C092",
-11904 => x"C0C0BFF9F990C099",
-11903 => x"C0C0BFF9F990C0B0",
-11902 => x"C0C0BFF9F990C0A4",
-11901 => x"C0C0BFF9F990C0F9",
-11900 => x"C0C0BFF9F990C0C0",
-11899 => x"C0C0BFF9F9809090",
-11898 => x"C0C0BFF9F9809080",
-11897 => x"C0C0BFF9F98090F8",
-11896 => x"C0C0BFF9F9809082",
-11895 => x"C0C0BFF9F9809092",
-11894 => x"C0C0BFF9F9809099",
-11893 => x"C0C0BFF9F98090B0",
-11892 => x"C0C0BFF9F98090A4",
-11891 => x"C0C0BFF9F98090F9",
-11890 => x"C0C0BFF9F98090C0",
-11889 => x"C0C0BFF9F9808090",
-11888 => x"C0C0BFF9F9808080",
-11887 => x"C0C0BFF9F98080F8",
-11886 => x"C0C0BFF9F9808082",
-11885 => x"C0C0BFF9F9808092",
-11884 => x"C0C0BFF9F9808099",
-11883 => x"C0C0BFF9F98080B0",
-11882 => x"C0C0BFF9F98080A4",
-11881 => x"C0C0BFF9F98080F9",
-11880 => x"C0C0BFF9F98080C0",
-11879 => x"C0C0BFF9F980F890",
-11878 => x"C0C0BFF9F980F880",
-11877 => x"C0C0BFF9F980F8F8",
-11876 => x"C0C0BFF9F980F882",
-11875 => x"C0C0BFF9F980F892",
-11874 => x"C0C0BFF9F980F899",
-11873 => x"C0C0BFF9F980F8B0",
-11872 => x"C0C0BFF9F980F8A4",
-11871 => x"C0C0BFF9F980F8F9",
-11870 => x"C0C0BFF9F980F8C0",
-11869 => x"C0C0BFF9F9808290",
-11868 => x"C0C0BFF9F9808280",
-11867 => x"C0C0BFF9F98082F8",
-11866 => x"C0C0BFF9F9808282",
-11865 => x"C0C0BFF9F9808292",
-11864 => x"C0C0BFF9F9808299",
-11863 => x"C0C0BFF9F98082B0",
-11862 => x"C0C0BFF9F98082A4",
-11861 => x"C0C0BFF9F98082F9",
-11860 => x"C0C0BFF9F98082C0",
-11859 => x"C0C0BFF9F9809290",
-11858 => x"C0C0BFF9F9809280",
-11857 => x"C0C0BFF9F98092F8",
-11856 => x"C0C0BFF9F9809282",
-11855 => x"C0C0BFF9F9809292",
-11854 => x"C0C0BFF9F9809299",
-11853 => x"C0C0BFF9F98092B0",
-11852 => x"C0C0BFF9F98092A4",
-11851 => x"C0C0BFF9F98092F9",
-11850 => x"C0C0BFF9F98092C0",
-11849 => x"C0C0BFF9F9809990",
-11848 => x"C0C0BFF9F9809980",
-11847 => x"C0C0BFF9F98099F8",
-11846 => x"C0C0BFF9F9809982",
-11845 => x"C0C0BFF9F9809992",
-11844 => x"C0C0BFF9F9809999",
-11843 => x"C0C0BFF9F98099B0",
-11842 => x"C0C0BFF9F98099A4",
-11841 => x"C0C0BFF9F98099F9",
-11840 => x"C0C0BFF9F98099C0",
-11839 => x"C0C0BFF9F980B090",
-11838 => x"C0C0BFF9F980B080",
-11837 => x"C0C0BFF9F980B0F8",
-11836 => x"C0C0BFF9F980B082",
-11835 => x"C0C0BFF9F980B092",
-11834 => x"C0C0BFF9F980B099",
-11833 => x"C0C0BFF9F980B0B0",
-11832 => x"C0C0BFF9F980B0A4",
-11831 => x"C0C0BFF9F980B0F9",
-11830 => x"C0C0BFF9F980B0C0",
-11829 => x"C0C0BFF9F980A490",
-11828 => x"C0C0BFF9F980A480",
-11827 => x"C0C0BFF9F980A4F8",
-11826 => x"C0C0BFF9F980A482",
-11825 => x"C0C0BFF9F980A492",
-11824 => x"C0C0BFF9F980A499",
-11823 => x"C0C0BFF9F980A4B0",
-11822 => x"C0C0BFF9F980A4A4",
-11821 => x"C0C0BFF9F980A4F9",
-11820 => x"C0C0BFF9F980A4C0",
-11819 => x"C0C0BFF9F980F990",
-11818 => x"C0C0BFF9F980F980",
-11817 => x"C0C0BFF9F980F9F8",
-11816 => x"C0C0BFF9F980F982",
-11815 => x"C0C0BFF9F980F992",
-11814 => x"C0C0BFF9F980F999",
-11813 => x"C0C0BFF9F980F9B0",
-11812 => x"C0C0BFF9F980F9A4",
-11811 => x"C0C0BFF9F980F9F9",
-11810 => x"C0C0BFF9F980F9C0",
-11809 => x"C0C0BFF9F980C090",
-11808 => x"C0C0BFF9F980C080",
-11807 => x"C0C0BFF9F980C0F8",
-11806 => x"C0C0BFF9F980C082",
-11805 => x"C0C0BFF9F980C092",
-11804 => x"C0C0BFF9F980C099",
-11803 => x"C0C0BFF9F980C0B0",
-11802 => x"C0C0BFF9F980C0A4",
-11801 => x"C0C0BFF9F980C0F9",
-11800 => x"C0C0BFF9F980C0C0",
-11799 => x"C0C0BFF9F9F89090",
-11798 => x"C0C0BFF9F9F89080",
-11797 => x"C0C0BFF9F9F890F8",
-11796 => x"C0C0BFF9F9F89082",
-11795 => x"C0C0BFF9F9F89092",
-11794 => x"C0C0BFF9F9F89099",
-11793 => x"C0C0BFF9F9F890B0",
-11792 => x"C0C0BFF9F9F890A4",
-11791 => x"C0C0BFF9F9F890F9",
-11790 => x"C0C0BFF9F9F890C0",
-11789 => x"C0C0BFF9F9F88090",
-11788 => x"C0C0BFF9F9F88080",
-11787 => x"C0C0BFF9F9F880F8",
-11786 => x"C0C0BFF9F9F88082",
-11785 => x"C0C0BFF9F9F88092",
-11784 => x"C0C0BFF9F9F88099",
-11783 => x"C0C0BFF9F9F880B0",
-11782 => x"C0C0BFF9F9F880A4",
-11781 => x"C0C0BFF9F9F880F9",
-11780 => x"C0C0BFF9F9F880C0",
-11779 => x"C0C0BFF9F9F8F890",
-11778 => x"C0C0BFF9F9F8F880",
-11777 => x"C0C0BFF9F9F8F8F8",
-11776 => x"C0C0BFF9F9F8F882",
-11775 => x"C0C0BFF9F9F8F892",
-11774 => x"C0C0BFF9F9F8F899",
-11773 => x"C0C0BFF9F9F8F8B0",
-11772 => x"C0C0BFF9F9F8F8A4",
-11771 => x"C0C0BFF9F9F8F8F9",
-11770 => x"C0C0BFF9F9F8F8C0",
-11769 => x"C0C0BFF9F9F88290",
-11768 => x"C0C0BFF9F9F88280",
-11767 => x"C0C0BFF9F9F882F8",
-11766 => x"C0C0BFF9F9F88282",
-11765 => x"C0C0BFF9F9F88292",
-11764 => x"C0C0BFF9F9F88299",
-11763 => x"C0C0BFF9F9F882B0",
-11762 => x"C0C0BFF9F9F882A4",
-11761 => x"C0C0BFF9F9F882F9",
-11760 => x"C0C0BFF9F9F882C0",
-11759 => x"C0C0BFF9F9F89290",
-11758 => x"C0C0BFF9F9F89280",
-11757 => x"C0C0BFF9F9F892F8",
-11756 => x"C0C0BFF9F9F89282",
-11755 => x"C0C0BFF9F9F89292",
-11754 => x"C0C0BFF9F9F89299",
-11753 => x"C0C0BFF9F9F892B0",
-11752 => x"C0C0BFF9F9F892A4",
-11751 => x"C0C0BFF9F9F892F9",
-11750 => x"C0C0BFF9F9F892C0",
-11749 => x"C0C0BFF9F9F89990",
-11748 => x"C0C0BFF9F9F89980",
-11747 => x"C0C0BFF9F9F899F8",
-11746 => x"C0C0BFF9F9F89982",
-11745 => x"C0C0BFF9F9F89992",
-11744 => x"C0C0BFF9F9F89999",
-11743 => x"C0C0BFF9F9F899B0",
-11742 => x"C0C0BFF9F9F899A4",
-11741 => x"C0C0BFF9F9F899F9",
-11740 => x"C0C0BFF9F9F899C0",
-11739 => x"C0C0BFF9F9F8B090",
-11738 => x"C0C0BFF9F9F8B080",
-11737 => x"C0C0BFF9F9F8B0F8",
-11736 => x"C0C0BFF9F9F8B082",
-11735 => x"C0C0BFF9F9F8B092",
-11734 => x"C0C0BFF9F9F8B099",
-11733 => x"C0C0BFF9F9F8B0B0",
-11732 => x"C0C0BFF9F9F8B0A4",
-11731 => x"C0C0BFF9F9F8B0F9",
-11730 => x"C0C0BFF9F9F8B0C0",
-11729 => x"C0C0BFF9F9F8A490",
-11728 => x"C0C0BFF9F9F8A480",
-11727 => x"C0C0BFF9F9F8A4F8",
-11726 => x"C0C0BFF9F9F8A482",
-11725 => x"C0C0BFF9F9F8A492",
-11724 => x"C0C0BFF9F9F8A499",
-11723 => x"C0C0BFF9F9F8A4B0",
-11722 => x"C0C0BFF9F9F8A4A4",
-11721 => x"C0C0BFF9F9F8A4F9",
-11720 => x"C0C0BFF9F9F8A4C0",
-11719 => x"C0C0BFF9F9F8F990",
-11718 => x"C0C0BFF9F9F8F980",
-11717 => x"C0C0BFF9F9F8F9F8",
-11716 => x"C0C0BFF9F9F8F982",
-11715 => x"C0C0BFF9F9F8F992",
-11714 => x"C0C0BFF9F9F8F999",
-11713 => x"C0C0BFF9F9F8F9B0",
-11712 => x"C0C0BFF9F9F8F9A4",
-11711 => x"C0C0BFF9F9F8F9F9",
-11710 => x"C0C0BFF9F9F8F9C0",
-11709 => x"C0C0BFF9F9F8C090",
-11708 => x"C0C0BFF9F9F8C080",
-11707 => x"C0C0BFF9F9F8C0F8",
-11706 => x"C0C0BFF9F9F8C082",
-11705 => x"C0C0BFF9F9F8C092",
-11704 => x"C0C0BFF9F9F8C099",
-11703 => x"C0C0BFF9F9F8C0B0",
-11702 => x"C0C0BFF9F9F8C0A4",
-11701 => x"C0C0BFF9F9F8C0F9",
-11700 => x"C0C0BFF9F9F8C0C0",
-11699 => x"C0C0BFF9F9829090",
-11698 => x"C0C0BFF9F9829080",
-11697 => x"C0C0BFF9F98290F8",
-11696 => x"C0C0BFF9F9829082",
-11695 => x"C0C0BFF9F9829092",
-11694 => x"C0C0BFF9F9829099",
-11693 => x"C0C0BFF9F98290B0",
-11692 => x"C0C0BFF9F98290A4",
-11691 => x"C0C0BFF9F98290F9",
-11690 => x"C0C0BFF9F98290C0",
-11689 => x"C0C0BFF9F9828090",
-11688 => x"C0C0BFF9F9828080",
-11687 => x"C0C0BFF9F98280F8",
-11686 => x"C0C0BFF9F9828082",
-11685 => x"C0C0BFF9F9828092",
-11684 => x"C0C0BFF9F9828099",
-11683 => x"C0C0BFF9F98280B0",
-11682 => x"C0C0BFF9F98280A4",
-11681 => x"C0C0BFF9F98280F9",
-11680 => x"C0C0BFF9F98280C0",
-11679 => x"C0C0BFF9F982F890",
-11678 => x"C0C0BFF9F982F880",
-11677 => x"C0C0BFF9F982F8F8",
-11676 => x"C0C0BFF9F982F882",
-11675 => x"C0C0BFF9F982F892",
-11674 => x"C0C0BFF9F982F899",
-11673 => x"C0C0BFF9F982F8B0",
-11672 => x"C0C0BFF9F982F8A4",
-11671 => x"C0C0BFF9F982F8F9",
-11670 => x"C0C0BFF9F982F8C0",
-11669 => x"C0C0BFF9F9828290",
-11668 => x"C0C0BFF9F9828280",
-11667 => x"C0C0BFF9F98282F8",
-11666 => x"C0C0BFF9F9828282",
-11665 => x"C0C0BFF9F9828292",
-11664 => x"C0C0BFF9F9828299",
-11663 => x"C0C0BFF9F98282B0",
-11662 => x"C0C0BFF9F98282A4",
-11661 => x"C0C0BFF9F98282F9",
-11660 => x"C0C0BFF9F98282C0",
-11659 => x"C0C0BFF9F9829290",
-11658 => x"C0C0BFF9F9829280",
-11657 => x"C0C0BFF9F98292F8",
-11656 => x"C0C0BFF9F9829282",
-11655 => x"C0C0BFF9F9829292",
-11654 => x"C0C0BFF9F9829299",
-11653 => x"C0C0BFF9F98292B0",
-11652 => x"C0C0BFF9F98292A4",
-11651 => x"C0C0BFF9F98292F9",
-11650 => x"C0C0BFF9F98292C0",
-11649 => x"C0C0BFF9F9829990",
-11648 => x"C0C0BFF9F9829980",
-11647 => x"C0C0BFF9F98299F8",
-11646 => x"C0C0BFF9F9829982",
-11645 => x"C0C0BFF9F9829992",
-11644 => x"C0C0BFF9F9829999",
-11643 => x"C0C0BFF9F98299B0",
-11642 => x"C0C0BFF9F98299A4",
-11641 => x"C0C0BFF9F98299F9",
-11640 => x"C0C0BFF9F98299C0",
-11639 => x"C0C0BFF9F982B090",
-11638 => x"C0C0BFF9F982B080",
-11637 => x"C0C0BFF9F982B0F8",
-11636 => x"C0C0BFF9F982B082",
-11635 => x"C0C0BFF9F982B092",
-11634 => x"C0C0BFF9F982B099",
-11633 => x"C0C0BFF9F982B0B0",
-11632 => x"C0C0BFF9F982B0A4",
-11631 => x"C0C0BFF9F982B0F9",
-11630 => x"C0C0BFF9F982B0C0",
-11629 => x"C0C0BFF9F982A490",
-11628 => x"C0C0BFF9F982A480",
-11627 => x"C0C0BFF9F982A4F8",
-11626 => x"C0C0BFF9F982A482",
-11625 => x"C0C0BFF9F982A492",
-11624 => x"C0C0BFF9F982A499",
-11623 => x"C0C0BFF9F982A4B0",
-11622 => x"C0C0BFF9F982A4A4",
-11621 => x"C0C0BFF9F982A4F9",
-11620 => x"C0C0BFF9F982A4C0",
-11619 => x"C0C0BFF9F982F990",
-11618 => x"C0C0BFF9F982F980",
-11617 => x"C0C0BFF9F982F9F8",
-11616 => x"C0C0BFF9F982F982",
-11615 => x"C0C0BFF9F982F992",
-11614 => x"C0C0BFF9F982F999",
-11613 => x"C0C0BFF9F982F9B0",
-11612 => x"C0C0BFF9F982F9A4",
-11611 => x"C0C0BFF9F982F9F9",
-11610 => x"C0C0BFF9F982F9C0",
-11609 => x"C0C0BFF9F982C090",
-11608 => x"C0C0BFF9F982C080",
-11607 => x"C0C0BFF9F982C0F8",
-11606 => x"C0C0BFF9F982C082",
-11605 => x"C0C0BFF9F982C092",
-11604 => x"C0C0BFF9F982C099",
-11603 => x"C0C0BFF9F982C0B0",
-11602 => x"C0C0BFF9F982C0A4",
-11601 => x"C0C0BFF9F982C0F9",
-11600 => x"C0C0BFF9F982C0C0",
-11599 => x"C0C0BFF9F9929090",
-11598 => x"C0C0BFF9F9929080",
-11597 => x"C0C0BFF9F99290F8",
-11596 => x"C0C0BFF9F9929082",
-11595 => x"C0C0BFF9F9929092",
-11594 => x"C0C0BFF9F9929099",
-11593 => x"C0C0BFF9F99290B0",
-11592 => x"C0C0BFF9F99290A4",
-11591 => x"C0C0BFF9F99290F9",
-11590 => x"C0C0BFF9F99290C0",
-11589 => x"C0C0BFF9F9928090",
-11588 => x"C0C0BFF9F9928080",
-11587 => x"C0C0BFF9F99280F8",
-11586 => x"C0C0BFF9F9928082",
-11585 => x"C0C0BFF9F9928092",
-11584 => x"C0C0BFF9F9928099",
-11583 => x"C0C0BFF9F99280B0",
-11582 => x"C0C0BFF9F99280A4",
-11581 => x"C0C0BFF9F99280F9",
-11580 => x"C0C0BFF9F99280C0",
-11579 => x"C0C0BFF9F992F890",
-11578 => x"C0C0BFF9F992F880",
-11577 => x"C0C0BFF9F992F8F8",
-11576 => x"C0C0BFF9F992F882",
-11575 => x"C0C0BFF9F992F892",
-11574 => x"C0C0BFF9F992F899",
-11573 => x"C0C0BFF9F992F8B0",
-11572 => x"C0C0BFF9F992F8A4",
-11571 => x"C0C0BFF9F992F8F9",
-11570 => x"C0C0BFF9F992F8C0",
-11569 => x"C0C0BFF9F9928290",
-11568 => x"C0C0BFF9F9928280",
-11567 => x"C0C0BFF9F99282F8",
-11566 => x"C0C0BFF9F9928282",
-11565 => x"C0C0BFF9F9928292",
-11564 => x"C0C0BFF9F9928299",
-11563 => x"C0C0BFF9F99282B0",
-11562 => x"C0C0BFF9F99282A4",
-11561 => x"C0C0BFF9F99282F9",
-11560 => x"C0C0BFF9F99282C0",
-11559 => x"C0C0BFF9F9929290",
-11558 => x"C0C0BFF9F9929280",
-11557 => x"C0C0BFF9F99292F8",
-11556 => x"C0C0BFF9F9929282",
-11555 => x"C0C0BFF9F9929292",
-11554 => x"C0C0BFF9F9929299",
-11553 => x"C0C0BFF9F99292B0",
-11552 => x"C0C0BFF9F99292A4",
-11551 => x"C0C0BFF9F99292F9",
-11550 => x"C0C0BFF9F99292C0",
-11549 => x"C0C0BFF9F9929990",
-11548 => x"C0C0BFF9F9929980",
-11547 => x"C0C0BFF9F99299F8",
-11546 => x"C0C0BFF9F9929982",
-11545 => x"C0C0BFF9F9929992",
-11544 => x"C0C0BFF9F9929999",
-11543 => x"C0C0BFF9F99299B0",
-11542 => x"C0C0BFF9F99299A4",
-11541 => x"C0C0BFF9F99299F9",
-11540 => x"C0C0BFF9F99299C0",
-11539 => x"C0C0BFF9F992B090",
-11538 => x"C0C0BFF9F992B080",
-11537 => x"C0C0BFF9F992B0F8",
-11536 => x"C0C0BFF9F992B082",
-11535 => x"C0C0BFF9F992B092",
-11534 => x"C0C0BFF9F992B099",
-11533 => x"C0C0BFF9F992B0B0",
-11532 => x"C0C0BFF9F992B0A4",
-11531 => x"C0C0BFF9F992B0F9",
-11530 => x"C0C0BFF9F992B0C0",
-11529 => x"C0C0BFF9F992A490",
-11528 => x"C0C0BFF9F992A480",
-11527 => x"C0C0BFF9F992A4F8",
-11526 => x"C0C0BFF9F992A482",
-11525 => x"C0C0BFF9F992A492",
-11524 => x"C0C0BFF9F992A499",
-11523 => x"C0C0BFF9F992A4B0",
-11522 => x"C0C0BFF9F992A4A4",
-11521 => x"C0C0BFF9F992A4F9",
-11520 => x"C0C0BFF9F992A4C0",
-11519 => x"C0C0BFF9F992F990",
-11518 => x"C0C0BFF9F992F980",
-11517 => x"C0C0BFF9F992F9F8",
-11516 => x"C0C0BFF9F992F982",
-11515 => x"C0C0BFF9F992F992",
-11514 => x"C0C0BFF9F992F999",
-11513 => x"C0C0BFF9F992F9B0",
-11512 => x"C0C0BFF9F992F9A4",
-11511 => x"C0C0BFF9F992F9F9",
-11510 => x"C0C0BFF9F992F9C0",
-11509 => x"C0C0BFF9F992C090",
-11508 => x"C0C0BFF9F992C080",
-11507 => x"C0C0BFF9F992C0F8",
-11506 => x"C0C0BFF9F992C082",
-11505 => x"C0C0BFF9F992C092",
-11504 => x"C0C0BFF9F992C099",
-11503 => x"C0C0BFF9F992C0B0",
-11502 => x"C0C0BFF9F992C0A4",
-11501 => x"C0C0BFF9F992C0F9",
-11500 => x"C0C0BFF9F992C0C0",
-11499 => x"C0C0BFF9F9999090",
-11498 => x"C0C0BFF9F9999080",
-11497 => x"C0C0BFF9F99990F8",
-11496 => x"C0C0BFF9F9999082",
-11495 => x"C0C0BFF9F9999092",
-11494 => x"C0C0BFF9F9999099",
-11493 => x"C0C0BFF9F99990B0",
-11492 => x"C0C0BFF9F99990A4",
-11491 => x"C0C0BFF9F99990F9",
-11490 => x"C0C0BFF9F99990C0",
-11489 => x"C0C0BFF9F9998090",
-11488 => x"C0C0BFF9F9998080",
-11487 => x"C0C0BFF9F99980F8",
-11486 => x"C0C0BFF9F9998082",
-11485 => x"C0C0BFF9F9998092",
-11484 => x"C0C0BFF9F9998099",
-11483 => x"C0C0BFF9F99980B0",
-11482 => x"C0C0BFF9F99980A4",
-11481 => x"C0C0BFF9F99980F9",
-11480 => x"C0C0BFF9F99980C0",
-11479 => x"C0C0BFF9F999F890",
-11478 => x"C0C0BFF9F999F880",
-11477 => x"C0C0BFF9F999F8F8",
-11476 => x"C0C0BFF9F999F882",
-11475 => x"C0C0BFF9F999F892",
-11474 => x"C0C0BFF9F999F899",
-11473 => x"C0C0BFF9F999F8B0",
-11472 => x"C0C0BFF9F999F8A4",
-11471 => x"C0C0BFF9F999F8F9",
-11470 => x"C0C0BFF9F999F8C0",
-11469 => x"C0C0BFF9F9998290",
-11468 => x"C0C0BFF9F9998280",
-11467 => x"C0C0BFF9F99982F8",
-11466 => x"C0C0BFF9F9998282",
-11465 => x"C0C0BFF9F9998292",
-11464 => x"C0C0BFF9F9998299",
-11463 => x"C0C0BFF9F99982B0",
-11462 => x"C0C0BFF9F99982A4",
-11461 => x"C0C0BFF9F99982F9",
-11460 => x"C0C0BFF9F99982C0",
-11459 => x"C0C0BFF9F9999290",
-11458 => x"C0C0BFF9F9999280",
-11457 => x"C0C0BFF9F99992F8",
-11456 => x"C0C0BFF9F9999282",
-11455 => x"C0C0BFF9F9999292",
-11454 => x"C0C0BFF9F9999299",
-11453 => x"C0C0BFF9F99992B0",
-11452 => x"C0C0BFF9F99992A4",
-11451 => x"C0C0BFF9F99992F9",
-11450 => x"C0C0BFF9F99992C0",
-11449 => x"C0C0BFF9F9999990",
-11448 => x"C0C0BFF9F9999980",
-11447 => x"C0C0BFF9F99999F8",
-11446 => x"C0C0BFF9F9999982",
-11445 => x"C0C0BFF9F9999992",
-11444 => x"C0C0BFF9F9999999",
-11443 => x"C0C0BFF9F99999B0",
-11442 => x"C0C0BFF9F99999A4",
-11441 => x"C0C0BFF9F99999F9",
-11440 => x"C0C0BFF9F99999C0",
-11439 => x"C0C0BFF9F999B090",
-11438 => x"C0C0BFF9F999B080",
-11437 => x"C0C0BFF9F999B0F8",
-11436 => x"C0C0BFF9F999B082",
-11435 => x"C0C0BFF9F999B092",
-11434 => x"C0C0BFF9F999B099",
-11433 => x"C0C0BFF9F999B0B0",
-11432 => x"C0C0BFF9F999B0A4",
-11431 => x"C0C0BFF9F999B0F9",
-11430 => x"C0C0BFF9F999B0C0",
-11429 => x"C0C0BFF9F999A490",
-11428 => x"C0C0BFF9F999A480",
-11427 => x"C0C0BFF9F999A4F8",
-11426 => x"C0C0BFF9F999A482",
-11425 => x"C0C0BFF9F999A492",
-11424 => x"C0C0BFF9F999A499",
-11423 => x"C0C0BFF9F999A4B0",
-11422 => x"C0C0BFF9F999A4A4",
-11421 => x"C0C0BFF9F999A4F9",
-11420 => x"C0C0BFF9F999A4C0",
-11419 => x"C0C0BFF9F999F990",
-11418 => x"C0C0BFF9F999F980",
-11417 => x"C0C0BFF9F999F9F8",
-11416 => x"C0C0BFF9F999F982",
-11415 => x"C0C0BFF9F999F992",
-11414 => x"C0C0BFF9F999F999",
-11413 => x"C0C0BFF9F999F9B0",
-11412 => x"C0C0BFF9F999F9A4",
-11411 => x"C0C0BFF9F999F9F9",
-11410 => x"C0C0BFF9F999F9C0",
-11409 => x"C0C0BFF9F999C090",
-11408 => x"C0C0BFF9F999C080",
-11407 => x"C0C0BFF9F999C0F8",
-11406 => x"C0C0BFF9F999C082",
-11405 => x"C0C0BFF9F999C092",
-11404 => x"C0C0BFF9F999C099",
-11403 => x"C0C0BFF9F999C0B0",
-11402 => x"C0C0BFF9F999C0A4",
-11401 => x"C0C0BFF9F999C0F9",
-11400 => x"C0C0BFF9F999C0C0",
-11399 => x"C0C0BFF9F9B09090",
-11398 => x"C0C0BFF9F9B09080",
-11397 => x"C0C0BFF9F9B090F8",
-11396 => x"C0C0BFF9F9B09082",
-11395 => x"C0C0BFF9F9B09092",
-11394 => x"C0C0BFF9F9B09099",
-11393 => x"C0C0BFF9F9B090B0",
-11392 => x"C0C0BFF9F9B090A4",
-11391 => x"C0C0BFF9F9B090F9",
-11390 => x"C0C0BFF9F9B090C0",
-11389 => x"C0C0BFF9F9B08090",
-11388 => x"C0C0BFF9F9B08080",
-11387 => x"C0C0BFF9F9B080F8",
-11386 => x"C0C0BFF9F9B08082",
-11385 => x"C0C0BFF9F9B08092",
-11384 => x"C0C0BFF9F9B08099",
-11383 => x"C0C0BFF9F9B080B0",
-11382 => x"C0C0BFF9F9B080A4",
-11381 => x"C0C0BFF9F9B080F9",
-11380 => x"C0C0BFF9F9B080C0",
-11379 => x"C0C0BFF9F9B0F890",
-11378 => x"C0C0BFF9F9B0F880",
-11377 => x"C0C0BFF9F9B0F8F8",
-11376 => x"C0C0BFF9F9B0F882",
-11375 => x"C0C0BFF9F9B0F892",
-11374 => x"C0C0BFF9F9B0F899",
-11373 => x"C0C0BFF9F9B0F8B0",
-11372 => x"C0C0BFF9F9B0F8A4",
-11371 => x"C0C0BFF9F9B0F8F9",
-11370 => x"C0C0BFF9F9B0F8C0",
-11369 => x"C0C0BFF9F9B08290",
-11368 => x"C0C0BFF9F9B08280",
-11367 => x"C0C0BFF9F9B082F8",
-11366 => x"C0C0BFF9F9B08282",
-11365 => x"C0C0BFF9F9B08292",
-11364 => x"C0C0BFF9F9B08299",
-11363 => x"C0C0BFF9F9B082B0",
-11362 => x"C0C0BFF9F9B082A4",
-11361 => x"C0C0BFF9F9B082F9",
-11360 => x"C0C0BFF9F9B082C0",
-11359 => x"C0C0BFF9F9B09290",
-11358 => x"C0C0BFF9F9B09280",
-11357 => x"C0C0BFF9F9B092F8",
-11356 => x"C0C0BFF9F9B09282",
-11355 => x"C0C0BFF9F9B09292",
-11354 => x"C0C0BFF9F9B09299",
-11353 => x"C0C0BFF9F9B092B0",
-11352 => x"C0C0BFF9F9B092A4",
-11351 => x"C0C0BFF9F9B092F9",
-11350 => x"C0C0BFF9F9B092C0",
-11349 => x"C0C0BFF9F9B09990",
-11348 => x"C0C0BFF9F9B09980",
-11347 => x"C0C0BFF9F9B099F8",
-11346 => x"C0C0BFF9F9B09982",
-11345 => x"C0C0BFF9F9B09992",
-11344 => x"C0C0BFF9F9B09999",
-11343 => x"C0C0BFF9F9B099B0",
-11342 => x"C0C0BFF9F9B099A4",
-11341 => x"C0C0BFF9F9B099F9",
-11340 => x"C0C0BFF9F9B099C0",
-11339 => x"C0C0BFF9F9B0B090",
-11338 => x"C0C0BFF9F9B0B080",
-11337 => x"C0C0BFF9F9B0B0F8",
-11336 => x"C0C0BFF9F9B0B082",
-11335 => x"C0C0BFF9F9B0B092",
-11334 => x"C0C0BFF9F9B0B099",
-11333 => x"C0C0BFF9F9B0B0B0",
-11332 => x"C0C0BFF9F9B0B0A4",
-11331 => x"C0C0BFF9F9B0B0F9",
-11330 => x"C0C0BFF9F9B0B0C0",
-11329 => x"C0C0BFF9F9B0A490",
-11328 => x"C0C0BFF9F9B0A480",
-11327 => x"C0C0BFF9F9B0A4F8",
-11326 => x"C0C0BFF9F9B0A482",
-11325 => x"C0C0BFF9F9B0A492",
-11324 => x"C0C0BFF9F9B0A499",
-11323 => x"C0C0BFF9F9B0A4B0",
-11322 => x"C0C0BFF9F9B0A4A4",
-11321 => x"C0C0BFF9F9B0A4F9",
-11320 => x"C0C0BFF9F9B0A4C0",
-11319 => x"C0C0BFF9F9B0F990",
-11318 => x"C0C0BFF9F9B0F980",
-11317 => x"C0C0BFF9F9B0F9F8",
-11316 => x"C0C0BFF9F9B0F982",
-11315 => x"C0C0BFF9F9B0F992",
-11314 => x"C0C0BFF9F9B0F999",
-11313 => x"C0C0BFF9F9B0F9B0",
-11312 => x"C0C0BFF9F9B0F9A4",
-11311 => x"C0C0BFF9F9B0F9F9",
-11310 => x"C0C0BFF9F9B0F9C0",
-11309 => x"C0C0BFF9F9B0C090",
-11308 => x"C0C0BFF9F9B0C080",
-11307 => x"C0C0BFF9F9B0C0F8",
-11306 => x"C0C0BFF9F9B0C082",
-11305 => x"C0C0BFF9F9B0C092",
-11304 => x"C0C0BFF9F9B0C099",
-11303 => x"C0C0BFF9F9B0C0B0",
-11302 => x"C0C0BFF9F9B0C0A4",
-11301 => x"C0C0BFF9F9B0C0F9",
-11300 => x"C0C0BFF9F9B0C0C0",
-11299 => x"C0C0BFF9F9A49090",
-11298 => x"C0C0BFF9F9A49080",
-11297 => x"C0C0BFF9F9A490F8",
-11296 => x"C0C0BFF9F9A49082",
-11295 => x"C0C0BFF9F9A49092",
-11294 => x"C0C0BFF9F9A49099",
-11293 => x"C0C0BFF9F9A490B0",
-11292 => x"C0C0BFF9F9A490A4",
-11291 => x"C0C0BFF9F9A490F9",
-11290 => x"C0C0BFF9F9A490C0",
-11289 => x"C0C0BFF9F9A48090",
-11288 => x"C0C0BFF9F9A48080",
-11287 => x"C0C0BFF9F9A480F8",
-11286 => x"C0C0BFF9F9A48082",
-11285 => x"C0C0BFF9F9A48092",
-11284 => x"C0C0BFF9F9A48099",
-11283 => x"C0C0BFF9F9A480B0",
-11282 => x"C0C0BFF9F9A480A4",
-11281 => x"C0C0BFF9F9A480F9",
-11280 => x"C0C0BFF9F9A480C0",
-11279 => x"C0C0BFF9F9A4F890",
-11278 => x"C0C0BFF9F9A4F880",
-11277 => x"C0C0BFF9F9A4F8F8",
-11276 => x"C0C0BFF9F9A4F882",
-11275 => x"C0C0BFF9F9A4F892",
-11274 => x"C0C0BFF9F9A4F899",
-11273 => x"C0C0BFF9F9A4F8B0",
-11272 => x"C0C0BFF9F9A4F8A4",
-11271 => x"C0C0BFF9F9A4F8F9",
-11270 => x"C0C0BFF9F9A4F8C0",
-11269 => x"C0C0BFF9F9A48290",
-11268 => x"C0C0BFF9F9A48280",
-11267 => x"C0C0BFF9F9A482F8",
-11266 => x"C0C0BFF9F9A48282",
-11265 => x"C0C0BFF9F9A48292",
-11264 => x"C0C0BFF9F9A48299",
-11263 => x"C0C0BFF9F9A482B0",
-11262 => x"C0C0BFF9F9A482A4",
-11261 => x"C0C0BFF9F9A482F9",
-11260 => x"C0C0BFF9F9A482C0",
-11259 => x"C0C0BFF9F9A49290",
-11258 => x"C0C0BFF9F9A49280",
-11257 => x"C0C0BFF9F9A492F8",
-11256 => x"C0C0BFF9F9A49282",
-11255 => x"C0C0BFF9F9A49292",
-11254 => x"C0C0BFF9F9A49299",
-11253 => x"C0C0BFF9F9A492B0",
-11252 => x"C0C0BFF9F9A492A4",
-11251 => x"C0C0BFF9F9A492F9",
-11250 => x"C0C0BFF9F9A492C0",
-11249 => x"C0C0BFF9F9A49990",
-11248 => x"C0C0BFF9F9A49980",
-11247 => x"C0C0BFF9F9A499F8",
-11246 => x"C0C0BFF9F9A49982",
-11245 => x"C0C0BFF9F9A49992",
-11244 => x"C0C0BFF9F9A49999",
-11243 => x"C0C0BFF9F9A499B0",
-11242 => x"C0C0BFF9F9A499A4",
-11241 => x"C0C0BFF9F9A499F9",
-11240 => x"C0C0BFF9F9A499C0",
-11239 => x"C0C0BFF9F9A4B090",
-11238 => x"C0C0BFF9F9A4B080",
-11237 => x"C0C0BFF9F9A4B0F8",
-11236 => x"C0C0BFF9F9A4B082",
-11235 => x"C0C0BFF9F9A4B092",
-11234 => x"C0C0BFF9F9A4B099",
-11233 => x"C0C0BFF9F9A4B0B0",
-11232 => x"C0C0BFF9F9A4B0A4",
-11231 => x"C0C0BFF9F9A4B0F9",
-11230 => x"C0C0BFF9F9A4B0C0",
-11229 => x"C0C0BFF9F9A4A490",
-11228 => x"C0C0BFF9F9A4A480",
-11227 => x"C0C0BFF9F9A4A4F8",
-11226 => x"C0C0BFF9F9A4A482",
-11225 => x"C0C0BFF9F9A4A492",
-11224 => x"C0C0BFF9F9A4A499",
-11223 => x"C0C0BFF9F9A4A4B0",
-11222 => x"C0C0BFF9F9A4A4A4",
-11221 => x"C0C0BFF9F9A4A4F9",
-11220 => x"C0C0BFF9F9A4A4C0",
-11219 => x"C0C0BFF9F9A4F990",
-11218 => x"C0C0BFF9F9A4F980",
-11217 => x"C0C0BFF9F9A4F9F8",
-11216 => x"C0C0BFF9F9A4F982",
-11215 => x"C0C0BFF9F9A4F992",
-11214 => x"C0C0BFF9F9A4F999",
-11213 => x"C0C0BFF9F9A4F9B0",
-11212 => x"C0C0BFF9F9A4F9A4",
-11211 => x"C0C0BFF9F9A4F9F9",
-11210 => x"C0C0BFF9F9A4F9C0",
-11209 => x"C0C0BFF9F9A4C090",
-11208 => x"C0C0BFF9F9A4C080",
-11207 => x"C0C0BFF9F9A4C0F8",
-11206 => x"C0C0BFF9F9A4C082",
-11205 => x"C0C0BFF9F9A4C092",
-11204 => x"C0C0BFF9F9A4C099",
-11203 => x"C0C0BFF9F9A4C0B0",
-11202 => x"C0C0BFF9F9A4C0A4",
-11201 => x"C0C0BFF9F9A4C0F9",
-11200 => x"C0C0BFF9F9A4C0C0",
-11199 => x"C0C0BFF9F9F99090",
-11198 => x"C0C0BFF9F9F99080",
-11197 => x"C0C0BFF9F9F990F8",
-11196 => x"C0C0BFF9F9F99082",
-11195 => x"C0C0BFF9F9F99092",
-11194 => x"C0C0BFF9F9F99099",
-11193 => x"C0C0BFF9F9F990B0",
-11192 => x"C0C0BFF9F9F990A4",
-11191 => x"C0C0BFF9F9F990F9",
-11190 => x"C0C0BFF9F9F990C0",
-11189 => x"C0C0BFF9F9F98090",
-11188 => x"C0C0BFF9F9F98080",
-11187 => x"C0C0BFF9F9F980F8",
-11186 => x"C0C0BFF9F9F98082",
-11185 => x"C0C0BFF9F9F98092",
-11184 => x"C0C0BFF9F9F98099",
-11183 => x"C0C0BFF9F9F980B0",
-11182 => x"C0C0BFF9F9F980A4",
-11181 => x"C0C0BFF9F9F980F9",
-11180 => x"C0C0BFF9F9F980C0",
-11179 => x"C0C0BFF9F9F9F890",
-11178 => x"C0C0BFF9F9F9F880",
-11177 => x"C0C0BFF9F9F9F8F8",
-11176 => x"C0C0BFF9F9F9F882",
-11175 => x"C0C0BFF9F9F9F892",
-11174 => x"C0C0BFF9F9F9F899",
-11173 => x"C0C0BFF9F9F9F8B0",
-11172 => x"C0C0BFF9F9F9F8A4",
-11171 => x"C0C0BFF9F9F9F8F9",
-11170 => x"C0C0BFF9F9F9F8C0",
-11169 => x"C0C0BFF9F9F98290",
-11168 => x"C0C0BFF9F9F98280",
-11167 => x"C0C0BFF9F9F982F8",
-11166 => x"C0C0BFF9F9F98282",
-11165 => x"C0C0BFF9F9F98292",
-11164 => x"C0C0BFF9F9F98299",
-11163 => x"C0C0BFF9F9F982B0",
-11162 => x"C0C0BFF9F9F982A4",
-11161 => x"C0C0BFF9F9F982F9",
-11160 => x"C0C0BFF9F9F982C0",
-11159 => x"C0C0BFF9F9F99290",
-11158 => x"C0C0BFF9F9F99280",
-11157 => x"C0C0BFF9F9F992F8",
-11156 => x"C0C0BFF9F9F99282",
-11155 => x"C0C0BFF9F9F99292",
-11154 => x"C0C0BFF9F9F99299",
-11153 => x"C0C0BFF9F9F992B0",
-11152 => x"C0C0BFF9F9F992A4",
-11151 => x"C0C0BFF9F9F992F9",
-11150 => x"C0C0BFF9F9F992C0",
-11149 => x"C0C0BFF9F9F99990",
-11148 => x"C0C0BFF9F9F99980",
-11147 => x"C0C0BFF9F9F999F8",
-11146 => x"C0C0BFF9F9F99982",
-11145 => x"C0C0BFF9F9F99992",
-11144 => x"C0C0BFF9F9F99999",
-11143 => x"C0C0BFF9F9F999B0",
-11142 => x"C0C0BFF9F9F999A4",
-11141 => x"C0C0BFF9F9F999F9",
-11140 => x"C0C0BFF9F9F999C0",
-11139 => x"C0C0BFF9F9F9B090",
-11138 => x"C0C0BFF9F9F9B080",
-11137 => x"C0C0BFF9F9F9B0F8",
-11136 => x"C0C0BFF9F9F9B082",
-11135 => x"C0C0BFF9F9F9B092",
-11134 => x"C0C0BFF9F9F9B099",
-11133 => x"C0C0BFF9F9F9B0B0",
-11132 => x"C0C0BFF9F9F9B0A4",
-11131 => x"C0C0BFF9F9F9B0F9",
-11130 => x"C0C0BFF9F9F9B0C0",
-11129 => x"C0C0BFF9F9F9A490",
-11128 => x"C0C0BFF9F9F9A480",
-11127 => x"C0C0BFF9F9F9A4F8",
-11126 => x"C0C0BFF9F9F9A482",
-11125 => x"C0C0BFF9F9F9A492",
-11124 => x"C0C0BFF9F9F9A499",
-11123 => x"C0C0BFF9F9F9A4B0",
-11122 => x"C0C0BFF9F9F9A4A4",
-11121 => x"C0C0BFF9F9F9A4F9",
-11120 => x"C0C0BFF9F9F9A4C0",
-11119 => x"C0C0BFF9F9F9F990",
-11118 => x"C0C0BFF9F9F9F980",
-11117 => x"C0C0BFF9F9F9F9F8",
-11116 => x"C0C0BFF9F9F9F982",
-11115 => x"C0C0BFF9F9F9F992",
-11114 => x"C0C0BFF9F9F9F999",
-11113 => x"C0C0BFF9F9F9F9B0",
-11112 => x"C0C0BFF9F9F9F9A4",
-11111 => x"C0C0BFF9F9F9F9F9",
-11110 => x"C0C0BFF9F9F9F9C0",
-11109 => x"C0C0BFF9F9F9C090",
-11108 => x"C0C0BFF9F9F9C080",
-11107 => x"C0C0BFF9F9F9C0F8",
-11106 => x"C0C0BFF9F9F9C082",
-11105 => x"C0C0BFF9F9F9C092",
-11104 => x"C0C0BFF9F9F9C099",
-11103 => x"C0C0BFF9F9F9C0B0",
-11102 => x"C0C0BFF9F9F9C0A4",
-11101 => x"C0C0BFF9F9F9C0F9",
-11100 => x"C0C0BFF9F9F9C0C0",
-11099 => x"C0C0BFF9F9C09090",
-11098 => x"C0C0BFF9F9C09080",
-11097 => x"C0C0BFF9F9C090F8",
-11096 => x"C0C0BFF9F9C09082",
-11095 => x"C0C0BFF9F9C09092",
-11094 => x"C0C0BFF9F9C09099",
-11093 => x"C0C0BFF9F9C090B0",
-11092 => x"C0C0BFF9F9C090A4",
-11091 => x"C0C0BFF9F9C090F9",
-11090 => x"C0C0BFF9F9C090C0",
-11089 => x"C0C0BFF9F9C08090",
-11088 => x"C0C0BFF9F9C08080",
-11087 => x"C0C0BFF9F9C080F8",
-11086 => x"C0C0BFF9F9C08082",
-11085 => x"C0C0BFF9F9C08092",
-11084 => x"C0C0BFF9F9C08099",
-11083 => x"C0C0BFF9F9C080B0",
-11082 => x"C0C0BFF9F9C080A4",
-11081 => x"C0C0BFF9F9C080F9",
-11080 => x"C0C0BFF9F9C080C0",
-11079 => x"C0C0BFF9F9C0F890",
-11078 => x"C0C0BFF9F9C0F880",
-11077 => x"C0C0BFF9F9C0F8F8",
-11076 => x"C0C0BFF9F9C0F882",
-11075 => x"C0C0BFF9F9C0F892",
-11074 => x"C0C0BFF9F9C0F899",
-11073 => x"C0C0BFF9F9C0F8B0",
-11072 => x"C0C0BFF9F9C0F8A4",
-11071 => x"C0C0BFF9F9C0F8F9",
-11070 => x"C0C0BFF9F9C0F8C0",
-11069 => x"C0C0BFF9F9C08290",
-11068 => x"C0C0BFF9F9C08280",
-11067 => x"C0C0BFF9F9C082F8",
-11066 => x"C0C0BFF9F9C08282",
-11065 => x"C0C0BFF9F9C08292",
-11064 => x"C0C0BFF9F9C08299",
-11063 => x"C0C0BFF9F9C082B0",
-11062 => x"C0C0BFF9F9C082A4",
-11061 => x"C0C0BFF9F9C082F9",
-11060 => x"C0C0BFF9F9C082C0",
-11059 => x"C0C0BFF9F9C09290",
-11058 => x"C0C0BFF9F9C09280",
-11057 => x"C0C0BFF9F9C092F8",
-11056 => x"C0C0BFF9F9C09282",
-11055 => x"C0C0BFF9F9C09292",
-11054 => x"C0C0BFF9F9C09299",
-11053 => x"C0C0BFF9F9C092B0",
-11052 => x"C0C0BFF9F9C092A4",
-11051 => x"C0C0BFF9F9C092F9",
-11050 => x"C0C0BFF9F9C092C0",
-11049 => x"C0C0BFF9F9C09990",
-11048 => x"C0C0BFF9F9C09980",
-11047 => x"C0C0BFF9F9C099F8",
-11046 => x"C0C0BFF9F9C09982",
-11045 => x"C0C0BFF9F9C09992",
-11044 => x"C0C0BFF9F9C09999",
-11043 => x"C0C0BFF9F9C099B0",
-11042 => x"C0C0BFF9F9C099A4",
-11041 => x"C0C0BFF9F9C099F9",
-11040 => x"C0C0BFF9F9C099C0",
-11039 => x"C0C0BFF9F9C0B090",
-11038 => x"C0C0BFF9F9C0B080",
-11037 => x"C0C0BFF9F9C0B0F8",
-11036 => x"C0C0BFF9F9C0B082",
-11035 => x"C0C0BFF9F9C0B092",
-11034 => x"C0C0BFF9F9C0B099",
-11033 => x"C0C0BFF9F9C0B0B0",
-11032 => x"C0C0BFF9F9C0B0A4",
-11031 => x"C0C0BFF9F9C0B0F9",
-11030 => x"C0C0BFF9F9C0B0C0",
-11029 => x"C0C0BFF9F9C0A490",
-11028 => x"C0C0BFF9F9C0A480",
-11027 => x"C0C0BFF9F9C0A4F8",
-11026 => x"C0C0BFF9F9C0A482",
-11025 => x"C0C0BFF9F9C0A492",
-11024 => x"C0C0BFF9F9C0A499",
-11023 => x"C0C0BFF9F9C0A4B0",
-11022 => x"C0C0BFF9F9C0A4A4",
-11021 => x"C0C0BFF9F9C0A4F9",
-11020 => x"C0C0BFF9F9C0A4C0",
-11019 => x"C0C0BFF9F9C0F990",
-11018 => x"C0C0BFF9F9C0F980",
-11017 => x"C0C0BFF9F9C0F9F8",
-11016 => x"C0C0BFF9F9C0F982",
-11015 => x"C0C0BFF9F9C0F992",
-11014 => x"C0C0BFF9F9C0F999",
-11013 => x"C0C0BFF9F9C0F9B0",
-11012 => x"C0C0BFF9F9C0F9A4",
-11011 => x"C0C0BFF9F9C0F9F9",
-11010 => x"C0C0BFF9F9C0F9C0",
-11009 => x"C0C0BFF9F9C0C090",
-11008 => x"C0C0BFF9F9C0C080",
-11007 => x"C0C0BFF9F9C0C0F8",
-11006 => x"C0C0BFF9F9C0C082",
-11005 => x"C0C0BFF9F9C0C092",
-11004 => x"C0C0BFF9F9C0C099",
-11003 => x"C0C0BFF9F9C0C0B0",
-11002 => x"C0C0BFF9F9C0C0A4",
-11001 => x"C0C0BFF9F9C0C0F9",
-11000 => x"C0C0BFF9F9C0C0C0",
-10999 => x"C0C0BFF9C0909090",
-10998 => x"C0C0BFF9C0909080",
-10997 => x"C0C0BFF9C09090F8",
-10996 => x"C0C0BFF9C0909082",
-10995 => x"C0C0BFF9C0909092",
-10994 => x"C0C0BFF9C0909099",
-10993 => x"C0C0BFF9C09090B0",
-10992 => x"C0C0BFF9C09090A4",
-10991 => x"C0C0BFF9C09090F9",
-10990 => x"C0C0BFF9C09090C0",
-10989 => x"C0C0BFF9C0908090",
-10988 => x"C0C0BFF9C0908080",
-10987 => x"C0C0BFF9C09080F8",
-10986 => x"C0C0BFF9C0908082",
-10985 => x"C0C0BFF9C0908092",
-10984 => x"C0C0BFF9C0908099",
-10983 => x"C0C0BFF9C09080B0",
-10982 => x"C0C0BFF9C09080A4",
-10981 => x"C0C0BFF9C09080F9",
-10980 => x"C0C0BFF9C09080C0",
-10979 => x"C0C0BFF9C090F890",
-10978 => x"C0C0BFF9C090F880",
-10977 => x"C0C0BFF9C090F8F8",
-10976 => x"C0C0BFF9C090F882",
-10975 => x"C0C0BFF9C090F892",
-10974 => x"C0C0BFF9C090F899",
-10973 => x"C0C0BFF9C090F8B0",
-10972 => x"C0C0BFF9C090F8A4",
-10971 => x"C0C0BFF9C090F8F9",
-10970 => x"C0C0BFF9C090F8C0",
-10969 => x"C0C0BFF9C0908290",
-10968 => x"C0C0BFF9C0908280",
-10967 => x"C0C0BFF9C09082F8",
-10966 => x"C0C0BFF9C0908282",
-10965 => x"C0C0BFF9C0908292",
-10964 => x"C0C0BFF9C0908299",
-10963 => x"C0C0BFF9C09082B0",
-10962 => x"C0C0BFF9C09082A4",
-10961 => x"C0C0BFF9C09082F9",
-10960 => x"C0C0BFF9C09082C0",
-10959 => x"C0C0BFF9C0909290",
-10958 => x"C0C0BFF9C0909280",
-10957 => x"C0C0BFF9C09092F8",
-10956 => x"C0C0BFF9C0909282",
-10955 => x"C0C0BFF9C0909292",
-10954 => x"C0C0BFF9C0909299",
-10953 => x"C0C0BFF9C09092B0",
-10952 => x"C0C0BFF9C09092A4",
-10951 => x"C0C0BFF9C09092F9",
-10950 => x"C0C0BFF9C09092C0",
-10949 => x"C0C0BFF9C0909990",
-10948 => x"C0C0BFF9C0909980",
-10947 => x"C0C0BFF9C09099F8",
-10946 => x"C0C0BFF9C0909982",
-10945 => x"C0C0BFF9C0909992",
-10944 => x"C0C0BFF9C0909999",
-10943 => x"C0C0BFF9C09099B0",
-10942 => x"C0C0BFF9C09099A4",
-10941 => x"C0C0BFF9C09099F9",
-10940 => x"C0C0BFF9C09099C0",
-10939 => x"C0C0BFF9C090B090",
-10938 => x"C0C0BFF9C090B080",
-10937 => x"C0C0BFF9C090B0F8",
-10936 => x"C0C0BFF9C090B082",
-10935 => x"C0C0BFF9C090B092",
-10934 => x"C0C0BFF9C090B099",
-10933 => x"C0C0BFF9C090B0B0",
-10932 => x"C0C0BFF9C090B0A4",
-10931 => x"C0C0BFF9C090B0F9",
-10930 => x"C0C0BFF9C090B0C0",
-10929 => x"C0C0BFF9C090A490",
-10928 => x"C0C0BFF9C090A480",
-10927 => x"C0C0BFF9C090A4F8",
-10926 => x"C0C0BFF9C090A482",
-10925 => x"C0C0BFF9C090A492",
-10924 => x"C0C0BFF9C090A499",
-10923 => x"C0C0BFF9C090A4B0",
-10922 => x"C0C0BFF9C090A4A4",
-10921 => x"C0C0BFF9C090A4F9",
-10920 => x"C0C0BFF9C090A4C0",
-10919 => x"C0C0BFF9C090F990",
-10918 => x"C0C0BFF9C090F980",
-10917 => x"C0C0BFF9C090F9F8",
-10916 => x"C0C0BFF9C090F982",
-10915 => x"C0C0BFF9C090F992",
-10914 => x"C0C0BFF9C090F999",
-10913 => x"C0C0BFF9C090F9B0",
-10912 => x"C0C0BFF9C090F9A4",
-10911 => x"C0C0BFF9C090F9F9",
-10910 => x"C0C0BFF9C090F9C0",
-10909 => x"C0C0BFF9C090C090",
-10908 => x"C0C0BFF9C090C080",
-10907 => x"C0C0BFF9C090C0F8",
-10906 => x"C0C0BFF9C090C082",
-10905 => x"C0C0BFF9C090C092",
-10904 => x"C0C0BFF9C090C099",
-10903 => x"C0C0BFF9C090C0B0",
-10902 => x"C0C0BFF9C090C0A4",
-10901 => x"C0C0BFF9C090C0F9",
-10900 => x"C0C0BFF9C090C0C0",
-10899 => x"C0C0BFF9C0809090",
-10898 => x"C0C0BFF9C0809080",
-10897 => x"C0C0BFF9C08090F8",
-10896 => x"C0C0BFF9C0809082",
-10895 => x"C0C0BFF9C0809092",
-10894 => x"C0C0BFF9C0809099",
-10893 => x"C0C0BFF9C08090B0",
-10892 => x"C0C0BFF9C08090A4",
-10891 => x"C0C0BFF9C08090F9",
-10890 => x"C0C0BFF9C08090C0",
-10889 => x"C0C0BFF9C0808090",
-10888 => x"C0C0BFF9C0808080",
-10887 => x"C0C0BFF9C08080F8",
-10886 => x"C0C0BFF9C0808082",
-10885 => x"C0C0BFF9C0808092",
-10884 => x"C0C0BFF9C0808099",
-10883 => x"C0C0BFF9C08080B0",
-10882 => x"C0C0BFF9C08080A4",
-10881 => x"C0C0BFF9C08080F9",
-10880 => x"C0C0BFF9C08080C0",
-10879 => x"C0C0BFF9C080F890",
-10878 => x"C0C0BFF9C080F880",
-10877 => x"C0C0BFF9C080F8F8",
-10876 => x"C0C0BFF9C080F882",
-10875 => x"C0C0BFF9C080F892",
-10874 => x"C0C0BFF9C080F899",
-10873 => x"C0C0BFF9C080F8B0",
-10872 => x"C0C0BFF9C080F8A4",
-10871 => x"C0C0BFF9C080F8F9",
-10870 => x"C0C0BFF9C080F8C0",
-10869 => x"C0C0BFF9C0808290",
-10868 => x"C0C0BFF9C0808280",
-10867 => x"C0C0BFF9C08082F8",
-10866 => x"C0C0BFF9C0808282",
-10865 => x"C0C0BFF9C0808292",
-10864 => x"C0C0BFF9C0808299",
-10863 => x"C0C0BFF9C08082B0",
-10862 => x"C0C0BFF9C08082A4",
-10861 => x"C0C0BFF9C08082F9",
-10860 => x"C0C0BFF9C08082C0",
-10859 => x"C0C0BFF9C0809290",
-10858 => x"C0C0BFF9C0809280",
-10857 => x"C0C0BFF9C08092F8",
-10856 => x"C0C0BFF9C0809282",
-10855 => x"C0C0BFF9C0809292",
-10854 => x"C0C0BFF9C0809299",
-10853 => x"C0C0BFF9C08092B0",
-10852 => x"C0C0BFF9C08092A4",
-10851 => x"C0C0BFF9C08092F9",
-10850 => x"C0C0BFF9C08092C0",
-10849 => x"C0C0BFF9C0809990",
-10848 => x"C0C0BFF9C0809980",
-10847 => x"C0C0BFF9C08099F8",
-10846 => x"C0C0BFF9C0809982",
-10845 => x"C0C0BFF9C0809992",
-10844 => x"C0C0BFF9C0809999",
-10843 => x"C0C0BFF9C08099B0",
-10842 => x"C0C0BFF9C08099A4",
-10841 => x"C0C0BFF9C08099F9",
-10840 => x"C0C0BFF9C08099C0",
-10839 => x"C0C0BFF9C080B090",
-10838 => x"C0C0BFF9C080B080",
-10837 => x"C0C0BFF9C080B0F8",
-10836 => x"C0C0BFF9C080B082",
-10835 => x"C0C0BFF9C080B092",
-10834 => x"C0C0BFF9C080B099",
-10833 => x"C0C0BFF9C080B0B0",
-10832 => x"C0C0BFF9C080B0A4",
-10831 => x"C0C0BFF9C080B0F9",
-10830 => x"C0C0BFF9C080B0C0",
-10829 => x"C0C0BFF9C080A490",
-10828 => x"C0C0BFF9C080A480",
-10827 => x"C0C0BFF9C080A4F8",
-10826 => x"C0C0BFF9C080A482",
-10825 => x"C0C0BFF9C080A492",
-10824 => x"C0C0BFF9C080A499",
-10823 => x"C0C0BFF9C080A4B0",
-10822 => x"C0C0BFF9C080A4A4",
-10821 => x"C0C0BFF9C080A4F9",
-10820 => x"C0C0BFF9C080A4C0",
-10819 => x"C0C0BFF9C080F990",
-10818 => x"C0C0BFF9C080F980",
-10817 => x"C0C0BFF9C080F9F8",
-10816 => x"C0C0BFF9C080F982",
-10815 => x"C0C0BFF9C080F992",
-10814 => x"C0C0BFF9C080F999",
-10813 => x"C0C0BFF9C080F9B0",
-10812 => x"C0C0BFF9C080F9A4",
-10811 => x"C0C0BFF9C080F9F9",
-10810 => x"C0C0BFF9C080F9C0",
-10809 => x"C0C0BFF9C080C090",
-10808 => x"C0C0BFF9C080C080",
-10807 => x"C0C0BFF9C080C0F8",
-10806 => x"C0C0BFF9C080C082",
-10805 => x"C0C0BFF9C080C092",
-10804 => x"C0C0BFF9C080C099",
-10803 => x"C0C0BFF9C080C0B0",
-10802 => x"C0C0BFF9C080C0A4",
-10801 => x"C0C0BFF9C080C0F9",
-10800 => x"C0C0BFF9C080C0C0",
-10799 => x"C0C0BFF9C0F89090",
-10798 => x"C0C0BFF9C0F89080",
-10797 => x"C0C0BFF9C0F890F8",
-10796 => x"C0C0BFF9C0F89082",
-10795 => x"C0C0BFF9C0F89092",
-10794 => x"C0C0BFF9C0F89099",
-10793 => x"C0C0BFF9C0F890B0",
-10792 => x"C0C0BFF9C0F890A4",
-10791 => x"C0C0BFF9C0F890F9",
-10790 => x"C0C0BFF9C0F890C0",
-10789 => x"C0C0BFF9C0F88090",
-10788 => x"C0C0BFF9C0F88080",
-10787 => x"C0C0BFF9C0F880F8",
-10786 => x"C0C0BFF9C0F88082",
-10785 => x"C0C0BFF9C0F88092",
-10784 => x"C0C0BFF9C0F88099",
-10783 => x"C0C0BFF9C0F880B0",
-10782 => x"C0C0BFF9C0F880A4",
-10781 => x"C0C0BFF9C0F880F9",
-10780 => x"C0C0BFF9C0F880C0",
-10779 => x"C0C0BFF9C0F8F890",
-10778 => x"C0C0BFF9C0F8F880",
-10777 => x"C0C0BFF9C0F8F8F8",
-10776 => x"C0C0BFF9C0F8F882",
-10775 => x"C0C0BFF9C0F8F892",
-10774 => x"C0C0BFF9C0F8F899",
-10773 => x"C0C0BFF9C0F8F8B0",
-10772 => x"C0C0BFF9C0F8F8A4",
-10771 => x"C0C0BFF9C0F8F8F9",
-10770 => x"C0C0BFF9C0F8F8C0",
-10769 => x"C0C0BFF9C0F88290",
-10768 => x"C0C0BFF9C0F88280",
-10767 => x"C0C0BFF9C0F882F8",
-10766 => x"C0C0BFF9C0F88282",
-10765 => x"C0C0BFF9C0F88292",
-10764 => x"C0C0BFF9C0F88299",
-10763 => x"C0C0BFF9C0F882B0",
-10762 => x"C0C0BFF9C0F882A4",
-10761 => x"C0C0BFF9C0F882F9",
-10760 => x"C0C0BFF9C0F882C0",
-10759 => x"C0C0BFF9C0F89290",
-10758 => x"C0C0BFF9C0F89280",
-10757 => x"C0C0BFF9C0F892F8",
-10756 => x"C0C0BFF9C0F89282",
-10755 => x"C0C0BFF9C0F89292",
-10754 => x"C0C0BFF9C0F89299",
-10753 => x"C0C0BFF9C0F892B0",
-10752 => x"C0C0BFF9C0F892A4",
-10751 => x"C0C0BFF9C0F892F9",
-10750 => x"C0C0BFF9C0F892C0",
-10749 => x"C0C0BFF9C0F89990",
-10748 => x"C0C0BFF9C0F89980",
-10747 => x"C0C0BFF9C0F899F8",
-10746 => x"C0C0BFF9C0F89982",
-10745 => x"C0C0BFF9C0F89992",
-10744 => x"C0C0BFF9C0F89999",
-10743 => x"C0C0BFF9C0F899B0",
-10742 => x"C0C0BFF9C0F899A4",
-10741 => x"C0C0BFF9C0F899F9",
-10740 => x"C0C0BFF9C0F899C0",
-10739 => x"C0C0BFF9C0F8B090",
-10738 => x"C0C0BFF9C0F8B080",
-10737 => x"C0C0BFF9C0F8B0F8",
-10736 => x"C0C0BFF9C0F8B082",
-10735 => x"C0C0BFF9C0F8B092",
-10734 => x"C0C0BFF9C0F8B099",
-10733 => x"C0C0BFF9C0F8B0B0",
-10732 => x"C0C0BFF9C0F8B0A4",
-10731 => x"C0C0BFF9C0F8B0F9",
-10730 => x"C0C0BFF9C0F8B0C0",
-10729 => x"C0C0BFF9C0F8A490",
-10728 => x"C0C0BFF9C0F8A480",
-10727 => x"C0C0BFF9C0F8A4F8",
-10726 => x"C0C0BFF9C0F8A482",
-10725 => x"C0C0BFF9C0F8A492",
-10724 => x"C0C0BFF9C0F8A499",
-10723 => x"C0C0BFF9C0F8A4B0",
-10722 => x"C0C0BFF9C0F8A4A4",
-10721 => x"C0C0BFF9C0F8A4F9",
-10720 => x"C0C0BFF9C0F8A4C0",
-10719 => x"C0C0BFF9C0F8F990",
-10718 => x"C0C0BFF9C0F8F980",
-10717 => x"C0C0BFF9C0F8F9F8",
-10716 => x"C0C0BFF9C0F8F982",
-10715 => x"C0C0BFF9C0F8F992",
-10714 => x"C0C0BFF9C0F8F999",
-10713 => x"C0C0BFF9C0F8F9B0",
-10712 => x"C0C0BFF9C0F8F9A4",
-10711 => x"C0C0BFF9C0F8F9F9",
-10710 => x"C0C0BFF9C0F8F9C0",
-10709 => x"C0C0BFF9C0F8C090",
-10708 => x"C0C0BFF9C0F8C080",
-10707 => x"C0C0BFF9C0F8C0F8",
-10706 => x"C0C0BFF9C0F8C082",
-10705 => x"C0C0BFF9C0F8C092",
-10704 => x"C0C0BFF9C0F8C099",
-10703 => x"C0C0BFF9C0F8C0B0",
-10702 => x"C0C0BFF9C0F8C0A4",
-10701 => x"C0C0BFF9C0F8C0F9",
-10700 => x"C0C0BFF9C0F8C0C0",
-10699 => x"C0C0BFF9C0829090",
-10698 => x"C0C0BFF9C0829080",
-10697 => x"C0C0BFF9C08290F8",
-10696 => x"C0C0BFF9C0829082",
-10695 => x"C0C0BFF9C0829092",
-10694 => x"C0C0BFF9C0829099",
-10693 => x"C0C0BFF9C08290B0",
-10692 => x"C0C0BFF9C08290A4",
-10691 => x"C0C0BFF9C08290F9",
-10690 => x"C0C0BFF9C08290C0",
-10689 => x"C0C0BFF9C0828090",
-10688 => x"C0C0BFF9C0828080",
-10687 => x"C0C0BFF9C08280F8",
-10686 => x"C0C0BFF9C0828082",
-10685 => x"C0C0BFF9C0828092",
-10684 => x"C0C0BFF9C0828099",
-10683 => x"C0C0BFF9C08280B0",
-10682 => x"C0C0BFF9C08280A4",
-10681 => x"C0C0BFF9C08280F9",
-10680 => x"C0C0BFF9C08280C0",
-10679 => x"C0C0BFF9C082F890",
-10678 => x"C0C0BFF9C082F880",
-10677 => x"C0C0BFF9C082F8F8",
-10676 => x"C0C0BFF9C082F882",
-10675 => x"C0C0BFF9C082F892",
-10674 => x"C0C0BFF9C082F899",
-10673 => x"C0C0BFF9C082F8B0",
-10672 => x"C0C0BFF9C082F8A4",
-10671 => x"C0C0BFF9C082F8F9",
-10670 => x"C0C0BFF9C082F8C0",
-10669 => x"C0C0BFF9C0828290",
-10668 => x"C0C0BFF9C0828280",
-10667 => x"C0C0BFF9C08282F8",
-10666 => x"C0C0BFF9C0828282",
-10665 => x"C0C0BFF9C0828292",
-10664 => x"C0C0BFF9C0828299",
-10663 => x"C0C0BFF9C08282B0",
-10662 => x"C0C0BFF9C08282A4",
-10661 => x"C0C0BFF9C08282F9",
-10660 => x"C0C0BFF9C08282C0",
-10659 => x"C0C0BFF9C0829290",
-10658 => x"C0C0BFF9C0829280",
-10657 => x"C0C0BFF9C08292F8",
-10656 => x"C0C0BFF9C0829282",
-10655 => x"C0C0BFF9C0829292",
-10654 => x"C0C0BFF9C0829299",
-10653 => x"C0C0BFF9C08292B0",
-10652 => x"C0C0BFF9C08292A4",
-10651 => x"C0C0BFF9C08292F9",
-10650 => x"C0C0BFF9C08292C0",
-10649 => x"C0C0BFF9C0829990",
-10648 => x"C0C0BFF9C0829980",
-10647 => x"C0C0BFF9C08299F8",
-10646 => x"C0C0BFF9C0829982",
-10645 => x"C0C0BFF9C0829992",
-10644 => x"C0C0BFF9C0829999",
-10643 => x"C0C0BFF9C08299B0",
-10642 => x"C0C0BFF9C08299A4",
-10641 => x"C0C0BFF9C08299F9",
-10640 => x"C0C0BFF9C08299C0",
-10639 => x"C0C0BFF9C082B090",
-10638 => x"C0C0BFF9C082B080",
-10637 => x"C0C0BFF9C082B0F8",
-10636 => x"C0C0BFF9C082B082",
-10635 => x"C0C0BFF9C082B092",
-10634 => x"C0C0BFF9C082B099",
-10633 => x"C0C0BFF9C082B0B0",
-10632 => x"C0C0BFF9C082B0A4",
-10631 => x"C0C0BFF9C082B0F9",
-10630 => x"C0C0BFF9C082B0C0",
-10629 => x"C0C0BFF9C082A490",
-10628 => x"C0C0BFF9C082A480",
-10627 => x"C0C0BFF9C082A4F8",
-10626 => x"C0C0BFF9C082A482",
-10625 => x"C0C0BFF9C082A492",
-10624 => x"C0C0BFF9C082A499",
-10623 => x"C0C0BFF9C082A4B0",
-10622 => x"C0C0BFF9C082A4A4",
-10621 => x"C0C0BFF9C082A4F9",
-10620 => x"C0C0BFF9C082A4C0",
-10619 => x"C0C0BFF9C082F990",
-10618 => x"C0C0BFF9C082F980",
-10617 => x"C0C0BFF9C082F9F8",
-10616 => x"C0C0BFF9C082F982",
-10615 => x"C0C0BFF9C082F992",
-10614 => x"C0C0BFF9C082F999",
-10613 => x"C0C0BFF9C082F9B0",
-10612 => x"C0C0BFF9C082F9A4",
-10611 => x"C0C0BFF9C082F9F9",
-10610 => x"C0C0BFF9C082F9C0",
-10609 => x"C0C0BFF9C082C090",
-10608 => x"C0C0BFF9C082C080",
-10607 => x"C0C0BFF9C082C0F8",
-10606 => x"C0C0BFF9C082C082",
-10605 => x"C0C0BFF9C082C092",
-10604 => x"C0C0BFF9C082C099",
-10603 => x"C0C0BFF9C082C0B0",
-10602 => x"C0C0BFF9C082C0A4",
-10601 => x"C0C0BFF9C082C0F9",
-10600 => x"C0C0BFF9C082C0C0",
-10599 => x"C0C0BFF9C0929090",
-10598 => x"C0C0BFF9C0929080",
-10597 => x"C0C0BFF9C09290F8",
-10596 => x"C0C0BFF9C0929082",
-10595 => x"C0C0BFF9C0929092",
-10594 => x"C0C0BFF9C0929099",
-10593 => x"C0C0BFF9C09290B0",
-10592 => x"C0C0BFF9C09290A4",
-10591 => x"C0C0BFF9C09290F9",
-10590 => x"C0C0BFF9C09290C0",
-10589 => x"C0C0BFF9C0928090",
-10588 => x"C0C0BFF9C0928080",
-10587 => x"C0C0BFF9C09280F8",
-10586 => x"C0C0BFF9C0928082",
-10585 => x"C0C0BFF9C0928092",
-10584 => x"C0C0BFF9C0928099",
-10583 => x"C0C0BFF9C09280B0",
-10582 => x"C0C0BFF9C09280A4",
-10581 => x"C0C0BFF9C09280F9",
-10580 => x"C0C0BFF9C09280C0",
-10579 => x"C0C0BFF9C092F890",
-10578 => x"C0C0BFF9C092F880",
-10577 => x"C0C0BFF9C092F8F8",
-10576 => x"C0C0BFF9C092F882",
-10575 => x"C0C0BFF9C092F892",
-10574 => x"C0C0BFF9C092F899",
-10573 => x"C0C0BFF9C092F8B0",
-10572 => x"C0C0BFF9C092F8A4",
-10571 => x"C0C0BFF9C092F8F9",
-10570 => x"C0C0BFF9C092F8C0",
-10569 => x"C0C0BFF9C0928290",
-10568 => x"C0C0BFF9C0928280",
-10567 => x"C0C0BFF9C09282F8",
-10566 => x"C0C0BFF9C0928282",
-10565 => x"C0C0BFF9C0928292",
-10564 => x"C0C0BFF9C0928299",
-10563 => x"C0C0BFF9C09282B0",
-10562 => x"C0C0BFF9C09282A4",
-10561 => x"C0C0BFF9C09282F9",
-10560 => x"C0C0BFF9C09282C0",
-10559 => x"C0C0BFF9C0929290",
-10558 => x"C0C0BFF9C0929280",
-10557 => x"C0C0BFF9C09292F8",
-10556 => x"C0C0BFF9C0929282",
-10555 => x"C0C0BFF9C0929292",
-10554 => x"C0C0BFF9C0929299",
-10553 => x"C0C0BFF9C09292B0",
-10552 => x"C0C0BFF9C09292A4",
-10551 => x"C0C0BFF9C09292F9",
-10550 => x"C0C0BFF9C09292C0",
-10549 => x"C0C0BFF9C0929990",
-10548 => x"C0C0BFF9C0929980",
-10547 => x"C0C0BFF9C09299F8",
-10546 => x"C0C0BFF9C0929982",
-10545 => x"C0C0BFF9C0929992",
-10544 => x"C0C0BFF9C0929999",
-10543 => x"C0C0BFF9C09299B0",
-10542 => x"C0C0BFF9C09299A4",
-10541 => x"C0C0BFF9C09299F9",
-10540 => x"C0C0BFF9C09299C0",
-10539 => x"C0C0BFF9C092B090",
-10538 => x"C0C0BFF9C092B080",
-10537 => x"C0C0BFF9C092B0F8",
-10536 => x"C0C0BFF9C092B082",
-10535 => x"C0C0BFF9C092B092",
-10534 => x"C0C0BFF9C092B099",
-10533 => x"C0C0BFF9C092B0B0",
-10532 => x"C0C0BFF9C092B0A4",
-10531 => x"C0C0BFF9C092B0F9",
-10530 => x"C0C0BFF9C092B0C0",
-10529 => x"C0C0BFF9C092A490",
-10528 => x"C0C0BFF9C092A480",
-10527 => x"C0C0BFF9C092A4F8",
-10526 => x"C0C0BFF9C092A482",
-10525 => x"C0C0BFF9C092A492",
-10524 => x"C0C0BFF9C092A499",
-10523 => x"C0C0BFF9C092A4B0",
-10522 => x"C0C0BFF9C092A4A4",
-10521 => x"C0C0BFF9C092A4F9",
-10520 => x"C0C0BFF9C092A4C0",
-10519 => x"C0C0BFF9C092F990",
-10518 => x"C0C0BFF9C092F980",
-10517 => x"C0C0BFF9C092F9F8",
-10516 => x"C0C0BFF9C092F982",
-10515 => x"C0C0BFF9C092F992",
-10514 => x"C0C0BFF9C092F999",
-10513 => x"C0C0BFF9C092F9B0",
-10512 => x"C0C0BFF9C092F9A4",
-10511 => x"C0C0BFF9C092F9F9",
-10510 => x"C0C0BFF9C092F9C0",
-10509 => x"C0C0BFF9C092C090",
-10508 => x"C0C0BFF9C092C080",
-10507 => x"C0C0BFF9C092C0F8",
-10506 => x"C0C0BFF9C092C082",
-10505 => x"C0C0BFF9C092C092",
-10504 => x"C0C0BFF9C092C099",
-10503 => x"C0C0BFF9C092C0B0",
-10502 => x"C0C0BFF9C092C0A4",
-10501 => x"C0C0BFF9C092C0F9",
-10500 => x"C0C0BFF9C092C0C0",
-10499 => x"C0C0BFF9C0999090",
-10498 => x"C0C0BFF9C0999080",
-10497 => x"C0C0BFF9C09990F8",
-10496 => x"C0C0BFF9C0999082",
-10495 => x"C0C0BFF9C0999092",
-10494 => x"C0C0BFF9C0999099",
-10493 => x"C0C0BFF9C09990B0",
-10492 => x"C0C0BFF9C09990A4",
-10491 => x"C0C0BFF9C09990F9",
-10490 => x"C0C0BFF9C09990C0",
-10489 => x"C0C0BFF9C0998090",
-10488 => x"C0C0BFF9C0998080",
-10487 => x"C0C0BFF9C09980F8",
-10486 => x"C0C0BFF9C0998082",
-10485 => x"C0C0BFF9C0998092",
-10484 => x"C0C0BFF9C0998099",
-10483 => x"C0C0BFF9C09980B0",
-10482 => x"C0C0BFF9C09980A4",
-10481 => x"C0C0BFF9C09980F9",
-10480 => x"C0C0BFF9C09980C0",
-10479 => x"C0C0BFF9C099F890",
-10478 => x"C0C0BFF9C099F880",
-10477 => x"C0C0BFF9C099F8F8",
-10476 => x"C0C0BFF9C099F882",
-10475 => x"C0C0BFF9C099F892",
-10474 => x"C0C0BFF9C099F899",
-10473 => x"C0C0BFF9C099F8B0",
-10472 => x"C0C0BFF9C099F8A4",
-10471 => x"C0C0BFF9C099F8F9",
-10470 => x"C0C0BFF9C099F8C0",
-10469 => x"C0C0BFF9C0998290",
-10468 => x"C0C0BFF9C0998280",
-10467 => x"C0C0BFF9C09982F8",
-10466 => x"C0C0BFF9C0998282",
-10465 => x"C0C0BFF9C0998292",
-10464 => x"C0C0BFF9C0998299",
-10463 => x"C0C0BFF9C09982B0",
-10462 => x"C0C0BFF9C09982A4",
-10461 => x"C0C0BFF9C09982F9",
-10460 => x"C0C0BFF9C09982C0",
-10459 => x"C0C0BFF9C0999290",
-10458 => x"C0C0BFF9C0999280",
-10457 => x"C0C0BFF9C09992F8",
-10456 => x"C0C0BFF9C0999282",
-10455 => x"C0C0BFF9C0999292",
-10454 => x"C0C0BFF9C0999299",
-10453 => x"C0C0BFF9C09992B0",
-10452 => x"C0C0BFF9C09992A4",
-10451 => x"C0C0BFF9C09992F9",
-10450 => x"C0C0BFF9C09992C0",
-10449 => x"C0C0BFF9C0999990",
-10448 => x"C0C0BFF9C0999980",
-10447 => x"C0C0BFF9C09999F8",
-10446 => x"C0C0BFF9C0999982",
-10445 => x"C0C0BFF9C0999992",
-10444 => x"C0C0BFF9C0999999",
-10443 => x"C0C0BFF9C09999B0",
-10442 => x"C0C0BFF9C09999A4",
-10441 => x"C0C0BFF9C09999F9",
-10440 => x"C0C0BFF9C09999C0",
-10439 => x"C0C0BFF9C099B090",
-10438 => x"C0C0BFF9C099B080",
-10437 => x"C0C0BFF9C099B0F8",
-10436 => x"C0C0BFF9C099B082",
-10435 => x"C0C0BFF9C099B092",
-10434 => x"C0C0BFF9C099B099",
-10433 => x"C0C0BFF9C099B0B0",
-10432 => x"C0C0BFF9C099B0A4",
-10431 => x"C0C0BFF9C099B0F9",
-10430 => x"C0C0BFF9C099B0C0",
-10429 => x"C0C0BFF9C099A490",
-10428 => x"C0C0BFF9C099A480",
-10427 => x"C0C0BFF9C099A4F8",
-10426 => x"C0C0BFF9C099A482",
-10425 => x"C0C0BFF9C099A492",
-10424 => x"C0C0BFF9C099A499",
-10423 => x"C0C0BFF9C099A4B0",
-10422 => x"C0C0BFF9C099A4A4",
-10421 => x"C0C0BFF9C099A4F9",
-10420 => x"C0C0BFF9C099A4C0",
-10419 => x"C0C0BFF9C099F990",
-10418 => x"C0C0BFF9C099F980",
-10417 => x"C0C0BFF9C099F9F8",
-10416 => x"C0C0BFF9C099F982",
-10415 => x"C0C0BFF9C099F992",
-10414 => x"C0C0BFF9C099F999",
-10413 => x"C0C0BFF9C099F9B0",
-10412 => x"C0C0BFF9C099F9A4",
-10411 => x"C0C0BFF9C099F9F9",
-10410 => x"C0C0BFF9C099F9C0",
-10409 => x"C0C0BFF9C099C090",
-10408 => x"C0C0BFF9C099C080",
-10407 => x"C0C0BFF9C099C0F8",
-10406 => x"C0C0BFF9C099C082",
-10405 => x"C0C0BFF9C099C092",
-10404 => x"C0C0BFF9C099C099",
-10403 => x"C0C0BFF9C099C0B0",
-10402 => x"C0C0BFF9C099C0A4",
-10401 => x"C0C0BFF9C099C0F9",
-10400 => x"C0C0BFF9C099C0C0",
-10399 => x"C0C0BFF9C0B09090",
-10398 => x"C0C0BFF9C0B09080",
-10397 => x"C0C0BFF9C0B090F8",
-10396 => x"C0C0BFF9C0B09082",
-10395 => x"C0C0BFF9C0B09092",
-10394 => x"C0C0BFF9C0B09099",
-10393 => x"C0C0BFF9C0B090B0",
-10392 => x"C0C0BFF9C0B090A4",
-10391 => x"C0C0BFF9C0B090F9",
-10390 => x"C0C0BFF9C0B090C0",
-10389 => x"C0C0BFF9C0B08090",
-10388 => x"C0C0BFF9C0B08080",
-10387 => x"C0C0BFF9C0B080F8",
-10386 => x"C0C0BFF9C0B08082",
-10385 => x"C0C0BFF9C0B08092",
-10384 => x"C0C0BFF9C0B08099",
-10383 => x"C0C0BFF9C0B080B0",
-10382 => x"C0C0BFF9C0B080A4",
-10381 => x"C0C0BFF9C0B080F9",
-10380 => x"C0C0BFF9C0B080C0",
-10379 => x"C0C0BFF9C0B0F890",
-10378 => x"C0C0BFF9C0B0F880",
-10377 => x"C0C0BFF9C0B0F8F8",
-10376 => x"C0C0BFF9C0B0F882",
-10375 => x"C0C0BFF9C0B0F892",
-10374 => x"C0C0BFF9C0B0F899",
-10373 => x"C0C0BFF9C0B0F8B0",
-10372 => x"C0C0BFF9C0B0F8A4",
-10371 => x"C0C0BFF9C0B0F8F9",
-10370 => x"C0C0BFF9C0B0F8C0",
-10369 => x"C0C0BFF9C0B08290",
-10368 => x"C0C0BFF9C0B08280",
-10367 => x"C0C0BFF9C0B082F8",
-10366 => x"C0C0BFF9C0B08282",
-10365 => x"C0C0BFF9C0B08292",
-10364 => x"C0C0BFF9C0B08299",
-10363 => x"C0C0BFF9C0B082B0",
-10362 => x"C0C0BFF9C0B082A4",
-10361 => x"C0C0BFF9C0B082F9",
-10360 => x"C0C0BFF9C0B082C0",
-10359 => x"C0C0BFF9C0B09290",
-10358 => x"C0C0BFF9C0B09280",
-10357 => x"C0C0BFF9C0B092F8",
-10356 => x"C0C0BFF9C0B09282",
-10355 => x"C0C0BFF9C0B09292",
-10354 => x"C0C0BFF9C0B09299",
-10353 => x"C0C0BFF9C0B092B0",
-10352 => x"C0C0BFF9C0B092A4",
-10351 => x"C0C0BFF9C0B092F9",
-10350 => x"C0C0BFF9C0B092C0",
-10349 => x"C0C0BFF9C0B09990",
-10348 => x"C0C0BFF9C0B09980",
-10347 => x"C0C0BFF9C0B099F8",
-10346 => x"C0C0BFF9C0B09982",
-10345 => x"C0C0BFF9C0B09992",
-10344 => x"C0C0BFF9C0B09999",
-10343 => x"C0C0BFF9C0B099B0",
-10342 => x"C0C0BFF9C0B099A4",
-10341 => x"C0C0BFF9C0B099F9",
-10340 => x"C0C0BFF9C0B099C0",
-10339 => x"C0C0BFF9C0B0B090",
-10338 => x"C0C0BFF9C0B0B080",
-10337 => x"C0C0BFF9C0B0B0F8",
-10336 => x"C0C0BFF9C0B0B082",
-10335 => x"C0C0BFF9C0B0B092",
-10334 => x"C0C0BFF9C0B0B099",
-10333 => x"C0C0BFF9C0B0B0B0",
-10332 => x"C0C0BFF9C0B0B0A4",
-10331 => x"C0C0BFF9C0B0B0F9",
-10330 => x"C0C0BFF9C0B0B0C0",
-10329 => x"C0C0BFF9C0B0A490",
-10328 => x"C0C0BFF9C0B0A480",
-10327 => x"C0C0BFF9C0B0A4F8",
-10326 => x"C0C0BFF9C0B0A482",
-10325 => x"C0C0BFF9C0B0A492",
-10324 => x"C0C0BFF9C0B0A499",
-10323 => x"C0C0BFF9C0B0A4B0",
-10322 => x"C0C0BFF9C0B0A4A4",
-10321 => x"C0C0BFF9C0B0A4F9",
-10320 => x"C0C0BFF9C0B0A4C0",
-10319 => x"C0C0BFF9C0B0F990",
-10318 => x"C0C0BFF9C0B0F980",
-10317 => x"C0C0BFF9C0B0F9F8",
-10316 => x"C0C0BFF9C0B0F982",
-10315 => x"C0C0BFF9C0B0F992",
-10314 => x"C0C0BFF9C0B0F999",
-10313 => x"C0C0BFF9C0B0F9B0",
-10312 => x"C0C0BFF9C0B0F9A4",
-10311 => x"C0C0BFF9C0B0F9F9",
-10310 => x"C0C0BFF9C0B0F9C0",
-10309 => x"C0C0BFF9C0B0C090",
-10308 => x"C0C0BFF9C0B0C080",
-10307 => x"C0C0BFF9C0B0C0F8",
-10306 => x"C0C0BFF9C0B0C082",
-10305 => x"C0C0BFF9C0B0C092",
-10304 => x"C0C0BFF9C0B0C099",
-10303 => x"C0C0BFF9C0B0C0B0",
-10302 => x"C0C0BFF9C0B0C0A4",
-10301 => x"C0C0BFF9C0B0C0F9",
-10300 => x"C0C0BFF9C0B0C0C0",
-10299 => x"C0C0BFF9C0A49090",
-10298 => x"C0C0BFF9C0A49080",
-10297 => x"C0C0BFF9C0A490F8",
-10296 => x"C0C0BFF9C0A49082",
-10295 => x"C0C0BFF9C0A49092",
-10294 => x"C0C0BFF9C0A49099",
-10293 => x"C0C0BFF9C0A490B0",
-10292 => x"C0C0BFF9C0A490A4",
-10291 => x"C0C0BFF9C0A490F9",
-10290 => x"C0C0BFF9C0A490C0",
-10289 => x"C0C0BFF9C0A48090",
-10288 => x"C0C0BFF9C0A48080",
-10287 => x"C0C0BFF9C0A480F8",
-10286 => x"C0C0BFF9C0A48082",
-10285 => x"C0C0BFF9C0A48092",
-10284 => x"C0C0BFF9C0A48099",
-10283 => x"C0C0BFF9C0A480B0",
-10282 => x"C0C0BFF9C0A480A4",
-10281 => x"C0C0BFF9C0A480F9",
-10280 => x"C0C0BFF9C0A480C0",
-10279 => x"C0C0BFF9C0A4F890",
-10278 => x"C0C0BFF9C0A4F880",
-10277 => x"C0C0BFF9C0A4F8F8",
-10276 => x"C0C0BFF9C0A4F882",
-10275 => x"C0C0BFF9C0A4F892",
-10274 => x"C0C0BFF9C0A4F899",
-10273 => x"C0C0BFF9C0A4F8B0",
-10272 => x"C0C0BFF9C0A4F8A4",
-10271 => x"C0C0BFF9C0A4F8F9",
-10270 => x"C0C0BFF9C0A4F8C0",
-10269 => x"C0C0BFF9C0A48290",
-10268 => x"C0C0BFF9C0A48280",
-10267 => x"C0C0BFF9C0A482F8",
-10266 => x"C0C0BFF9C0A48282",
-10265 => x"C0C0BFF9C0A48292",
-10264 => x"C0C0BFF9C0A48299",
-10263 => x"C0C0BFF9C0A482B0",
-10262 => x"C0C0BFF9C0A482A4",
-10261 => x"C0C0BFF9C0A482F9",
-10260 => x"C0C0BFF9C0A482C0",
-10259 => x"C0C0BFF9C0A49290",
-10258 => x"C0C0BFF9C0A49280",
-10257 => x"C0C0BFF9C0A492F8",
-10256 => x"C0C0BFF9C0A49282",
-10255 => x"C0C0BFF9C0A49292",
-10254 => x"C0C0BFF9C0A49299",
-10253 => x"C0C0BFF9C0A492B0",
-10252 => x"C0C0BFF9C0A492A4",
-10251 => x"C0C0BFF9C0A492F9",
-10250 => x"C0C0BFF9C0A492C0",
-10249 => x"C0C0BFF9C0A49990",
-10248 => x"C0C0BFF9C0A49980",
-10247 => x"C0C0BFF9C0A499F8",
-10246 => x"C0C0BFF9C0A49982",
-10245 => x"C0C0BFF9C0A49992",
-10244 => x"C0C0BFF9C0A49999",
-10243 => x"C0C0BFF9C0A499B0",
-10242 => x"C0C0BFF9C0A499A4",
-10241 => x"C0C0BFF9C0A499F9",
-10240 => x"C0C0BFF9C0A499C0",
-10239 => x"C0C0BFF9C0A4B090",
-10238 => x"C0C0BFF9C0A4B080",
-10237 => x"C0C0BFF9C0A4B0F8",
-10236 => x"C0C0BFF9C0A4B082",
-10235 => x"C0C0BFF9C0A4B092",
-10234 => x"C0C0BFF9C0A4B099",
-10233 => x"C0C0BFF9C0A4B0B0",
-10232 => x"C0C0BFF9C0A4B0A4",
-10231 => x"C0C0BFF9C0A4B0F9",
-10230 => x"C0C0BFF9C0A4B0C0",
-10229 => x"C0C0BFF9C0A4A490",
-10228 => x"C0C0BFF9C0A4A480",
-10227 => x"C0C0BFF9C0A4A4F8",
-10226 => x"C0C0BFF9C0A4A482",
-10225 => x"C0C0BFF9C0A4A492",
-10224 => x"C0C0BFF9C0A4A499",
-10223 => x"C0C0BFF9C0A4A4B0",
-10222 => x"C0C0BFF9C0A4A4A4",
-10221 => x"C0C0BFF9C0A4A4F9",
-10220 => x"C0C0BFF9C0A4A4C0",
-10219 => x"C0C0BFF9C0A4F990",
-10218 => x"C0C0BFF9C0A4F980",
-10217 => x"C0C0BFF9C0A4F9F8",
-10216 => x"C0C0BFF9C0A4F982",
-10215 => x"C0C0BFF9C0A4F992",
-10214 => x"C0C0BFF9C0A4F999",
-10213 => x"C0C0BFF9C0A4F9B0",
-10212 => x"C0C0BFF9C0A4F9A4",
-10211 => x"C0C0BFF9C0A4F9F9",
-10210 => x"C0C0BFF9C0A4F9C0",
-10209 => x"C0C0BFF9C0A4C090",
-10208 => x"C0C0BFF9C0A4C080",
-10207 => x"C0C0BFF9C0A4C0F8",
-10206 => x"C0C0BFF9C0A4C082",
-10205 => x"C0C0BFF9C0A4C092",
-10204 => x"C0C0BFF9C0A4C099",
-10203 => x"C0C0BFF9C0A4C0B0",
-10202 => x"C0C0BFF9C0A4C0A4",
-10201 => x"C0C0BFF9C0A4C0F9",
-10200 => x"C0C0BFF9C0A4C0C0",
-10199 => x"C0C0BFF9C0F99090",
-10198 => x"C0C0BFF9C0F99080",
-10197 => x"C0C0BFF9C0F990F8",
-10196 => x"C0C0BFF9C0F99082",
-10195 => x"C0C0BFF9C0F99092",
-10194 => x"C0C0BFF9C0F99099",
-10193 => x"C0C0BFF9C0F990B0",
-10192 => x"C0C0BFF9C0F990A4",
-10191 => x"C0C0BFF9C0F990F9",
-10190 => x"C0C0BFF9C0F990C0",
-10189 => x"C0C0BFF9C0F98090",
-10188 => x"C0C0BFF9C0F98080",
-10187 => x"C0C0BFF9C0F980F8",
-10186 => x"C0C0BFF9C0F98082",
-10185 => x"C0C0BFF9C0F98092",
-10184 => x"C0C0BFF9C0F98099",
-10183 => x"C0C0BFF9C0F980B0",
-10182 => x"C0C0BFF9C0F980A4",
-10181 => x"C0C0BFF9C0F980F9",
-10180 => x"C0C0BFF9C0F980C0",
-10179 => x"C0C0BFF9C0F9F890",
-10178 => x"C0C0BFF9C0F9F880",
-10177 => x"C0C0BFF9C0F9F8F8",
-10176 => x"C0C0BFF9C0F9F882",
-10175 => x"C0C0BFF9C0F9F892",
-10174 => x"C0C0BFF9C0F9F899",
-10173 => x"C0C0BFF9C0F9F8B0",
-10172 => x"C0C0BFF9C0F9F8A4",
-10171 => x"C0C0BFF9C0F9F8F9",
-10170 => x"C0C0BFF9C0F9F8C0",
-10169 => x"C0C0BFF9C0F98290",
-10168 => x"C0C0BFF9C0F98280",
-10167 => x"C0C0BFF9C0F982F8",
-10166 => x"C0C0BFF9C0F98282",
-10165 => x"C0C0BFF9C0F98292",
-10164 => x"C0C0BFF9C0F98299",
-10163 => x"C0C0BFF9C0F982B0",
-10162 => x"C0C0BFF9C0F982A4",
-10161 => x"C0C0BFF9C0F982F9",
-10160 => x"C0C0BFF9C0F982C0",
-10159 => x"C0C0BFF9C0F99290",
-10158 => x"C0C0BFF9C0F99280",
-10157 => x"C0C0BFF9C0F992F8",
-10156 => x"C0C0BFF9C0F99282",
-10155 => x"C0C0BFF9C0F99292",
-10154 => x"C0C0BFF9C0F99299",
-10153 => x"C0C0BFF9C0F992B0",
-10152 => x"C0C0BFF9C0F992A4",
-10151 => x"C0C0BFF9C0F992F9",
-10150 => x"C0C0BFF9C0F992C0",
-10149 => x"C0C0BFF9C0F99990",
-10148 => x"C0C0BFF9C0F99980",
-10147 => x"C0C0BFF9C0F999F8",
-10146 => x"C0C0BFF9C0F99982",
-10145 => x"C0C0BFF9C0F99992",
-10144 => x"C0C0BFF9C0F99999",
-10143 => x"C0C0BFF9C0F999B0",
-10142 => x"C0C0BFF9C0F999A4",
-10141 => x"C0C0BFF9C0F999F9",
-10140 => x"C0C0BFF9C0F999C0",
-10139 => x"C0C0BFF9C0F9B090",
-10138 => x"C0C0BFF9C0F9B080",
-10137 => x"C0C0BFF9C0F9B0F8",
-10136 => x"C0C0BFF9C0F9B082",
-10135 => x"C0C0BFF9C0F9B092",
-10134 => x"C0C0BFF9C0F9B099",
-10133 => x"C0C0BFF9C0F9B0B0",
-10132 => x"C0C0BFF9C0F9B0A4",
-10131 => x"C0C0BFF9C0F9B0F9",
-10130 => x"C0C0BFF9C0F9B0C0",
-10129 => x"C0C0BFF9C0F9A490",
-10128 => x"C0C0BFF9C0F9A480",
-10127 => x"C0C0BFF9C0F9A4F8",
-10126 => x"C0C0BFF9C0F9A482",
-10125 => x"C0C0BFF9C0F9A492",
-10124 => x"C0C0BFF9C0F9A499",
-10123 => x"C0C0BFF9C0F9A4B0",
-10122 => x"C0C0BFF9C0F9A4A4",
-10121 => x"C0C0BFF9C0F9A4F9",
-10120 => x"C0C0BFF9C0F9A4C0",
-10119 => x"C0C0BFF9C0F9F990",
-10118 => x"C0C0BFF9C0F9F980",
-10117 => x"C0C0BFF9C0F9F9F8",
-10116 => x"C0C0BFF9C0F9F982",
-10115 => x"C0C0BFF9C0F9F992",
-10114 => x"C0C0BFF9C0F9F999",
-10113 => x"C0C0BFF9C0F9F9B0",
-10112 => x"C0C0BFF9C0F9F9A4",
-10111 => x"C0C0BFF9C0F9F9F9",
-10110 => x"C0C0BFF9C0F9F9C0",
-10109 => x"C0C0BFF9C0F9C090",
-10108 => x"C0C0BFF9C0F9C080",
-10107 => x"C0C0BFF9C0F9C0F8",
-10106 => x"C0C0BFF9C0F9C082",
-10105 => x"C0C0BFF9C0F9C092",
-10104 => x"C0C0BFF9C0F9C099",
-10103 => x"C0C0BFF9C0F9C0B0",
-10102 => x"C0C0BFF9C0F9C0A4",
-10101 => x"C0C0BFF9C0F9C0F9",
-10100 => x"C0C0BFF9C0F9C0C0",
-10099 => x"C0C0BFF9C0C09090",
-10098 => x"C0C0BFF9C0C09080",
-10097 => x"C0C0BFF9C0C090F8",
-10096 => x"C0C0BFF9C0C09082",
-10095 => x"C0C0BFF9C0C09092",
-10094 => x"C0C0BFF9C0C09099",
-10093 => x"C0C0BFF9C0C090B0",
-10092 => x"C0C0BFF9C0C090A4",
-10091 => x"C0C0BFF9C0C090F9",
-10090 => x"C0C0BFF9C0C090C0",
-10089 => x"C0C0BFF9C0C08090",
-10088 => x"C0C0BFF9C0C08080",
-10087 => x"C0C0BFF9C0C080F8",
-10086 => x"C0C0BFF9C0C08082",
-10085 => x"C0C0BFF9C0C08092",
-10084 => x"C0C0BFF9C0C08099",
-10083 => x"C0C0BFF9C0C080B0",
-10082 => x"C0C0BFF9C0C080A4",
-10081 => x"C0C0BFF9C0C080F9",
-10080 => x"C0C0BFF9C0C080C0",
-10079 => x"C0C0BFF9C0C0F890",
-10078 => x"C0C0BFF9C0C0F880",
-10077 => x"C0C0BFF9C0C0F8F8",
-10076 => x"C0C0BFF9C0C0F882",
-10075 => x"C0C0BFF9C0C0F892",
-10074 => x"C0C0BFF9C0C0F899",
-10073 => x"C0C0BFF9C0C0F8B0",
-10072 => x"C0C0BFF9C0C0F8A4",
-10071 => x"C0C0BFF9C0C0F8F9",
-10070 => x"C0C0BFF9C0C0F8C0",
-10069 => x"C0C0BFF9C0C08290",
-10068 => x"C0C0BFF9C0C08280",
-10067 => x"C0C0BFF9C0C082F8",
-10066 => x"C0C0BFF9C0C08282",
-10065 => x"C0C0BFF9C0C08292",
-10064 => x"C0C0BFF9C0C08299",
-10063 => x"C0C0BFF9C0C082B0",
-10062 => x"C0C0BFF9C0C082A4",
-10061 => x"C0C0BFF9C0C082F9",
-10060 => x"C0C0BFF9C0C082C0",
-10059 => x"C0C0BFF9C0C09290",
-10058 => x"C0C0BFF9C0C09280",
-10057 => x"C0C0BFF9C0C092F8",
-10056 => x"C0C0BFF9C0C09282",
-10055 => x"C0C0BFF9C0C09292",
-10054 => x"C0C0BFF9C0C09299",
-10053 => x"C0C0BFF9C0C092B0",
-10052 => x"C0C0BFF9C0C092A4",
-10051 => x"C0C0BFF9C0C092F9",
-10050 => x"C0C0BFF9C0C092C0",
-10049 => x"C0C0BFF9C0C09990",
-10048 => x"C0C0BFF9C0C09980",
-10047 => x"C0C0BFF9C0C099F8",
-10046 => x"C0C0BFF9C0C09982",
-10045 => x"C0C0BFF9C0C09992",
-10044 => x"C0C0BFF9C0C09999",
-10043 => x"C0C0BFF9C0C099B0",
-10042 => x"C0C0BFF9C0C099A4",
-10041 => x"C0C0BFF9C0C099F9",
-10040 => x"C0C0BFF9C0C099C0",
-10039 => x"C0C0BFF9C0C0B090",
-10038 => x"C0C0BFF9C0C0B080",
-10037 => x"C0C0BFF9C0C0B0F8",
-10036 => x"C0C0BFF9C0C0B082",
-10035 => x"C0C0BFF9C0C0B092",
-10034 => x"C0C0BFF9C0C0B099",
-10033 => x"C0C0BFF9C0C0B0B0",
-10032 => x"C0C0BFF9C0C0B0A4",
-10031 => x"C0C0BFF9C0C0B0F9",
-10030 => x"C0C0BFF9C0C0B0C0",
-10029 => x"C0C0BFF9C0C0A490",
-10028 => x"C0C0BFF9C0C0A480",
-10027 => x"C0C0BFF9C0C0A4F8",
-10026 => x"C0C0BFF9C0C0A482",
-10025 => x"C0C0BFF9C0C0A492",
-10024 => x"C0C0BFF9C0C0A499",
-10023 => x"C0C0BFF9C0C0A4B0",
-10022 => x"C0C0BFF9C0C0A4A4",
-10021 => x"C0C0BFF9C0C0A4F9",
-10020 => x"C0C0BFF9C0C0A4C0",
-10019 => x"C0C0BFF9C0C0F990",
-10018 => x"C0C0BFF9C0C0F980",
-10017 => x"C0C0BFF9C0C0F9F8",
-10016 => x"C0C0BFF9C0C0F982",
-10015 => x"C0C0BFF9C0C0F992",
-10014 => x"C0C0BFF9C0C0F999",
-10013 => x"C0C0BFF9C0C0F9B0",
-10012 => x"C0C0BFF9C0C0F9A4",
-10011 => x"C0C0BFF9C0C0F9F9",
-10010 => x"C0C0BFF9C0C0F9C0",
-10009 => x"C0C0BFF9C0C0C090",
-10008 => x"C0C0BFF9C0C0C080",
-10007 => x"C0C0BFF9C0C0C0F8",
-10006 => x"C0C0BFF9C0C0C082",
-10005 => x"C0C0BFF9C0C0C092",
-10004 => x"C0C0BFF9C0C0C099",
-10003 => x"C0C0BFF9C0C0C0B0",
-10002 => x"C0C0BFF9C0C0C0A4",
-10001 => x"C0C0BFF9C0C0C0F9",
-10000 => x"C0C0BFF9C0C0C0C0",
 -9999 => x"C0C0C0BF90909090",
 -9998 => x"C0C0C0BF90909080",
 -9997 => x"C0C0C0BF909090F8",
 -9996 => x"C0C0C0BF90909082",
 -9995 => x"C0C0C0BF90909092",
 -9994 => x"C0C0C0BF90909099",
 -9993 => x"C0C0C0BF909090B0",
 -9992 => x"C0C0C0BF909090A4",
 -9991 => x"C0C0C0BF909090F9",
 -9990 => x"C0C0C0BF909090C0",
 -9989 => x"C0C0C0BF90908090",
 -9988 => x"C0C0C0BF90908080",
 -9987 => x"C0C0C0BF909080F8",
 -9986 => x"C0C0C0BF90908082",
 -9985 => x"C0C0C0BF90908092",
 -9984 => x"C0C0C0BF90908099",
 -9983 => x"C0C0C0BF909080B0",
 -9982 => x"C0C0C0BF909080A4",
 -9981 => x"C0C0C0BF909080F9",
 -9980 => x"C0C0C0BF909080C0",
 -9979 => x"C0C0C0BF9090F890",
 -9978 => x"C0C0C0BF9090F880",
 -9977 => x"C0C0C0BF9090F8F8",
 -9976 => x"C0C0C0BF9090F882",
 -9975 => x"C0C0C0BF9090F892",
 -9974 => x"C0C0C0BF9090F899",
 -9973 => x"C0C0C0BF9090F8B0",
 -9972 => x"C0C0C0BF9090F8A4",
 -9971 => x"C0C0C0BF9090F8F9",
 -9970 => x"C0C0C0BF9090F8C0",
 -9969 => x"C0C0C0BF90908290",
 -9968 => x"C0C0C0BF90908280",
 -9967 => x"C0C0C0BF909082F8",
 -9966 => x"C0C0C0BF90908282",
 -9965 => x"C0C0C0BF90908292",
 -9964 => x"C0C0C0BF90908299",
 -9963 => x"C0C0C0BF909082B0",
 -9962 => x"C0C0C0BF909082A4",
 -9961 => x"C0C0C0BF909082F9",
 -9960 => x"C0C0C0BF909082C0",
 -9959 => x"C0C0C0BF90909290",
 -9958 => x"C0C0C0BF90909280",
 -9957 => x"C0C0C0BF909092F8",
 -9956 => x"C0C0C0BF90909282",
 -9955 => x"C0C0C0BF90909292",
 -9954 => x"C0C0C0BF90909299",
 -9953 => x"C0C0C0BF909092B0",
 -9952 => x"C0C0C0BF909092A4",
 -9951 => x"C0C0C0BF909092F9",
 -9950 => x"C0C0C0BF909092C0",
 -9949 => x"C0C0C0BF90909990",
 -9948 => x"C0C0C0BF90909980",
 -9947 => x"C0C0C0BF909099F8",
 -9946 => x"C0C0C0BF90909982",
 -9945 => x"C0C0C0BF90909992",
 -9944 => x"C0C0C0BF90909999",
 -9943 => x"C0C0C0BF909099B0",
 -9942 => x"C0C0C0BF909099A4",
 -9941 => x"C0C0C0BF909099F9",
 -9940 => x"C0C0C0BF909099C0",
 -9939 => x"C0C0C0BF9090B090",
 -9938 => x"C0C0C0BF9090B080",
 -9937 => x"C0C0C0BF9090B0F8",
 -9936 => x"C0C0C0BF9090B082",
 -9935 => x"C0C0C0BF9090B092",
 -9934 => x"C0C0C0BF9090B099",
 -9933 => x"C0C0C0BF9090B0B0",
 -9932 => x"C0C0C0BF9090B0A4",
 -9931 => x"C0C0C0BF9090B0F9",
 -9930 => x"C0C0C0BF9090B0C0",
 -9929 => x"C0C0C0BF9090A490",
 -9928 => x"C0C0C0BF9090A480",
 -9927 => x"C0C0C0BF9090A4F8",
 -9926 => x"C0C0C0BF9090A482",
 -9925 => x"C0C0C0BF9090A492",
 -9924 => x"C0C0C0BF9090A499",
 -9923 => x"C0C0C0BF9090A4B0",
 -9922 => x"C0C0C0BF9090A4A4",
 -9921 => x"C0C0C0BF9090A4F9",
 -9920 => x"C0C0C0BF9090A4C0",
 -9919 => x"C0C0C0BF9090F990",
 -9918 => x"C0C0C0BF9090F980",
 -9917 => x"C0C0C0BF9090F9F8",
 -9916 => x"C0C0C0BF9090F982",
 -9915 => x"C0C0C0BF9090F992",
 -9914 => x"C0C0C0BF9090F999",
 -9913 => x"C0C0C0BF9090F9B0",
 -9912 => x"C0C0C0BF9090F9A4",
 -9911 => x"C0C0C0BF9090F9F9",
 -9910 => x"C0C0C0BF9090F9C0",
 -9909 => x"C0C0C0BF9090C090",
 -9908 => x"C0C0C0BF9090C080",
 -9907 => x"C0C0C0BF9090C0F8",
 -9906 => x"C0C0C0BF9090C082",
 -9905 => x"C0C0C0BF9090C092",
 -9904 => x"C0C0C0BF9090C099",
 -9903 => x"C0C0C0BF9090C0B0",
 -9902 => x"C0C0C0BF9090C0A4",
 -9901 => x"C0C0C0BF9090C0F9",
 -9900 => x"C0C0C0BF9090C0C0",
 -9899 => x"C0C0C0BF90809090",
 -9898 => x"C0C0C0BF90809080",
 -9897 => x"C0C0C0BF908090F8",
 -9896 => x"C0C0C0BF90809082",
 -9895 => x"C0C0C0BF90809092",
 -9894 => x"C0C0C0BF90809099",
 -9893 => x"C0C0C0BF908090B0",
 -9892 => x"C0C0C0BF908090A4",
 -9891 => x"C0C0C0BF908090F9",
 -9890 => x"C0C0C0BF908090C0",
 -9889 => x"C0C0C0BF90808090",
 -9888 => x"C0C0C0BF90808080",
 -9887 => x"C0C0C0BF908080F8",
 -9886 => x"C0C0C0BF90808082",
 -9885 => x"C0C0C0BF90808092",
 -9884 => x"C0C0C0BF90808099",
 -9883 => x"C0C0C0BF908080B0",
 -9882 => x"C0C0C0BF908080A4",
 -9881 => x"C0C0C0BF908080F9",
 -9880 => x"C0C0C0BF908080C0",
 -9879 => x"C0C0C0BF9080F890",
 -9878 => x"C0C0C0BF9080F880",
 -9877 => x"C0C0C0BF9080F8F8",
 -9876 => x"C0C0C0BF9080F882",
 -9875 => x"C0C0C0BF9080F892",
 -9874 => x"C0C0C0BF9080F899",
 -9873 => x"C0C0C0BF9080F8B0",
 -9872 => x"C0C0C0BF9080F8A4",
 -9871 => x"C0C0C0BF9080F8F9",
 -9870 => x"C0C0C0BF9080F8C0",
 -9869 => x"C0C0C0BF90808290",
 -9868 => x"C0C0C0BF90808280",
 -9867 => x"C0C0C0BF908082F8",
 -9866 => x"C0C0C0BF90808282",
 -9865 => x"C0C0C0BF90808292",
 -9864 => x"C0C0C0BF90808299",
 -9863 => x"C0C0C0BF908082B0",
 -9862 => x"C0C0C0BF908082A4",
 -9861 => x"C0C0C0BF908082F9",
 -9860 => x"C0C0C0BF908082C0",
 -9859 => x"C0C0C0BF90809290",
 -9858 => x"C0C0C0BF90809280",
 -9857 => x"C0C0C0BF908092F8",
 -9856 => x"C0C0C0BF90809282",
 -9855 => x"C0C0C0BF90809292",
 -9854 => x"C0C0C0BF90809299",
 -9853 => x"C0C0C0BF908092B0",
 -9852 => x"C0C0C0BF908092A4",
 -9851 => x"C0C0C0BF908092F9",
 -9850 => x"C0C0C0BF908092C0",
 -9849 => x"C0C0C0BF90809990",
 -9848 => x"C0C0C0BF90809980",
 -9847 => x"C0C0C0BF908099F8",
 -9846 => x"C0C0C0BF90809982",
 -9845 => x"C0C0C0BF90809992",
 -9844 => x"C0C0C0BF90809999",
 -9843 => x"C0C0C0BF908099B0",
 -9842 => x"C0C0C0BF908099A4",
 -9841 => x"C0C0C0BF908099F9",
 -9840 => x"C0C0C0BF908099C0",
 -9839 => x"C0C0C0BF9080B090",
 -9838 => x"C0C0C0BF9080B080",
 -9837 => x"C0C0C0BF9080B0F8",
 -9836 => x"C0C0C0BF9080B082",
 -9835 => x"C0C0C0BF9080B092",
 -9834 => x"C0C0C0BF9080B099",
 -9833 => x"C0C0C0BF9080B0B0",
 -9832 => x"C0C0C0BF9080B0A4",
 -9831 => x"C0C0C0BF9080B0F9",
 -9830 => x"C0C0C0BF9080B0C0",
 -9829 => x"C0C0C0BF9080A490",
 -9828 => x"C0C0C0BF9080A480",
 -9827 => x"C0C0C0BF9080A4F8",
 -9826 => x"C0C0C0BF9080A482",
 -9825 => x"C0C0C0BF9080A492",
 -9824 => x"C0C0C0BF9080A499",
 -9823 => x"C0C0C0BF9080A4B0",
 -9822 => x"C0C0C0BF9080A4A4",
 -9821 => x"C0C0C0BF9080A4F9",
 -9820 => x"C0C0C0BF9080A4C0",
 -9819 => x"C0C0C0BF9080F990",
 -9818 => x"C0C0C0BF9080F980",
 -9817 => x"C0C0C0BF9080F9F8",
 -9816 => x"C0C0C0BF9080F982",
 -9815 => x"C0C0C0BF9080F992",
 -9814 => x"C0C0C0BF9080F999",
 -9813 => x"C0C0C0BF9080F9B0",
 -9812 => x"C0C0C0BF9080F9A4",
 -9811 => x"C0C0C0BF9080F9F9",
 -9810 => x"C0C0C0BF9080F9C0",
 -9809 => x"C0C0C0BF9080C090",
 -9808 => x"C0C0C0BF9080C080",
 -9807 => x"C0C0C0BF9080C0F8",
 -9806 => x"C0C0C0BF9080C082",
 -9805 => x"C0C0C0BF9080C092",
 -9804 => x"C0C0C0BF9080C099",
 -9803 => x"C0C0C0BF9080C0B0",
 -9802 => x"C0C0C0BF9080C0A4",
 -9801 => x"C0C0C0BF9080C0F9",
 -9800 => x"C0C0C0BF9080C0C0",
 -9799 => x"C0C0C0BF90F89090",
 -9798 => x"C0C0C0BF90F89080",
 -9797 => x"C0C0C0BF90F890F8",
 -9796 => x"C0C0C0BF90F89082",
 -9795 => x"C0C0C0BF90F89092",
 -9794 => x"C0C0C0BF90F89099",
 -9793 => x"C0C0C0BF90F890B0",
 -9792 => x"C0C0C0BF90F890A4",
 -9791 => x"C0C0C0BF90F890F9",
 -9790 => x"C0C0C0BF90F890C0",
 -9789 => x"C0C0C0BF90F88090",
 -9788 => x"C0C0C0BF90F88080",
 -9787 => x"C0C0C0BF90F880F8",
 -9786 => x"C0C0C0BF90F88082",
 -9785 => x"C0C0C0BF90F88092",
 -9784 => x"C0C0C0BF90F88099",
 -9783 => x"C0C0C0BF90F880B0",
 -9782 => x"C0C0C0BF90F880A4",
 -9781 => x"C0C0C0BF90F880F9",
 -9780 => x"C0C0C0BF90F880C0",
 -9779 => x"C0C0C0BF90F8F890",
 -9778 => x"C0C0C0BF90F8F880",
 -9777 => x"C0C0C0BF90F8F8F8",
 -9776 => x"C0C0C0BF90F8F882",
 -9775 => x"C0C0C0BF90F8F892",
 -9774 => x"C0C0C0BF90F8F899",
 -9773 => x"C0C0C0BF90F8F8B0",
 -9772 => x"C0C0C0BF90F8F8A4",
 -9771 => x"C0C0C0BF90F8F8F9",
 -9770 => x"C0C0C0BF90F8F8C0",
 -9769 => x"C0C0C0BF90F88290",
 -9768 => x"C0C0C0BF90F88280",
 -9767 => x"C0C0C0BF90F882F8",
 -9766 => x"C0C0C0BF90F88282",
 -9765 => x"C0C0C0BF90F88292",
 -9764 => x"C0C0C0BF90F88299",
 -9763 => x"C0C0C0BF90F882B0",
 -9762 => x"C0C0C0BF90F882A4",
 -9761 => x"C0C0C0BF90F882F9",
 -9760 => x"C0C0C0BF90F882C0",
 -9759 => x"C0C0C0BF90F89290",
 -9758 => x"C0C0C0BF90F89280",
 -9757 => x"C0C0C0BF90F892F8",
 -9756 => x"C0C0C0BF90F89282",
 -9755 => x"C0C0C0BF90F89292",
 -9754 => x"C0C0C0BF90F89299",
 -9753 => x"C0C0C0BF90F892B0",
 -9752 => x"C0C0C0BF90F892A4",
 -9751 => x"C0C0C0BF90F892F9",
 -9750 => x"C0C0C0BF90F892C0",
 -9749 => x"C0C0C0BF90F89990",
 -9748 => x"C0C0C0BF90F89980",
 -9747 => x"C0C0C0BF90F899F8",
 -9746 => x"C0C0C0BF90F89982",
 -9745 => x"C0C0C0BF90F89992",
 -9744 => x"C0C0C0BF90F89999",
 -9743 => x"C0C0C0BF90F899B0",
 -9742 => x"C0C0C0BF90F899A4",
 -9741 => x"C0C0C0BF90F899F9",
 -9740 => x"C0C0C0BF90F899C0",
 -9739 => x"C0C0C0BF90F8B090",
 -9738 => x"C0C0C0BF90F8B080",
 -9737 => x"C0C0C0BF90F8B0F8",
 -9736 => x"C0C0C0BF90F8B082",
 -9735 => x"C0C0C0BF90F8B092",
 -9734 => x"C0C0C0BF90F8B099",
 -9733 => x"C0C0C0BF90F8B0B0",
 -9732 => x"C0C0C0BF90F8B0A4",
 -9731 => x"C0C0C0BF90F8B0F9",
 -9730 => x"C0C0C0BF90F8B0C0",
 -9729 => x"C0C0C0BF90F8A490",
 -9728 => x"C0C0C0BF90F8A480",
 -9727 => x"C0C0C0BF90F8A4F8",
 -9726 => x"C0C0C0BF90F8A482",
 -9725 => x"C0C0C0BF90F8A492",
 -9724 => x"C0C0C0BF90F8A499",
 -9723 => x"C0C0C0BF90F8A4B0",
 -9722 => x"C0C0C0BF90F8A4A4",
 -9721 => x"C0C0C0BF90F8A4F9",
 -9720 => x"C0C0C0BF90F8A4C0",
 -9719 => x"C0C0C0BF90F8F990",
 -9718 => x"C0C0C0BF90F8F980",
 -9717 => x"C0C0C0BF90F8F9F8",
 -9716 => x"C0C0C0BF90F8F982",
 -9715 => x"C0C0C0BF90F8F992",
 -9714 => x"C0C0C0BF90F8F999",
 -9713 => x"C0C0C0BF90F8F9B0",
 -9712 => x"C0C0C0BF90F8F9A4",
 -9711 => x"C0C0C0BF90F8F9F9",
 -9710 => x"C0C0C0BF90F8F9C0",
 -9709 => x"C0C0C0BF90F8C090",
 -9708 => x"C0C0C0BF90F8C080",
 -9707 => x"C0C0C0BF90F8C0F8",
 -9706 => x"C0C0C0BF90F8C082",
 -9705 => x"C0C0C0BF90F8C092",
 -9704 => x"C0C0C0BF90F8C099",
 -9703 => x"C0C0C0BF90F8C0B0",
 -9702 => x"C0C0C0BF90F8C0A4",
 -9701 => x"C0C0C0BF90F8C0F9",
 -9700 => x"C0C0C0BF90F8C0C0",
 -9699 => x"C0C0C0BF90829090",
 -9698 => x"C0C0C0BF90829080",
 -9697 => x"C0C0C0BF908290F8",
 -9696 => x"C0C0C0BF90829082",
 -9695 => x"C0C0C0BF90829092",
 -9694 => x"C0C0C0BF90829099",
 -9693 => x"C0C0C0BF908290B0",
 -9692 => x"C0C0C0BF908290A4",
 -9691 => x"C0C0C0BF908290F9",
 -9690 => x"C0C0C0BF908290C0",
 -9689 => x"C0C0C0BF90828090",
 -9688 => x"C0C0C0BF90828080",
 -9687 => x"C0C0C0BF908280F8",
 -9686 => x"C0C0C0BF90828082",
 -9685 => x"C0C0C0BF90828092",
 -9684 => x"C0C0C0BF90828099",
 -9683 => x"C0C0C0BF908280B0",
 -9682 => x"C0C0C0BF908280A4",
 -9681 => x"C0C0C0BF908280F9",
 -9680 => x"C0C0C0BF908280C0",
 -9679 => x"C0C0C0BF9082F890",
 -9678 => x"C0C0C0BF9082F880",
 -9677 => x"C0C0C0BF9082F8F8",
 -9676 => x"C0C0C0BF9082F882",
 -9675 => x"C0C0C0BF9082F892",
 -9674 => x"C0C0C0BF9082F899",
 -9673 => x"C0C0C0BF9082F8B0",
 -9672 => x"C0C0C0BF9082F8A4",
 -9671 => x"C0C0C0BF9082F8F9",
 -9670 => x"C0C0C0BF9082F8C0",
 -9669 => x"C0C0C0BF90828290",
 -9668 => x"C0C0C0BF90828280",
 -9667 => x"C0C0C0BF908282F8",
 -9666 => x"C0C0C0BF90828282",
 -9665 => x"C0C0C0BF90828292",
 -9664 => x"C0C0C0BF90828299",
 -9663 => x"C0C0C0BF908282B0",
 -9662 => x"C0C0C0BF908282A4",
 -9661 => x"C0C0C0BF908282F9",
 -9660 => x"C0C0C0BF908282C0",
 -9659 => x"C0C0C0BF90829290",
 -9658 => x"C0C0C0BF90829280",
 -9657 => x"C0C0C0BF908292F8",
 -9656 => x"C0C0C0BF90829282",
 -9655 => x"C0C0C0BF90829292",
 -9654 => x"C0C0C0BF90829299",
 -9653 => x"C0C0C0BF908292B0",
 -9652 => x"C0C0C0BF908292A4",
 -9651 => x"C0C0C0BF908292F9",
 -9650 => x"C0C0C0BF908292C0",
 -9649 => x"C0C0C0BF90829990",
 -9648 => x"C0C0C0BF90829980",
 -9647 => x"C0C0C0BF908299F8",
 -9646 => x"C0C0C0BF90829982",
 -9645 => x"C0C0C0BF90829992",
 -9644 => x"C0C0C0BF90829999",
 -9643 => x"C0C0C0BF908299B0",
 -9642 => x"C0C0C0BF908299A4",
 -9641 => x"C0C0C0BF908299F9",
 -9640 => x"C0C0C0BF908299C0",
 -9639 => x"C0C0C0BF9082B090",
 -9638 => x"C0C0C0BF9082B080",
 -9637 => x"C0C0C0BF9082B0F8",
 -9636 => x"C0C0C0BF9082B082",
 -9635 => x"C0C0C0BF9082B092",
 -9634 => x"C0C0C0BF9082B099",
 -9633 => x"C0C0C0BF9082B0B0",
 -9632 => x"C0C0C0BF9082B0A4",
 -9631 => x"C0C0C0BF9082B0F9",
 -9630 => x"C0C0C0BF9082B0C0",
 -9629 => x"C0C0C0BF9082A490",
 -9628 => x"C0C0C0BF9082A480",
 -9627 => x"C0C0C0BF9082A4F8",
 -9626 => x"C0C0C0BF9082A482",
 -9625 => x"C0C0C0BF9082A492",
 -9624 => x"C0C0C0BF9082A499",
 -9623 => x"C0C0C0BF9082A4B0",
 -9622 => x"C0C0C0BF9082A4A4",
 -9621 => x"C0C0C0BF9082A4F9",
 -9620 => x"C0C0C0BF9082A4C0",
 -9619 => x"C0C0C0BF9082F990",
 -9618 => x"C0C0C0BF9082F980",
 -9617 => x"C0C0C0BF9082F9F8",
 -9616 => x"C0C0C0BF9082F982",
 -9615 => x"C0C0C0BF9082F992",
 -9614 => x"C0C0C0BF9082F999",
 -9613 => x"C0C0C0BF9082F9B0",
 -9612 => x"C0C0C0BF9082F9A4",
 -9611 => x"C0C0C0BF9082F9F9",
 -9610 => x"C0C0C0BF9082F9C0",
 -9609 => x"C0C0C0BF9082C090",
 -9608 => x"C0C0C0BF9082C080",
 -9607 => x"C0C0C0BF9082C0F8",
 -9606 => x"C0C0C0BF9082C082",
 -9605 => x"C0C0C0BF9082C092",
 -9604 => x"C0C0C0BF9082C099",
 -9603 => x"C0C0C0BF9082C0B0",
 -9602 => x"C0C0C0BF9082C0A4",
 -9601 => x"C0C0C0BF9082C0F9",
 -9600 => x"C0C0C0BF9082C0C0",
 -9599 => x"C0C0C0BF90929090",
 -9598 => x"C0C0C0BF90929080",
 -9597 => x"C0C0C0BF909290F8",
 -9596 => x"C0C0C0BF90929082",
 -9595 => x"C0C0C0BF90929092",
 -9594 => x"C0C0C0BF90929099",
 -9593 => x"C0C0C0BF909290B0",
 -9592 => x"C0C0C0BF909290A4",
 -9591 => x"C0C0C0BF909290F9",
 -9590 => x"C0C0C0BF909290C0",
 -9589 => x"C0C0C0BF90928090",
 -9588 => x"C0C0C0BF90928080",
 -9587 => x"C0C0C0BF909280F8",
 -9586 => x"C0C0C0BF90928082",
 -9585 => x"C0C0C0BF90928092",
 -9584 => x"C0C0C0BF90928099",
 -9583 => x"C0C0C0BF909280B0",
 -9582 => x"C0C0C0BF909280A4",
 -9581 => x"C0C0C0BF909280F9",
 -9580 => x"C0C0C0BF909280C0",
 -9579 => x"C0C0C0BF9092F890",
 -9578 => x"C0C0C0BF9092F880",
 -9577 => x"C0C0C0BF9092F8F8",
 -9576 => x"C0C0C0BF9092F882",
 -9575 => x"C0C0C0BF9092F892",
 -9574 => x"C0C0C0BF9092F899",
 -9573 => x"C0C0C0BF9092F8B0",
 -9572 => x"C0C0C0BF9092F8A4",
 -9571 => x"C0C0C0BF9092F8F9",
 -9570 => x"C0C0C0BF9092F8C0",
 -9569 => x"C0C0C0BF90928290",
 -9568 => x"C0C0C0BF90928280",
 -9567 => x"C0C0C0BF909282F8",
 -9566 => x"C0C0C0BF90928282",
 -9565 => x"C0C0C0BF90928292",
 -9564 => x"C0C0C0BF90928299",
 -9563 => x"C0C0C0BF909282B0",
 -9562 => x"C0C0C0BF909282A4",
 -9561 => x"C0C0C0BF909282F9",
 -9560 => x"C0C0C0BF909282C0",
 -9559 => x"C0C0C0BF90929290",
 -9558 => x"C0C0C0BF90929280",
 -9557 => x"C0C0C0BF909292F8",
 -9556 => x"C0C0C0BF90929282",
 -9555 => x"C0C0C0BF90929292",
 -9554 => x"C0C0C0BF90929299",
 -9553 => x"C0C0C0BF909292B0",
 -9552 => x"C0C0C0BF909292A4",
 -9551 => x"C0C0C0BF909292F9",
 -9550 => x"C0C0C0BF909292C0",
 -9549 => x"C0C0C0BF90929990",
 -9548 => x"C0C0C0BF90929980",
 -9547 => x"C0C0C0BF909299F8",
 -9546 => x"C0C0C0BF90929982",
 -9545 => x"C0C0C0BF90929992",
 -9544 => x"C0C0C0BF90929999",
 -9543 => x"C0C0C0BF909299B0",
 -9542 => x"C0C0C0BF909299A4",
 -9541 => x"C0C0C0BF909299F9",
 -9540 => x"C0C0C0BF909299C0",
 -9539 => x"C0C0C0BF9092B090",
 -9538 => x"C0C0C0BF9092B080",
 -9537 => x"C0C0C0BF9092B0F8",
 -9536 => x"C0C0C0BF9092B082",
 -9535 => x"C0C0C0BF9092B092",
 -9534 => x"C0C0C0BF9092B099",
 -9533 => x"C0C0C0BF9092B0B0",
 -9532 => x"C0C0C0BF9092B0A4",
 -9531 => x"C0C0C0BF9092B0F9",
 -9530 => x"C0C0C0BF9092B0C0",
 -9529 => x"C0C0C0BF9092A490",
 -9528 => x"C0C0C0BF9092A480",
 -9527 => x"C0C0C0BF9092A4F8",
 -9526 => x"C0C0C0BF9092A482",
 -9525 => x"C0C0C0BF9092A492",
 -9524 => x"C0C0C0BF9092A499",
 -9523 => x"C0C0C0BF9092A4B0",
 -9522 => x"C0C0C0BF9092A4A4",
 -9521 => x"C0C0C0BF9092A4F9",
 -9520 => x"C0C0C0BF9092A4C0",
 -9519 => x"C0C0C0BF9092F990",
 -9518 => x"C0C0C0BF9092F980",
 -9517 => x"C0C0C0BF9092F9F8",
 -9516 => x"C0C0C0BF9092F982",
 -9515 => x"C0C0C0BF9092F992",
 -9514 => x"C0C0C0BF9092F999",
 -9513 => x"C0C0C0BF9092F9B0",
 -9512 => x"C0C0C0BF9092F9A4",
 -9511 => x"C0C0C0BF9092F9F9",
 -9510 => x"C0C0C0BF9092F9C0",
 -9509 => x"C0C0C0BF9092C090",
 -9508 => x"C0C0C0BF9092C080",
 -9507 => x"C0C0C0BF9092C0F8",
 -9506 => x"C0C0C0BF9092C082",
 -9505 => x"C0C0C0BF9092C092",
 -9504 => x"C0C0C0BF9092C099",
 -9503 => x"C0C0C0BF9092C0B0",
 -9502 => x"C0C0C0BF9092C0A4",
 -9501 => x"C0C0C0BF9092C0F9",
 -9500 => x"C0C0C0BF9092C0C0",
 -9499 => x"C0C0C0BF90999090",
 -9498 => x"C0C0C0BF90999080",
 -9497 => x"C0C0C0BF909990F8",
 -9496 => x"C0C0C0BF90999082",
 -9495 => x"C0C0C0BF90999092",
 -9494 => x"C0C0C0BF90999099",
 -9493 => x"C0C0C0BF909990B0",
 -9492 => x"C0C0C0BF909990A4",
 -9491 => x"C0C0C0BF909990F9",
 -9490 => x"C0C0C0BF909990C0",
 -9489 => x"C0C0C0BF90998090",
 -9488 => x"C0C0C0BF90998080",
 -9487 => x"C0C0C0BF909980F8",
 -9486 => x"C0C0C0BF90998082",
 -9485 => x"C0C0C0BF90998092",
 -9484 => x"C0C0C0BF90998099",
 -9483 => x"C0C0C0BF909980B0",
 -9482 => x"C0C0C0BF909980A4",
 -9481 => x"C0C0C0BF909980F9",
 -9480 => x"C0C0C0BF909980C0",
 -9479 => x"C0C0C0BF9099F890",
 -9478 => x"C0C0C0BF9099F880",
 -9477 => x"C0C0C0BF9099F8F8",
 -9476 => x"C0C0C0BF9099F882",
 -9475 => x"C0C0C0BF9099F892",
 -9474 => x"C0C0C0BF9099F899",
 -9473 => x"C0C0C0BF9099F8B0",
 -9472 => x"C0C0C0BF9099F8A4",
 -9471 => x"C0C0C0BF9099F8F9",
 -9470 => x"C0C0C0BF9099F8C0",
 -9469 => x"C0C0C0BF90998290",
 -9468 => x"C0C0C0BF90998280",
 -9467 => x"C0C0C0BF909982F8",
 -9466 => x"C0C0C0BF90998282",
 -9465 => x"C0C0C0BF90998292",
 -9464 => x"C0C0C0BF90998299",
 -9463 => x"C0C0C0BF909982B0",
 -9462 => x"C0C0C0BF909982A4",
 -9461 => x"C0C0C0BF909982F9",
 -9460 => x"C0C0C0BF909982C0",
 -9459 => x"C0C0C0BF90999290",
 -9458 => x"C0C0C0BF90999280",
 -9457 => x"C0C0C0BF909992F8",
 -9456 => x"C0C0C0BF90999282",
 -9455 => x"C0C0C0BF90999292",
 -9454 => x"C0C0C0BF90999299",
 -9453 => x"C0C0C0BF909992B0",
 -9452 => x"C0C0C0BF909992A4",
 -9451 => x"C0C0C0BF909992F9",
 -9450 => x"C0C0C0BF909992C0",
 -9449 => x"C0C0C0BF90999990",
 -9448 => x"C0C0C0BF90999980",
 -9447 => x"C0C0C0BF909999F8",
 -9446 => x"C0C0C0BF90999982",
 -9445 => x"C0C0C0BF90999992",
 -9444 => x"C0C0C0BF90999999",
 -9443 => x"C0C0C0BF909999B0",
 -9442 => x"C0C0C0BF909999A4",
 -9441 => x"C0C0C0BF909999F9",
 -9440 => x"C0C0C0BF909999C0",
 -9439 => x"C0C0C0BF9099B090",
 -9438 => x"C0C0C0BF9099B080",
 -9437 => x"C0C0C0BF9099B0F8",
 -9436 => x"C0C0C0BF9099B082",
 -9435 => x"C0C0C0BF9099B092",
 -9434 => x"C0C0C0BF9099B099",
 -9433 => x"C0C0C0BF9099B0B0",
 -9432 => x"C0C0C0BF9099B0A4",
 -9431 => x"C0C0C0BF9099B0F9",
 -9430 => x"C0C0C0BF9099B0C0",
 -9429 => x"C0C0C0BF9099A490",
 -9428 => x"C0C0C0BF9099A480",
 -9427 => x"C0C0C0BF9099A4F8",
 -9426 => x"C0C0C0BF9099A482",
 -9425 => x"C0C0C0BF9099A492",
 -9424 => x"C0C0C0BF9099A499",
 -9423 => x"C0C0C0BF9099A4B0",
 -9422 => x"C0C0C0BF9099A4A4",
 -9421 => x"C0C0C0BF9099A4F9",
 -9420 => x"C0C0C0BF9099A4C0",
 -9419 => x"C0C0C0BF9099F990",
 -9418 => x"C0C0C0BF9099F980",
 -9417 => x"C0C0C0BF9099F9F8",
 -9416 => x"C0C0C0BF9099F982",
 -9415 => x"C0C0C0BF9099F992",
 -9414 => x"C0C0C0BF9099F999",
 -9413 => x"C0C0C0BF9099F9B0",
 -9412 => x"C0C0C0BF9099F9A4",
 -9411 => x"C0C0C0BF9099F9F9",
 -9410 => x"C0C0C0BF9099F9C0",
 -9409 => x"C0C0C0BF9099C090",
 -9408 => x"C0C0C0BF9099C080",
 -9407 => x"C0C0C0BF9099C0F8",
 -9406 => x"C0C0C0BF9099C082",
 -9405 => x"C0C0C0BF9099C092",
 -9404 => x"C0C0C0BF9099C099",
 -9403 => x"C0C0C0BF9099C0B0",
 -9402 => x"C0C0C0BF9099C0A4",
 -9401 => x"C0C0C0BF9099C0F9",
 -9400 => x"C0C0C0BF9099C0C0",
 -9399 => x"C0C0C0BF90B09090",
 -9398 => x"C0C0C0BF90B09080",
 -9397 => x"C0C0C0BF90B090F8",
 -9396 => x"C0C0C0BF90B09082",
 -9395 => x"C0C0C0BF90B09092",
 -9394 => x"C0C0C0BF90B09099",
 -9393 => x"C0C0C0BF90B090B0",
 -9392 => x"C0C0C0BF90B090A4",
 -9391 => x"C0C0C0BF90B090F9",
 -9390 => x"C0C0C0BF90B090C0",
 -9389 => x"C0C0C0BF90B08090",
 -9388 => x"C0C0C0BF90B08080",
 -9387 => x"C0C0C0BF90B080F8",
 -9386 => x"C0C0C0BF90B08082",
 -9385 => x"C0C0C0BF90B08092",
 -9384 => x"C0C0C0BF90B08099",
 -9383 => x"C0C0C0BF90B080B0",
 -9382 => x"C0C0C0BF90B080A4",
 -9381 => x"C0C0C0BF90B080F9",
 -9380 => x"C0C0C0BF90B080C0",
 -9379 => x"C0C0C0BF90B0F890",
 -9378 => x"C0C0C0BF90B0F880",
 -9377 => x"C0C0C0BF90B0F8F8",
 -9376 => x"C0C0C0BF90B0F882",
 -9375 => x"C0C0C0BF90B0F892",
 -9374 => x"C0C0C0BF90B0F899",
 -9373 => x"C0C0C0BF90B0F8B0",
 -9372 => x"C0C0C0BF90B0F8A4",
 -9371 => x"C0C0C0BF90B0F8F9",
 -9370 => x"C0C0C0BF90B0F8C0",
 -9369 => x"C0C0C0BF90B08290",
 -9368 => x"C0C0C0BF90B08280",
 -9367 => x"C0C0C0BF90B082F8",
 -9366 => x"C0C0C0BF90B08282",
 -9365 => x"C0C0C0BF90B08292",
 -9364 => x"C0C0C0BF90B08299",
 -9363 => x"C0C0C0BF90B082B0",
 -9362 => x"C0C0C0BF90B082A4",
 -9361 => x"C0C0C0BF90B082F9",
 -9360 => x"C0C0C0BF90B082C0",
 -9359 => x"C0C0C0BF90B09290",
 -9358 => x"C0C0C0BF90B09280",
 -9357 => x"C0C0C0BF90B092F8",
 -9356 => x"C0C0C0BF90B09282",
 -9355 => x"C0C0C0BF90B09292",
 -9354 => x"C0C0C0BF90B09299",
 -9353 => x"C0C0C0BF90B092B0",
 -9352 => x"C0C0C0BF90B092A4",
 -9351 => x"C0C0C0BF90B092F9",
 -9350 => x"C0C0C0BF90B092C0",
 -9349 => x"C0C0C0BF90B09990",
 -9348 => x"C0C0C0BF90B09980",
 -9347 => x"C0C0C0BF90B099F8",
 -9346 => x"C0C0C0BF90B09982",
 -9345 => x"C0C0C0BF90B09992",
 -9344 => x"C0C0C0BF90B09999",
 -9343 => x"C0C0C0BF90B099B0",
 -9342 => x"C0C0C0BF90B099A4",
 -9341 => x"C0C0C0BF90B099F9",
 -9340 => x"C0C0C0BF90B099C0",
 -9339 => x"C0C0C0BF90B0B090",
 -9338 => x"C0C0C0BF90B0B080",
 -9337 => x"C0C0C0BF90B0B0F8",
 -9336 => x"C0C0C0BF90B0B082",
 -9335 => x"C0C0C0BF90B0B092",
 -9334 => x"C0C0C0BF90B0B099",
 -9333 => x"C0C0C0BF90B0B0B0",
 -9332 => x"C0C0C0BF90B0B0A4",
 -9331 => x"C0C0C0BF90B0B0F9",
 -9330 => x"C0C0C0BF90B0B0C0",
 -9329 => x"C0C0C0BF90B0A490",
 -9328 => x"C0C0C0BF90B0A480",
 -9327 => x"C0C0C0BF90B0A4F8",
 -9326 => x"C0C0C0BF90B0A482",
 -9325 => x"C0C0C0BF90B0A492",
 -9324 => x"C0C0C0BF90B0A499",
 -9323 => x"C0C0C0BF90B0A4B0",
 -9322 => x"C0C0C0BF90B0A4A4",
 -9321 => x"C0C0C0BF90B0A4F9",
 -9320 => x"C0C0C0BF90B0A4C0",
 -9319 => x"C0C0C0BF90B0F990",
 -9318 => x"C0C0C0BF90B0F980",
 -9317 => x"C0C0C0BF90B0F9F8",
 -9316 => x"C0C0C0BF90B0F982",
 -9315 => x"C0C0C0BF90B0F992",
 -9314 => x"C0C0C0BF90B0F999",
 -9313 => x"C0C0C0BF90B0F9B0",
 -9312 => x"C0C0C0BF90B0F9A4",
 -9311 => x"C0C0C0BF90B0F9F9",
 -9310 => x"C0C0C0BF90B0F9C0",
 -9309 => x"C0C0C0BF90B0C090",
 -9308 => x"C0C0C0BF90B0C080",
 -9307 => x"C0C0C0BF90B0C0F8",
 -9306 => x"C0C0C0BF90B0C082",
 -9305 => x"C0C0C0BF90B0C092",
 -9304 => x"C0C0C0BF90B0C099",
 -9303 => x"C0C0C0BF90B0C0B0",
 -9302 => x"C0C0C0BF90B0C0A4",
 -9301 => x"C0C0C0BF90B0C0F9",
 -9300 => x"C0C0C0BF90B0C0C0",
 -9299 => x"C0C0C0BF90A49090",
 -9298 => x"C0C0C0BF90A49080",
 -9297 => x"C0C0C0BF90A490F8",
 -9296 => x"C0C0C0BF90A49082",
 -9295 => x"C0C0C0BF90A49092",
 -9294 => x"C0C0C0BF90A49099",
 -9293 => x"C0C0C0BF90A490B0",
 -9292 => x"C0C0C0BF90A490A4",
 -9291 => x"C0C0C0BF90A490F9",
 -9290 => x"C0C0C0BF90A490C0",
 -9289 => x"C0C0C0BF90A48090",
 -9288 => x"C0C0C0BF90A48080",
 -9287 => x"C0C0C0BF90A480F8",
 -9286 => x"C0C0C0BF90A48082",
 -9285 => x"C0C0C0BF90A48092",
 -9284 => x"C0C0C0BF90A48099",
 -9283 => x"C0C0C0BF90A480B0",
 -9282 => x"C0C0C0BF90A480A4",
 -9281 => x"C0C0C0BF90A480F9",
 -9280 => x"C0C0C0BF90A480C0",
 -9279 => x"C0C0C0BF90A4F890",
 -9278 => x"C0C0C0BF90A4F880",
 -9277 => x"C0C0C0BF90A4F8F8",
 -9276 => x"C0C0C0BF90A4F882",
 -9275 => x"C0C0C0BF90A4F892",
 -9274 => x"C0C0C0BF90A4F899",
 -9273 => x"C0C0C0BF90A4F8B0",
 -9272 => x"C0C0C0BF90A4F8A4",
 -9271 => x"C0C0C0BF90A4F8F9",
 -9270 => x"C0C0C0BF90A4F8C0",
 -9269 => x"C0C0C0BF90A48290",
 -9268 => x"C0C0C0BF90A48280",
 -9267 => x"C0C0C0BF90A482F8",
 -9266 => x"C0C0C0BF90A48282",
 -9265 => x"C0C0C0BF90A48292",
 -9264 => x"C0C0C0BF90A48299",
 -9263 => x"C0C0C0BF90A482B0",
 -9262 => x"C0C0C0BF90A482A4",
 -9261 => x"C0C0C0BF90A482F9",
 -9260 => x"C0C0C0BF90A482C0",
 -9259 => x"C0C0C0BF90A49290",
 -9258 => x"C0C0C0BF90A49280",
 -9257 => x"C0C0C0BF90A492F8",
 -9256 => x"C0C0C0BF90A49282",
 -9255 => x"C0C0C0BF90A49292",
 -9254 => x"C0C0C0BF90A49299",
 -9253 => x"C0C0C0BF90A492B0",
 -9252 => x"C0C0C0BF90A492A4",
 -9251 => x"C0C0C0BF90A492F9",
 -9250 => x"C0C0C0BF90A492C0",
 -9249 => x"C0C0C0BF90A49990",
 -9248 => x"C0C0C0BF90A49980",
 -9247 => x"C0C0C0BF90A499F8",
 -9246 => x"C0C0C0BF90A49982",
 -9245 => x"C0C0C0BF90A49992",
 -9244 => x"C0C0C0BF90A49999",
 -9243 => x"C0C0C0BF90A499B0",
 -9242 => x"C0C0C0BF90A499A4",
 -9241 => x"C0C0C0BF90A499F9",
 -9240 => x"C0C0C0BF90A499C0",
 -9239 => x"C0C0C0BF90A4B090",
 -9238 => x"C0C0C0BF90A4B080",
 -9237 => x"C0C0C0BF90A4B0F8",
 -9236 => x"C0C0C0BF90A4B082",
 -9235 => x"C0C0C0BF90A4B092",
 -9234 => x"C0C0C0BF90A4B099",
 -9233 => x"C0C0C0BF90A4B0B0",
 -9232 => x"C0C0C0BF90A4B0A4",
 -9231 => x"C0C0C0BF90A4B0F9",
 -9230 => x"C0C0C0BF90A4B0C0",
 -9229 => x"C0C0C0BF90A4A490",
 -9228 => x"C0C0C0BF90A4A480",
 -9227 => x"C0C0C0BF90A4A4F8",
 -9226 => x"C0C0C0BF90A4A482",
 -9225 => x"C0C0C0BF90A4A492",
 -9224 => x"C0C0C0BF90A4A499",
 -9223 => x"C0C0C0BF90A4A4B0",
 -9222 => x"C0C0C0BF90A4A4A4",
 -9221 => x"C0C0C0BF90A4A4F9",
 -9220 => x"C0C0C0BF90A4A4C0",
 -9219 => x"C0C0C0BF90A4F990",
 -9218 => x"C0C0C0BF90A4F980",
 -9217 => x"C0C0C0BF90A4F9F8",
 -9216 => x"C0C0C0BF90A4F982",
 -9215 => x"C0C0C0BF90A4F992",
 -9214 => x"C0C0C0BF90A4F999",
 -9213 => x"C0C0C0BF90A4F9B0",
 -9212 => x"C0C0C0BF90A4F9A4",
 -9211 => x"C0C0C0BF90A4F9F9",
 -9210 => x"C0C0C0BF90A4F9C0",
 -9209 => x"C0C0C0BF90A4C090",
 -9208 => x"C0C0C0BF90A4C080",
 -9207 => x"C0C0C0BF90A4C0F8",
 -9206 => x"C0C0C0BF90A4C082",
 -9205 => x"C0C0C0BF90A4C092",
 -9204 => x"C0C0C0BF90A4C099",
 -9203 => x"C0C0C0BF90A4C0B0",
 -9202 => x"C0C0C0BF90A4C0A4",
 -9201 => x"C0C0C0BF90A4C0F9",
 -9200 => x"C0C0C0BF90A4C0C0",
 -9199 => x"C0C0C0BF90F99090",
 -9198 => x"C0C0C0BF90F99080",
 -9197 => x"C0C0C0BF90F990F8",
 -9196 => x"C0C0C0BF90F99082",
 -9195 => x"C0C0C0BF90F99092",
 -9194 => x"C0C0C0BF90F99099",
 -9193 => x"C0C0C0BF90F990B0",
 -9192 => x"C0C0C0BF90F990A4",
 -9191 => x"C0C0C0BF90F990F9",
 -9190 => x"C0C0C0BF90F990C0",
 -9189 => x"C0C0C0BF90F98090",
 -9188 => x"C0C0C0BF90F98080",
 -9187 => x"C0C0C0BF90F980F8",
 -9186 => x"C0C0C0BF90F98082",
 -9185 => x"C0C0C0BF90F98092",
 -9184 => x"C0C0C0BF90F98099",
 -9183 => x"C0C0C0BF90F980B0",
 -9182 => x"C0C0C0BF90F980A4",
 -9181 => x"C0C0C0BF90F980F9",
 -9180 => x"C0C0C0BF90F980C0",
 -9179 => x"C0C0C0BF90F9F890",
 -9178 => x"C0C0C0BF90F9F880",
 -9177 => x"C0C0C0BF90F9F8F8",
 -9176 => x"C0C0C0BF90F9F882",
 -9175 => x"C0C0C0BF90F9F892",
 -9174 => x"C0C0C0BF90F9F899",
 -9173 => x"C0C0C0BF90F9F8B0",
 -9172 => x"C0C0C0BF90F9F8A4",
 -9171 => x"C0C0C0BF90F9F8F9",
 -9170 => x"C0C0C0BF90F9F8C0",
 -9169 => x"C0C0C0BF90F98290",
 -9168 => x"C0C0C0BF90F98280",
 -9167 => x"C0C0C0BF90F982F8",
 -9166 => x"C0C0C0BF90F98282",
 -9165 => x"C0C0C0BF90F98292",
 -9164 => x"C0C0C0BF90F98299",
 -9163 => x"C0C0C0BF90F982B0",
 -9162 => x"C0C0C0BF90F982A4",
 -9161 => x"C0C0C0BF90F982F9",
 -9160 => x"C0C0C0BF90F982C0",
 -9159 => x"C0C0C0BF90F99290",
 -9158 => x"C0C0C0BF90F99280",
 -9157 => x"C0C0C0BF90F992F8",
 -9156 => x"C0C0C0BF90F99282",
 -9155 => x"C0C0C0BF90F99292",
 -9154 => x"C0C0C0BF90F99299",
 -9153 => x"C0C0C0BF90F992B0",
 -9152 => x"C0C0C0BF90F992A4",
 -9151 => x"C0C0C0BF90F992F9",
 -9150 => x"C0C0C0BF90F992C0",
 -9149 => x"C0C0C0BF90F99990",
 -9148 => x"C0C0C0BF90F99980",
 -9147 => x"C0C0C0BF90F999F8",
 -9146 => x"C0C0C0BF90F99982",
 -9145 => x"C0C0C0BF90F99992",
 -9144 => x"C0C0C0BF90F99999",
 -9143 => x"C0C0C0BF90F999B0",
 -9142 => x"C0C0C0BF90F999A4",
 -9141 => x"C0C0C0BF90F999F9",
 -9140 => x"C0C0C0BF90F999C0",
 -9139 => x"C0C0C0BF90F9B090",
 -9138 => x"C0C0C0BF90F9B080",
 -9137 => x"C0C0C0BF90F9B0F8",
 -9136 => x"C0C0C0BF90F9B082",
 -9135 => x"C0C0C0BF90F9B092",
 -9134 => x"C0C0C0BF90F9B099",
 -9133 => x"C0C0C0BF90F9B0B0",
 -9132 => x"C0C0C0BF90F9B0A4",
 -9131 => x"C0C0C0BF90F9B0F9",
 -9130 => x"C0C0C0BF90F9B0C0",
 -9129 => x"C0C0C0BF90F9A490",
 -9128 => x"C0C0C0BF90F9A480",
 -9127 => x"C0C0C0BF90F9A4F8",
 -9126 => x"C0C0C0BF90F9A482",
 -9125 => x"C0C0C0BF90F9A492",
 -9124 => x"C0C0C0BF90F9A499",
 -9123 => x"C0C0C0BF90F9A4B0",
 -9122 => x"C0C0C0BF90F9A4A4",
 -9121 => x"C0C0C0BF90F9A4F9",
 -9120 => x"C0C0C0BF90F9A4C0",
 -9119 => x"C0C0C0BF90F9F990",
 -9118 => x"C0C0C0BF90F9F980",
 -9117 => x"C0C0C0BF90F9F9F8",
 -9116 => x"C0C0C0BF90F9F982",
 -9115 => x"C0C0C0BF90F9F992",
 -9114 => x"C0C0C0BF90F9F999",
 -9113 => x"C0C0C0BF90F9F9B0",
 -9112 => x"C0C0C0BF90F9F9A4",
 -9111 => x"C0C0C0BF90F9F9F9",
 -9110 => x"C0C0C0BF90F9F9C0",
 -9109 => x"C0C0C0BF90F9C090",
 -9108 => x"C0C0C0BF90F9C080",
 -9107 => x"C0C0C0BF90F9C0F8",
 -9106 => x"C0C0C0BF90F9C082",
 -9105 => x"C0C0C0BF90F9C092",
 -9104 => x"C0C0C0BF90F9C099",
 -9103 => x"C0C0C0BF90F9C0B0",
 -9102 => x"C0C0C0BF90F9C0A4",
 -9101 => x"C0C0C0BF90F9C0F9",
 -9100 => x"C0C0C0BF90F9C0C0",
 -9099 => x"C0C0C0BF90C09090",
 -9098 => x"C0C0C0BF90C09080",
 -9097 => x"C0C0C0BF90C090F8",
 -9096 => x"C0C0C0BF90C09082",
 -9095 => x"C0C0C0BF90C09092",
 -9094 => x"C0C0C0BF90C09099",
 -9093 => x"C0C0C0BF90C090B0",
 -9092 => x"C0C0C0BF90C090A4",
 -9091 => x"C0C0C0BF90C090F9",
 -9090 => x"C0C0C0BF90C090C0",
 -9089 => x"C0C0C0BF90C08090",
 -9088 => x"C0C0C0BF90C08080",
 -9087 => x"C0C0C0BF90C080F8",
 -9086 => x"C0C0C0BF90C08082",
 -9085 => x"C0C0C0BF90C08092",
 -9084 => x"C0C0C0BF90C08099",
 -9083 => x"C0C0C0BF90C080B0",
 -9082 => x"C0C0C0BF90C080A4",
 -9081 => x"C0C0C0BF90C080F9",
 -9080 => x"C0C0C0BF90C080C0",
 -9079 => x"C0C0C0BF90C0F890",
 -9078 => x"C0C0C0BF90C0F880",
 -9077 => x"C0C0C0BF90C0F8F8",
 -9076 => x"C0C0C0BF90C0F882",
 -9075 => x"C0C0C0BF90C0F892",
 -9074 => x"C0C0C0BF90C0F899",
 -9073 => x"C0C0C0BF90C0F8B0",
 -9072 => x"C0C0C0BF90C0F8A4",
 -9071 => x"C0C0C0BF90C0F8F9",
 -9070 => x"C0C0C0BF90C0F8C0",
 -9069 => x"C0C0C0BF90C08290",
 -9068 => x"C0C0C0BF90C08280",
 -9067 => x"C0C0C0BF90C082F8",
 -9066 => x"C0C0C0BF90C08282",
 -9065 => x"C0C0C0BF90C08292",
 -9064 => x"C0C0C0BF90C08299",
 -9063 => x"C0C0C0BF90C082B0",
 -9062 => x"C0C0C0BF90C082A4",
 -9061 => x"C0C0C0BF90C082F9",
 -9060 => x"C0C0C0BF90C082C0",
 -9059 => x"C0C0C0BF90C09290",
 -9058 => x"C0C0C0BF90C09280",
 -9057 => x"C0C0C0BF90C092F8",
 -9056 => x"C0C0C0BF90C09282",
 -9055 => x"C0C0C0BF90C09292",
 -9054 => x"C0C0C0BF90C09299",
 -9053 => x"C0C0C0BF90C092B0",
 -9052 => x"C0C0C0BF90C092A4",
 -9051 => x"C0C0C0BF90C092F9",
 -9050 => x"C0C0C0BF90C092C0",
 -9049 => x"C0C0C0BF90C09990",
 -9048 => x"C0C0C0BF90C09980",
 -9047 => x"C0C0C0BF90C099F8",
 -9046 => x"C0C0C0BF90C09982",
 -9045 => x"C0C0C0BF90C09992",
 -9044 => x"C0C0C0BF90C09999",
 -9043 => x"C0C0C0BF90C099B0",
 -9042 => x"C0C0C0BF90C099A4",
 -9041 => x"C0C0C0BF90C099F9",
 -9040 => x"C0C0C0BF90C099C0",
 -9039 => x"C0C0C0BF90C0B090",
 -9038 => x"C0C0C0BF90C0B080",
 -9037 => x"C0C0C0BF90C0B0F8",
 -9036 => x"C0C0C0BF90C0B082",
 -9035 => x"C0C0C0BF90C0B092",
 -9034 => x"C0C0C0BF90C0B099",
 -9033 => x"C0C0C0BF90C0B0B0",
 -9032 => x"C0C0C0BF90C0B0A4",
 -9031 => x"C0C0C0BF90C0B0F9",
 -9030 => x"C0C0C0BF90C0B0C0",
 -9029 => x"C0C0C0BF90C0A490",
 -9028 => x"C0C0C0BF90C0A480",
 -9027 => x"C0C0C0BF90C0A4F8",
 -9026 => x"C0C0C0BF90C0A482",
 -9025 => x"C0C0C0BF90C0A492",
 -9024 => x"C0C0C0BF90C0A499",
 -9023 => x"C0C0C0BF90C0A4B0",
 -9022 => x"C0C0C0BF90C0A4A4",
 -9021 => x"C0C0C0BF90C0A4F9",
 -9020 => x"C0C0C0BF90C0A4C0",
 -9019 => x"C0C0C0BF90C0F990",
 -9018 => x"C0C0C0BF90C0F980",
 -9017 => x"C0C0C0BF90C0F9F8",
 -9016 => x"C0C0C0BF90C0F982",
 -9015 => x"C0C0C0BF90C0F992",
 -9014 => x"C0C0C0BF90C0F999",
 -9013 => x"C0C0C0BF90C0F9B0",
 -9012 => x"C0C0C0BF90C0F9A4",
 -9011 => x"C0C0C0BF90C0F9F9",
 -9010 => x"C0C0C0BF90C0F9C0",
 -9009 => x"C0C0C0BF90C0C090",
 -9008 => x"C0C0C0BF90C0C080",
 -9007 => x"C0C0C0BF90C0C0F8",
 -9006 => x"C0C0C0BF90C0C082",
 -9005 => x"C0C0C0BF90C0C092",
 -9004 => x"C0C0C0BF90C0C099",
 -9003 => x"C0C0C0BF90C0C0B0",
 -9002 => x"C0C0C0BF90C0C0A4",
 -9001 => x"C0C0C0BF90C0C0F9",
 -9000 => x"C0C0C0BF90C0C0C0",
 -8999 => x"C0C0C0BF80909090",
 -8998 => x"C0C0C0BF80909080",
 -8997 => x"C0C0C0BF809090F8",
 -8996 => x"C0C0C0BF80909082",
 -8995 => x"C0C0C0BF80909092",
 -8994 => x"C0C0C0BF80909099",
 -8993 => x"C0C0C0BF809090B0",
 -8992 => x"C0C0C0BF809090A4",
 -8991 => x"C0C0C0BF809090F9",
 -8990 => x"C0C0C0BF809090C0",
 -8989 => x"C0C0C0BF80908090",
 -8988 => x"C0C0C0BF80908080",
 -8987 => x"C0C0C0BF809080F8",
 -8986 => x"C0C0C0BF80908082",
 -8985 => x"C0C0C0BF80908092",
 -8984 => x"C0C0C0BF80908099",
 -8983 => x"C0C0C0BF809080B0",
 -8982 => x"C0C0C0BF809080A4",
 -8981 => x"C0C0C0BF809080F9",
 -8980 => x"C0C0C0BF809080C0",
 -8979 => x"C0C0C0BF8090F890",
 -8978 => x"C0C0C0BF8090F880",
 -8977 => x"C0C0C0BF8090F8F8",
 -8976 => x"C0C0C0BF8090F882",
 -8975 => x"C0C0C0BF8090F892",
 -8974 => x"C0C0C0BF8090F899",
 -8973 => x"C0C0C0BF8090F8B0",
 -8972 => x"C0C0C0BF8090F8A4",
 -8971 => x"C0C0C0BF8090F8F9",
 -8970 => x"C0C0C0BF8090F8C0",
 -8969 => x"C0C0C0BF80908290",
 -8968 => x"C0C0C0BF80908280",
 -8967 => x"C0C0C0BF809082F8",
 -8966 => x"C0C0C0BF80908282",
 -8965 => x"C0C0C0BF80908292",
 -8964 => x"C0C0C0BF80908299",
 -8963 => x"C0C0C0BF809082B0",
 -8962 => x"C0C0C0BF809082A4",
 -8961 => x"C0C0C0BF809082F9",
 -8960 => x"C0C0C0BF809082C0",
 -8959 => x"C0C0C0BF80909290",
 -8958 => x"C0C0C0BF80909280",
 -8957 => x"C0C0C0BF809092F8",
 -8956 => x"C0C0C0BF80909282",
 -8955 => x"C0C0C0BF80909292",
 -8954 => x"C0C0C0BF80909299",
 -8953 => x"C0C0C0BF809092B0",
 -8952 => x"C0C0C0BF809092A4",
 -8951 => x"C0C0C0BF809092F9",
 -8950 => x"C0C0C0BF809092C0",
 -8949 => x"C0C0C0BF80909990",
 -8948 => x"C0C0C0BF80909980",
 -8947 => x"C0C0C0BF809099F8",
 -8946 => x"C0C0C0BF80909982",
 -8945 => x"C0C0C0BF80909992",
 -8944 => x"C0C0C0BF80909999",
 -8943 => x"C0C0C0BF809099B0",
 -8942 => x"C0C0C0BF809099A4",
 -8941 => x"C0C0C0BF809099F9",
 -8940 => x"C0C0C0BF809099C0",
 -8939 => x"C0C0C0BF8090B090",
 -8938 => x"C0C0C0BF8090B080",
 -8937 => x"C0C0C0BF8090B0F8",
 -8936 => x"C0C0C0BF8090B082",
 -8935 => x"C0C0C0BF8090B092",
 -8934 => x"C0C0C0BF8090B099",
 -8933 => x"C0C0C0BF8090B0B0",
 -8932 => x"C0C0C0BF8090B0A4",
 -8931 => x"C0C0C0BF8090B0F9",
 -8930 => x"C0C0C0BF8090B0C0",
 -8929 => x"C0C0C0BF8090A490",
 -8928 => x"C0C0C0BF8090A480",
 -8927 => x"C0C0C0BF8090A4F8",
 -8926 => x"C0C0C0BF8090A482",
 -8925 => x"C0C0C0BF8090A492",
 -8924 => x"C0C0C0BF8090A499",
 -8923 => x"C0C0C0BF8090A4B0",
 -8922 => x"C0C0C0BF8090A4A4",
 -8921 => x"C0C0C0BF8090A4F9",
 -8920 => x"C0C0C0BF8090A4C0",
 -8919 => x"C0C0C0BF8090F990",
 -8918 => x"C0C0C0BF8090F980",
 -8917 => x"C0C0C0BF8090F9F8",
 -8916 => x"C0C0C0BF8090F982",
 -8915 => x"C0C0C0BF8090F992",
 -8914 => x"C0C0C0BF8090F999",
 -8913 => x"C0C0C0BF8090F9B0",
 -8912 => x"C0C0C0BF8090F9A4",
 -8911 => x"C0C0C0BF8090F9F9",
 -8910 => x"C0C0C0BF8090F9C0",
 -8909 => x"C0C0C0BF8090C090",
 -8908 => x"C0C0C0BF8090C080",
 -8907 => x"C0C0C0BF8090C0F8",
 -8906 => x"C0C0C0BF8090C082",
 -8905 => x"C0C0C0BF8090C092",
 -8904 => x"C0C0C0BF8090C099",
 -8903 => x"C0C0C0BF8090C0B0",
 -8902 => x"C0C0C0BF8090C0A4",
 -8901 => x"C0C0C0BF8090C0F9",
 -8900 => x"C0C0C0BF8090C0C0",
 -8899 => x"C0C0C0BF80809090",
 -8898 => x"C0C0C0BF80809080",
 -8897 => x"C0C0C0BF808090F8",
 -8896 => x"C0C0C0BF80809082",
 -8895 => x"C0C0C0BF80809092",
 -8894 => x"C0C0C0BF80809099",
 -8893 => x"C0C0C0BF808090B0",
 -8892 => x"C0C0C0BF808090A4",
 -8891 => x"C0C0C0BF808090F9",
 -8890 => x"C0C0C0BF808090C0",
 -8889 => x"C0C0C0BF80808090",
 -8888 => x"C0C0C0BF80808080",
 -8887 => x"C0C0C0BF808080F8",
 -8886 => x"C0C0C0BF80808082",
 -8885 => x"C0C0C0BF80808092",
 -8884 => x"C0C0C0BF80808099",
 -8883 => x"C0C0C0BF808080B0",
 -8882 => x"C0C0C0BF808080A4",
 -8881 => x"C0C0C0BF808080F9",
 -8880 => x"C0C0C0BF808080C0",
 -8879 => x"C0C0C0BF8080F890",
 -8878 => x"C0C0C0BF8080F880",
 -8877 => x"C0C0C0BF8080F8F8",
 -8876 => x"C0C0C0BF8080F882",
 -8875 => x"C0C0C0BF8080F892",
 -8874 => x"C0C0C0BF8080F899",
 -8873 => x"C0C0C0BF8080F8B0",
 -8872 => x"C0C0C0BF8080F8A4",
 -8871 => x"C0C0C0BF8080F8F9",
 -8870 => x"C0C0C0BF8080F8C0",
 -8869 => x"C0C0C0BF80808290",
 -8868 => x"C0C0C0BF80808280",
 -8867 => x"C0C0C0BF808082F8",
 -8866 => x"C0C0C0BF80808282",
 -8865 => x"C0C0C0BF80808292",
 -8864 => x"C0C0C0BF80808299",
 -8863 => x"C0C0C0BF808082B0",
 -8862 => x"C0C0C0BF808082A4",
 -8861 => x"C0C0C0BF808082F9",
 -8860 => x"C0C0C0BF808082C0",
 -8859 => x"C0C0C0BF80809290",
 -8858 => x"C0C0C0BF80809280",
 -8857 => x"C0C0C0BF808092F8",
 -8856 => x"C0C0C0BF80809282",
 -8855 => x"C0C0C0BF80809292",
 -8854 => x"C0C0C0BF80809299",
 -8853 => x"C0C0C0BF808092B0",
 -8852 => x"C0C0C0BF808092A4",
 -8851 => x"C0C0C0BF808092F9",
 -8850 => x"C0C0C0BF808092C0",
 -8849 => x"C0C0C0BF80809990",
 -8848 => x"C0C0C0BF80809980",
 -8847 => x"C0C0C0BF808099F8",
 -8846 => x"C0C0C0BF80809982",
 -8845 => x"C0C0C0BF80809992",
 -8844 => x"C0C0C0BF80809999",
 -8843 => x"C0C0C0BF808099B0",
 -8842 => x"C0C0C0BF808099A4",
 -8841 => x"C0C0C0BF808099F9",
 -8840 => x"C0C0C0BF808099C0",
 -8839 => x"C0C0C0BF8080B090",
 -8838 => x"C0C0C0BF8080B080",
 -8837 => x"C0C0C0BF8080B0F8",
 -8836 => x"C0C0C0BF8080B082",
 -8835 => x"C0C0C0BF8080B092",
 -8834 => x"C0C0C0BF8080B099",
 -8833 => x"C0C0C0BF8080B0B0",
 -8832 => x"C0C0C0BF8080B0A4",
 -8831 => x"C0C0C0BF8080B0F9",
 -8830 => x"C0C0C0BF8080B0C0",
 -8829 => x"C0C0C0BF8080A490",
 -8828 => x"C0C0C0BF8080A480",
 -8827 => x"C0C0C0BF8080A4F8",
 -8826 => x"C0C0C0BF8080A482",
 -8825 => x"C0C0C0BF8080A492",
 -8824 => x"C0C0C0BF8080A499",
 -8823 => x"C0C0C0BF8080A4B0",
 -8822 => x"C0C0C0BF8080A4A4",
 -8821 => x"C0C0C0BF8080A4F9",
 -8820 => x"C0C0C0BF8080A4C0",
 -8819 => x"C0C0C0BF8080F990",
 -8818 => x"C0C0C0BF8080F980",
 -8817 => x"C0C0C0BF8080F9F8",
 -8816 => x"C0C0C0BF8080F982",
 -8815 => x"C0C0C0BF8080F992",
 -8814 => x"C0C0C0BF8080F999",
 -8813 => x"C0C0C0BF8080F9B0",
 -8812 => x"C0C0C0BF8080F9A4",
 -8811 => x"C0C0C0BF8080F9F9",
 -8810 => x"C0C0C0BF8080F9C0",
 -8809 => x"C0C0C0BF8080C090",
 -8808 => x"C0C0C0BF8080C080",
 -8807 => x"C0C0C0BF8080C0F8",
 -8806 => x"C0C0C0BF8080C082",
 -8805 => x"C0C0C0BF8080C092",
 -8804 => x"C0C0C0BF8080C099",
 -8803 => x"C0C0C0BF8080C0B0",
 -8802 => x"C0C0C0BF8080C0A4",
 -8801 => x"C0C0C0BF8080C0F9",
 -8800 => x"C0C0C0BF8080C0C0",
 -8799 => x"C0C0C0BF80F89090",
 -8798 => x"C0C0C0BF80F89080",
 -8797 => x"C0C0C0BF80F890F8",
 -8796 => x"C0C0C0BF80F89082",
 -8795 => x"C0C0C0BF80F89092",
 -8794 => x"C0C0C0BF80F89099",
 -8793 => x"C0C0C0BF80F890B0",
 -8792 => x"C0C0C0BF80F890A4",
 -8791 => x"C0C0C0BF80F890F9",
 -8790 => x"C0C0C0BF80F890C0",
 -8789 => x"C0C0C0BF80F88090",
 -8788 => x"C0C0C0BF80F88080",
 -8787 => x"C0C0C0BF80F880F8",
 -8786 => x"C0C0C0BF80F88082",
 -8785 => x"C0C0C0BF80F88092",
 -8784 => x"C0C0C0BF80F88099",
 -8783 => x"C0C0C0BF80F880B0",
 -8782 => x"C0C0C0BF80F880A4",
 -8781 => x"C0C0C0BF80F880F9",
 -8780 => x"C0C0C0BF80F880C0",
 -8779 => x"C0C0C0BF80F8F890",
 -8778 => x"C0C0C0BF80F8F880",
 -8777 => x"C0C0C0BF80F8F8F8",
 -8776 => x"C0C0C0BF80F8F882",
 -8775 => x"C0C0C0BF80F8F892",
 -8774 => x"C0C0C0BF80F8F899",
 -8773 => x"C0C0C0BF80F8F8B0",
 -8772 => x"C0C0C0BF80F8F8A4",
 -8771 => x"C0C0C0BF80F8F8F9",
 -8770 => x"C0C0C0BF80F8F8C0",
 -8769 => x"C0C0C0BF80F88290",
 -8768 => x"C0C0C0BF80F88280",
 -8767 => x"C0C0C0BF80F882F8",
 -8766 => x"C0C0C0BF80F88282",
 -8765 => x"C0C0C0BF80F88292",
 -8764 => x"C0C0C0BF80F88299",
 -8763 => x"C0C0C0BF80F882B0",
 -8762 => x"C0C0C0BF80F882A4",
 -8761 => x"C0C0C0BF80F882F9",
 -8760 => x"C0C0C0BF80F882C0",
 -8759 => x"C0C0C0BF80F89290",
 -8758 => x"C0C0C0BF80F89280",
 -8757 => x"C0C0C0BF80F892F8",
 -8756 => x"C0C0C0BF80F89282",
 -8755 => x"C0C0C0BF80F89292",
 -8754 => x"C0C0C0BF80F89299",
 -8753 => x"C0C0C0BF80F892B0",
 -8752 => x"C0C0C0BF80F892A4",
 -8751 => x"C0C0C0BF80F892F9",
 -8750 => x"C0C0C0BF80F892C0",
 -8749 => x"C0C0C0BF80F89990",
 -8748 => x"C0C0C0BF80F89980",
 -8747 => x"C0C0C0BF80F899F8",
 -8746 => x"C0C0C0BF80F89982",
 -8745 => x"C0C0C0BF80F89992",
 -8744 => x"C0C0C0BF80F89999",
 -8743 => x"C0C0C0BF80F899B0",
 -8742 => x"C0C0C0BF80F899A4",
 -8741 => x"C0C0C0BF80F899F9",
 -8740 => x"C0C0C0BF80F899C0",
 -8739 => x"C0C0C0BF80F8B090",
 -8738 => x"C0C0C0BF80F8B080",
 -8737 => x"C0C0C0BF80F8B0F8",
 -8736 => x"C0C0C0BF80F8B082",
 -8735 => x"C0C0C0BF80F8B092",
 -8734 => x"C0C0C0BF80F8B099",
 -8733 => x"C0C0C0BF80F8B0B0",
 -8732 => x"C0C0C0BF80F8B0A4",
 -8731 => x"C0C0C0BF80F8B0F9",
 -8730 => x"C0C0C0BF80F8B0C0",
 -8729 => x"C0C0C0BF80F8A490",
 -8728 => x"C0C0C0BF80F8A480",
 -8727 => x"C0C0C0BF80F8A4F8",
 -8726 => x"C0C0C0BF80F8A482",
 -8725 => x"C0C0C0BF80F8A492",
 -8724 => x"C0C0C0BF80F8A499",
 -8723 => x"C0C0C0BF80F8A4B0",
 -8722 => x"C0C0C0BF80F8A4A4",
 -8721 => x"C0C0C0BF80F8A4F9",
 -8720 => x"C0C0C0BF80F8A4C0",
 -8719 => x"C0C0C0BF80F8F990",
 -8718 => x"C0C0C0BF80F8F980",
 -8717 => x"C0C0C0BF80F8F9F8",
 -8716 => x"C0C0C0BF80F8F982",
 -8715 => x"C0C0C0BF80F8F992",
 -8714 => x"C0C0C0BF80F8F999",
 -8713 => x"C0C0C0BF80F8F9B0",
 -8712 => x"C0C0C0BF80F8F9A4",
 -8711 => x"C0C0C0BF80F8F9F9",
 -8710 => x"C0C0C0BF80F8F9C0",
 -8709 => x"C0C0C0BF80F8C090",
 -8708 => x"C0C0C0BF80F8C080",
 -8707 => x"C0C0C0BF80F8C0F8",
 -8706 => x"C0C0C0BF80F8C082",
 -8705 => x"C0C0C0BF80F8C092",
 -8704 => x"C0C0C0BF80F8C099",
 -8703 => x"C0C0C0BF80F8C0B0",
 -8702 => x"C0C0C0BF80F8C0A4",
 -8701 => x"C0C0C0BF80F8C0F9",
 -8700 => x"C0C0C0BF80F8C0C0",
 -8699 => x"C0C0C0BF80829090",
 -8698 => x"C0C0C0BF80829080",
 -8697 => x"C0C0C0BF808290F8",
 -8696 => x"C0C0C0BF80829082",
 -8695 => x"C0C0C0BF80829092",
 -8694 => x"C0C0C0BF80829099",
 -8693 => x"C0C0C0BF808290B0",
 -8692 => x"C0C0C0BF808290A4",
 -8691 => x"C0C0C0BF808290F9",
 -8690 => x"C0C0C0BF808290C0",
 -8689 => x"C0C0C0BF80828090",
 -8688 => x"C0C0C0BF80828080",
 -8687 => x"C0C0C0BF808280F8",
 -8686 => x"C0C0C0BF80828082",
 -8685 => x"C0C0C0BF80828092",
 -8684 => x"C0C0C0BF80828099",
 -8683 => x"C0C0C0BF808280B0",
 -8682 => x"C0C0C0BF808280A4",
 -8681 => x"C0C0C0BF808280F9",
 -8680 => x"C0C0C0BF808280C0",
 -8679 => x"C0C0C0BF8082F890",
 -8678 => x"C0C0C0BF8082F880",
 -8677 => x"C0C0C0BF8082F8F8",
 -8676 => x"C0C0C0BF8082F882",
 -8675 => x"C0C0C0BF8082F892",
 -8674 => x"C0C0C0BF8082F899",
 -8673 => x"C0C0C0BF8082F8B0",
 -8672 => x"C0C0C0BF8082F8A4",
 -8671 => x"C0C0C0BF8082F8F9",
 -8670 => x"C0C0C0BF8082F8C0",
 -8669 => x"C0C0C0BF80828290",
 -8668 => x"C0C0C0BF80828280",
 -8667 => x"C0C0C0BF808282F8",
 -8666 => x"C0C0C0BF80828282",
 -8665 => x"C0C0C0BF80828292",
 -8664 => x"C0C0C0BF80828299",
 -8663 => x"C0C0C0BF808282B0",
 -8662 => x"C0C0C0BF808282A4",
 -8661 => x"C0C0C0BF808282F9",
 -8660 => x"C0C0C0BF808282C0",
 -8659 => x"C0C0C0BF80829290",
 -8658 => x"C0C0C0BF80829280",
 -8657 => x"C0C0C0BF808292F8",
 -8656 => x"C0C0C0BF80829282",
 -8655 => x"C0C0C0BF80829292",
 -8654 => x"C0C0C0BF80829299",
 -8653 => x"C0C0C0BF808292B0",
 -8652 => x"C0C0C0BF808292A4",
 -8651 => x"C0C0C0BF808292F9",
 -8650 => x"C0C0C0BF808292C0",
 -8649 => x"C0C0C0BF80829990",
 -8648 => x"C0C0C0BF80829980",
 -8647 => x"C0C0C0BF808299F8",
 -8646 => x"C0C0C0BF80829982",
 -8645 => x"C0C0C0BF80829992",
 -8644 => x"C0C0C0BF80829999",
 -8643 => x"C0C0C0BF808299B0",
 -8642 => x"C0C0C0BF808299A4",
 -8641 => x"C0C0C0BF808299F9",
 -8640 => x"C0C0C0BF808299C0",
 -8639 => x"C0C0C0BF8082B090",
 -8638 => x"C0C0C0BF8082B080",
 -8637 => x"C0C0C0BF8082B0F8",
 -8636 => x"C0C0C0BF8082B082",
 -8635 => x"C0C0C0BF8082B092",
 -8634 => x"C0C0C0BF8082B099",
 -8633 => x"C0C0C0BF8082B0B0",
 -8632 => x"C0C0C0BF8082B0A4",
 -8631 => x"C0C0C0BF8082B0F9",
 -8630 => x"C0C0C0BF8082B0C0",
 -8629 => x"C0C0C0BF8082A490",
 -8628 => x"C0C0C0BF8082A480",
 -8627 => x"C0C0C0BF8082A4F8",
 -8626 => x"C0C0C0BF8082A482",
 -8625 => x"C0C0C0BF8082A492",
 -8624 => x"C0C0C0BF8082A499",
 -8623 => x"C0C0C0BF8082A4B0",
 -8622 => x"C0C0C0BF8082A4A4",
 -8621 => x"C0C0C0BF8082A4F9",
 -8620 => x"C0C0C0BF8082A4C0",
 -8619 => x"C0C0C0BF8082F990",
 -8618 => x"C0C0C0BF8082F980",
 -8617 => x"C0C0C0BF8082F9F8",
 -8616 => x"C0C0C0BF8082F982",
 -8615 => x"C0C0C0BF8082F992",
 -8614 => x"C0C0C0BF8082F999",
 -8613 => x"C0C0C0BF8082F9B0",
 -8612 => x"C0C0C0BF8082F9A4",
 -8611 => x"C0C0C0BF8082F9F9",
 -8610 => x"C0C0C0BF8082F9C0",
 -8609 => x"C0C0C0BF8082C090",
 -8608 => x"C0C0C0BF8082C080",
 -8607 => x"C0C0C0BF8082C0F8",
 -8606 => x"C0C0C0BF8082C082",
 -8605 => x"C0C0C0BF8082C092",
 -8604 => x"C0C0C0BF8082C099",
 -8603 => x"C0C0C0BF8082C0B0",
 -8602 => x"C0C0C0BF8082C0A4",
 -8601 => x"C0C0C0BF8082C0F9",
 -8600 => x"C0C0C0BF8082C0C0",
 -8599 => x"C0C0C0BF80929090",
 -8598 => x"C0C0C0BF80929080",
 -8597 => x"C0C0C0BF809290F8",
 -8596 => x"C0C0C0BF80929082",
 -8595 => x"C0C0C0BF80929092",
 -8594 => x"C0C0C0BF80929099",
 -8593 => x"C0C0C0BF809290B0",
 -8592 => x"C0C0C0BF809290A4",
 -8591 => x"C0C0C0BF809290F9",
 -8590 => x"C0C0C0BF809290C0",
 -8589 => x"C0C0C0BF80928090",
 -8588 => x"C0C0C0BF80928080",
 -8587 => x"C0C0C0BF809280F8",
 -8586 => x"C0C0C0BF80928082",
 -8585 => x"C0C0C0BF80928092",
 -8584 => x"C0C0C0BF80928099",
 -8583 => x"C0C0C0BF809280B0",
 -8582 => x"C0C0C0BF809280A4",
 -8581 => x"C0C0C0BF809280F9",
 -8580 => x"C0C0C0BF809280C0",
 -8579 => x"C0C0C0BF8092F890",
 -8578 => x"C0C0C0BF8092F880",
 -8577 => x"C0C0C0BF8092F8F8",
 -8576 => x"C0C0C0BF8092F882",
 -8575 => x"C0C0C0BF8092F892",
 -8574 => x"C0C0C0BF8092F899",
 -8573 => x"C0C0C0BF8092F8B0",
 -8572 => x"C0C0C0BF8092F8A4",
 -8571 => x"C0C0C0BF8092F8F9",
 -8570 => x"C0C0C0BF8092F8C0",
 -8569 => x"C0C0C0BF80928290",
 -8568 => x"C0C0C0BF80928280",
 -8567 => x"C0C0C0BF809282F8",
 -8566 => x"C0C0C0BF80928282",
 -8565 => x"C0C0C0BF80928292",
 -8564 => x"C0C0C0BF80928299",
 -8563 => x"C0C0C0BF809282B0",
 -8562 => x"C0C0C0BF809282A4",
 -8561 => x"C0C0C0BF809282F9",
 -8560 => x"C0C0C0BF809282C0",
 -8559 => x"C0C0C0BF80929290",
 -8558 => x"C0C0C0BF80929280",
 -8557 => x"C0C0C0BF809292F8",
 -8556 => x"C0C0C0BF80929282",
 -8555 => x"C0C0C0BF80929292",
 -8554 => x"C0C0C0BF80929299",
 -8553 => x"C0C0C0BF809292B0",
 -8552 => x"C0C0C0BF809292A4",
 -8551 => x"C0C0C0BF809292F9",
 -8550 => x"C0C0C0BF809292C0",
 -8549 => x"C0C0C0BF80929990",
 -8548 => x"C0C0C0BF80929980",
 -8547 => x"C0C0C0BF809299F8",
 -8546 => x"C0C0C0BF80929982",
 -8545 => x"C0C0C0BF80929992",
 -8544 => x"C0C0C0BF80929999",
 -8543 => x"C0C0C0BF809299B0",
 -8542 => x"C0C0C0BF809299A4",
 -8541 => x"C0C0C0BF809299F9",
 -8540 => x"C0C0C0BF809299C0",
 -8539 => x"C0C0C0BF8092B090",
 -8538 => x"C0C0C0BF8092B080",
 -8537 => x"C0C0C0BF8092B0F8",
 -8536 => x"C0C0C0BF8092B082",
 -8535 => x"C0C0C0BF8092B092",
 -8534 => x"C0C0C0BF8092B099",
 -8533 => x"C0C0C0BF8092B0B0",
 -8532 => x"C0C0C0BF8092B0A4",
 -8531 => x"C0C0C0BF8092B0F9",
 -8530 => x"C0C0C0BF8092B0C0",
 -8529 => x"C0C0C0BF8092A490",
 -8528 => x"C0C0C0BF8092A480",
 -8527 => x"C0C0C0BF8092A4F8",
 -8526 => x"C0C0C0BF8092A482",
 -8525 => x"C0C0C0BF8092A492",
 -8524 => x"C0C0C0BF8092A499",
 -8523 => x"C0C0C0BF8092A4B0",
 -8522 => x"C0C0C0BF8092A4A4",
 -8521 => x"C0C0C0BF8092A4F9",
 -8520 => x"C0C0C0BF8092A4C0",
 -8519 => x"C0C0C0BF8092F990",
 -8518 => x"C0C0C0BF8092F980",
 -8517 => x"C0C0C0BF8092F9F8",
 -8516 => x"C0C0C0BF8092F982",
 -8515 => x"C0C0C0BF8092F992",
 -8514 => x"C0C0C0BF8092F999",
 -8513 => x"C0C0C0BF8092F9B0",
 -8512 => x"C0C0C0BF8092F9A4",
 -8511 => x"C0C0C0BF8092F9F9",
 -8510 => x"C0C0C0BF8092F9C0",
 -8509 => x"C0C0C0BF8092C090",
 -8508 => x"C0C0C0BF8092C080",
 -8507 => x"C0C0C0BF8092C0F8",
 -8506 => x"C0C0C0BF8092C082",
 -8505 => x"C0C0C0BF8092C092",
 -8504 => x"C0C0C0BF8092C099",
 -8503 => x"C0C0C0BF8092C0B0",
 -8502 => x"C0C0C0BF8092C0A4",
 -8501 => x"C0C0C0BF8092C0F9",
 -8500 => x"C0C0C0BF8092C0C0",
 -8499 => x"C0C0C0BF80999090",
 -8498 => x"C0C0C0BF80999080",
 -8497 => x"C0C0C0BF809990F8",
 -8496 => x"C0C0C0BF80999082",
 -8495 => x"C0C0C0BF80999092",
 -8494 => x"C0C0C0BF80999099",
 -8493 => x"C0C0C0BF809990B0",
 -8492 => x"C0C0C0BF809990A4",
 -8491 => x"C0C0C0BF809990F9",
 -8490 => x"C0C0C0BF809990C0",
 -8489 => x"C0C0C0BF80998090",
 -8488 => x"C0C0C0BF80998080",
 -8487 => x"C0C0C0BF809980F8",
 -8486 => x"C0C0C0BF80998082",
 -8485 => x"C0C0C0BF80998092",
 -8484 => x"C0C0C0BF80998099",
 -8483 => x"C0C0C0BF809980B0",
 -8482 => x"C0C0C0BF809980A4",
 -8481 => x"C0C0C0BF809980F9",
 -8480 => x"C0C0C0BF809980C0",
 -8479 => x"C0C0C0BF8099F890",
 -8478 => x"C0C0C0BF8099F880",
 -8477 => x"C0C0C0BF8099F8F8",
 -8476 => x"C0C0C0BF8099F882",
 -8475 => x"C0C0C0BF8099F892",
 -8474 => x"C0C0C0BF8099F899",
 -8473 => x"C0C0C0BF8099F8B0",
 -8472 => x"C0C0C0BF8099F8A4",
 -8471 => x"C0C0C0BF8099F8F9",
 -8470 => x"C0C0C0BF8099F8C0",
 -8469 => x"C0C0C0BF80998290",
 -8468 => x"C0C0C0BF80998280",
 -8467 => x"C0C0C0BF809982F8",
 -8466 => x"C0C0C0BF80998282",
 -8465 => x"C0C0C0BF80998292",
 -8464 => x"C0C0C0BF80998299",
 -8463 => x"C0C0C0BF809982B0",
 -8462 => x"C0C0C0BF809982A4",
 -8461 => x"C0C0C0BF809982F9",
 -8460 => x"C0C0C0BF809982C0",
 -8459 => x"C0C0C0BF80999290",
 -8458 => x"C0C0C0BF80999280",
 -8457 => x"C0C0C0BF809992F8",
 -8456 => x"C0C0C0BF80999282",
 -8455 => x"C0C0C0BF80999292",
 -8454 => x"C0C0C0BF80999299",
 -8453 => x"C0C0C0BF809992B0",
 -8452 => x"C0C0C0BF809992A4",
 -8451 => x"C0C0C0BF809992F9",
 -8450 => x"C0C0C0BF809992C0",
 -8449 => x"C0C0C0BF80999990",
 -8448 => x"C0C0C0BF80999980",
 -8447 => x"C0C0C0BF809999F8",
 -8446 => x"C0C0C0BF80999982",
 -8445 => x"C0C0C0BF80999992",
 -8444 => x"C0C0C0BF80999999",
 -8443 => x"C0C0C0BF809999B0",
 -8442 => x"C0C0C0BF809999A4",
 -8441 => x"C0C0C0BF809999F9",
 -8440 => x"C0C0C0BF809999C0",
 -8439 => x"C0C0C0BF8099B090",
 -8438 => x"C0C0C0BF8099B080",
 -8437 => x"C0C0C0BF8099B0F8",
 -8436 => x"C0C0C0BF8099B082",
 -8435 => x"C0C0C0BF8099B092",
 -8434 => x"C0C0C0BF8099B099",
 -8433 => x"C0C0C0BF8099B0B0",
 -8432 => x"C0C0C0BF8099B0A4",
 -8431 => x"C0C0C0BF8099B0F9",
 -8430 => x"C0C0C0BF8099B0C0",
 -8429 => x"C0C0C0BF8099A490",
 -8428 => x"C0C0C0BF8099A480",
 -8427 => x"C0C0C0BF8099A4F8",
 -8426 => x"C0C0C0BF8099A482",
 -8425 => x"C0C0C0BF8099A492",
 -8424 => x"C0C0C0BF8099A499",
 -8423 => x"C0C0C0BF8099A4B0",
 -8422 => x"C0C0C0BF8099A4A4",
 -8421 => x"C0C0C0BF8099A4F9",
 -8420 => x"C0C0C0BF8099A4C0",
 -8419 => x"C0C0C0BF8099F990",
 -8418 => x"C0C0C0BF8099F980",
 -8417 => x"C0C0C0BF8099F9F8",
 -8416 => x"C0C0C0BF8099F982",
 -8415 => x"C0C0C0BF8099F992",
 -8414 => x"C0C0C0BF8099F999",
 -8413 => x"C0C0C0BF8099F9B0",
 -8412 => x"C0C0C0BF8099F9A4",
 -8411 => x"C0C0C0BF8099F9F9",
 -8410 => x"C0C0C0BF8099F9C0",
 -8409 => x"C0C0C0BF8099C090",
 -8408 => x"C0C0C0BF8099C080",
 -8407 => x"C0C0C0BF8099C0F8",
 -8406 => x"C0C0C0BF8099C082",
 -8405 => x"C0C0C0BF8099C092",
 -8404 => x"C0C0C0BF8099C099",
 -8403 => x"C0C0C0BF8099C0B0",
 -8402 => x"C0C0C0BF8099C0A4",
 -8401 => x"C0C0C0BF8099C0F9",
 -8400 => x"C0C0C0BF8099C0C0",
 -8399 => x"C0C0C0BF80B09090",
 -8398 => x"C0C0C0BF80B09080",
 -8397 => x"C0C0C0BF80B090F8",
 -8396 => x"C0C0C0BF80B09082",
 -8395 => x"C0C0C0BF80B09092",
 -8394 => x"C0C0C0BF80B09099",
 -8393 => x"C0C0C0BF80B090B0",
 -8392 => x"C0C0C0BF80B090A4",
 -8391 => x"C0C0C0BF80B090F9",
 -8390 => x"C0C0C0BF80B090C0",
 -8389 => x"C0C0C0BF80B08090",
 -8388 => x"C0C0C0BF80B08080",
 -8387 => x"C0C0C0BF80B080F8",
 -8386 => x"C0C0C0BF80B08082",
 -8385 => x"C0C0C0BF80B08092",
 -8384 => x"C0C0C0BF80B08099",
 -8383 => x"C0C0C0BF80B080B0",
 -8382 => x"C0C0C0BF80B080A4",
 -8381 => x"C0C0C0BF80B080F9",
 -8380 => x"C0C0C0BF80B080C0",
 -8379 => x"C0C0C0BF80B0F890",
 -8378 => x"C0C0C0BF80B0F880",
 -8377 => x"C0C0C0BF80B0F8F8",
 -8376 => x"C0C0C0BF80B0F882",
 -8375 => x"C0C0C0BF80B0F892",
 -8374 => x"C0C0C0BF80B0F899",
 -8373 => x"C0C0C0BF80B0F8B0",
 -8372 => x"C0C0C0BF80B0F8A4",
 -8371 => x"C0C0C0BF80B0F8F9",
 -8370 => x"C0C0C0BF80B0F8C0",
 -8369 => x"C0C0C0BF80B08290",
 -8368 => x"C0C0C0BF80B08280",
 -8367 => x"C0C0C0BF80B082F8",
 -8366 => x"C0C0C0BF80B08282",
 -8365 => x"C0C0C0BF80B08292",
 -8364 => x"C0C0C0BF80B08299",
 -8363 => x"C0C0C0BF80B082B0",
 -8362 => x"C0C0C0BF80B082A4",
 -8361 => x"C0C0C0BF80B082F9",
 -8360 => x"C0C0C0BF80B082C0",
 -8359 => x"C0C0C0BF80B09290",
 -8358 => x"C0C0C0BF80B09280",
 -8357 => x"C0C0C0BF80B092F8",
 -8356 => x"C0C0C0BF80B09282",
 -8355 => x"C0C0C0BF80B09292",
 -8354 => x"C0C0C0BF80B09299",
 -8353 => x"C0C0C0BF80B092B0",
 -8352 => x"C0C0C0BF80B092A4",
 -8351 => x"C0C0C0BF80B092F9",
 -8350 => x"C0C0C0BF80B092C0",
 -8349 => x"C0C0C0BF80B09990",
 -8348 => x"C0C0C0BF80B09980",
 -8347 => x"C0C0C0BF80B099F8",
 -8346 => x"C0C0C0BF80B09982",
 -8345 => x"C0C0C0BF80B09992",
 -8344 => x"C0C0C0BF80B09999",
 -8343 => x"C0C0C0BF80B099B0",
 -8342 => x"C0C0C0BF80B099A4",
 -8341 => x"C0C0C0BF80B099F9",
 -8340 => x"C0C0C0BF80B099C0",
 -8339 => x"C0C0C0BF80B0B090",
 -8338 => x"C0C0C0BF80B0B080",
 -8337 => x"C0C0C0BF80B0B0F8",
 -8336 => x"C0C0C0BF80B0B082",
 -8335 => x"C0C0C0BF80B0B092",
 -8334 => x"C0C0C0BF80B0B099",
 -8333 => x"C0C0C0BF80B0B0B0",
 -8332 => x"C0C0C0BF80B0B0A4",
 -8331 => x"C0C0C0BF80B0B0F9",
 -8330 => x"C0C0C0BF80B0B0C0",
 -8329 => x"C0C0C0BF80B0A490",
 -8328 => x"C0C0C0BF80B0A480",
 -8327 => x"C0C0C0BF80B0A4F8",
 -8326 => x"C0C0C0BF80B0A482",
 -8325 => x"C0C0C0BF80B0A492",
 -8324 => x"C0C0C0BF80B0A499",
 -8323 => x"C0C0C0BF80B0A4B0",
 -8322 => x"C0C0C0BF80B0A4A4",
 -8321 => x"C0C0C0BF80B0A4F9",
 -8320 => x"C0C0C0BF80B0A4C0",
 -8319 => x"C0C0C0BF80B0F990",
 -8318 => x"C0C0C0BF80B0F980",
 -8317 => x"C0C0C0BF80B0F9F8",
 -8316 => x"C0C0C0BF80B0F982",
 -8315 => x"C0C0C0BF80B0F992",
 -8314 => x"C0C0C0BF80B0F999",
 -8313 => x"C0C0C0BF80B0F9B0",
 -8312 => x"C0C0C0BF80B0F9A4",
 -8311 => x"C0C0C0BF80B0F9F9",
 -8310 => x"C0C0C0BF80B0F9C0",
 -8309 => x"C0C0C0BF80B0C090",
 -8308 => x"C0C0C0BF80B0C080",
 -8307 => x"C0C0C0BF80B0C0F8",
 -8306 => x"C0C0C0BF80B0C082",
 -8305 => x"C0C0C0BF80B0C092",
 -8304 => x"C0C0C0BF80B0C099",
 -8303 => x"C0C0C0BF80B0C0B0",
 -8302 => x"C0C0C0BF80B0C0A4",
 -8301 => x"C0C0C0BF80B0C0F9",
 -8300 => x"C0C0C0BF80B0C0C0",
 -8299 => x"C0C0C0BF80A49090",
 -8298 => x"C0C0C0BF80A49080",
 -8297 => x"C0C0C0BF80A490F8",
 -8296 => x"C0C0C0BF80A49082",
 -8295 => x"C0C0C0BF80A49092",
 -8294 => x"C0C0C0BF80A49099",
 -8293 => x"C0C0C0BF80A490B0",
 -8292 => x"C0C0C0BF80A490A4",
 -8291 => x"C0C0C0BF80A490F9",
 -8290 => x"C0C0C0BF80A490C0",
 -8289 => x"C0C0C0BF80A48090",
 -8288 => x"C0C0C0BF80A48080",
 -8287 => x"C0C0C0BF80A480F8",
 -8286 => x"C0C0C0BF80A48082",
 -8285 => x"C0C0C0BF80A48092",
 -8284 => x"C0C0C0BF80A48099",
 -8283 => x"C0C0C0BF80A480B0",
 -8282 => x"C0C0C0BF80A480A4",
 -8281 => x"C0C0C0BF80A480F9",
 -8280 => x"C0C0C0BF80A480C0",
 -8279 => x"C0C0C0BF80A4F890",
 -8278 => x"C0C0C0BF80A4F880",
 -8277 => x"C0C0C0BF80A4F8F8",
 -8276 => x"C0C0C0BF80A4F882",
 -8275 => x"C0C0C0BF80A4F892",
 -8274 => x"C0C0C0BF80A4F899",
 -8273 => x"C0C0C0BF80A4F8B0",
 -8272 => x"C0C0C0BF80A4F8A4",
 -8271 => x"C0C0C0BF80A4F8F9",
 -8270 => x"C0C0C0BF80A4F8C0",
 -8269 => x"C0C0C0BF80A48290",
 -8268 => x"C0C0C0BF80A48280",
 -8267 => x"C0C0C0BF80A482F8",
 -8266 => x"C0C0C0BF80A48282",
 -8265 => x"C0C0C0BF80A48292",
 -8264 => x"C0C0C0BF80A48299",
 -8263 => x"C0C0C0BF80A482B0",
 -8262 => x"C0C0C0BF80A482A4",
 -8261 => x"C0C0C0BF80A482F9",
 -8260 => x"C0C0C0BF80A482C0",
 -8259 => x"C0C0C0BF80A49290",
 -8258 => x"C0C0C0BF80A49280",
 -8257 => x"C0C0C0BF80A492F8",
 -8256 => x"C0C0C0BF80A49282",
 -8255 => x"C0C0C0BF80A49292",
 -8254 => x"C0C0C0BF80A49299",
 -8253 => x"C0C0C0BF80A492B0",
 -8252 => x"C0C0C0BF80A492A4",
 -8251 => x"C0C0C0BF80A492F9",
 -8250 => x"C0C0C0BF80A492C0",
 -8249 => x"C0C0C0BF80A49990",
 -8248 => x"C0C0C0BF80A49980",
 -8247 => x"C0C0C0BF80A499F8",
 -8246 => x"C0C0C0BF80A49982",
 -8245 => x"C0C0C0BF80A49992",
 -8244 => x"C0C0C0BF80A49999",
 -8243 => x"C0C0C0BF80A499B0",
 -8242 => x"C0C0C0BF80A499A4",
 -8241 => x"C0C0C0BF80A499F9",
 -8240 => x"C0C0C0BF80A499C0",
 -8239 => x"C0C0C0BF80A4B090",
 -8238 => x"C0C0C0BF80A4B080",
 -8237 => x"C0C0C0BF80A4B0F8",
 -8236 => x"C0C0C0BF80A4B082",
 -8235 => x"C0C0C0BF80A4B092",
 -8234 => x"C0C0C0BF80A4B099",
 -8233 => x"C0C0C0BF80A4B0B0",
 -8232 => x"C0C0C0BF80A4B0A4",
 -8231 => x"C0C0C0BF80A4B0F9",
 -8230 => x"C0C0C0BF80A4B0C0",
 -8229 => x"C0C0C0BF80A4A490",
 -8228 => x"C0C0C0BF80A4A480",
 -8227 => x"C0C0C0BF80A4A4F8",
 -8226 => x"C0C0C0BF80A4A482",
 -8225 => x"C0C0C0BF80A4A492",
 -8224 => x"C0C0C0BF80A4A499",
 -8223 => x"C0C0C0BF80A4A4B0",
 -8222 => x"C0C0C0BF80A4A4A4",
 -8221 => x"C0C0C0BF80A4A4F9",
 -8220 => x"C0C0C0BF80A4A4C0",
 -8219 => x"C0C0C0BF80A4F990",
 -8218 => x"C0C0C0BF80A4F980",
 -8217 => x"C0C0C0BF80A4F9F8",
 -8216 => x"C0C0C0BF80A4F982",
 -8215 => x"C0C0C0BF80A4F992",
 -8214 => x"C0C0C0BF80A4F999",
 -8213 => x"C0C0C0BF80A4F9B0",
 -8212 => x"C0C0C0BF80A4F9A4",
 -8211 => x"C0C0C0BF80A4F9F9",
 -8210 => x"C0C0C0BF80A4F9C0",
 -8209 => x"C0C0C0BF80A4C090",
 -8208 => x"C0C0C0BF80A4C080",
 -8207 => x"C0C0C0BF80A4C0F8",
 -8206 => x"C0C0C0BF80A4C082",
 -8205 => x"C0C0C0BF80A4C092",
 -8204 => x"C0C0C0BF80A4C099",
 -8203 => x"C0C0C0BF80A4C0B0",
 -8202 => x"C0C0C0BF80A4C0A4",
 -8201 => x"C0C0C0BF80A4C0F9",
 -8200 => x"C0C0C0BF80A4C0C0",
 -8199 => x"C0C0C0BF80F99090",
 -8198 => x"C0C0C0BF80F99080",
 -8197 => x"C0C0C0BF80F990F8",
 -8196 => x"C0C0C0BF80F99082",
 -8195 => x"C0C0C0BF80F99092",
 -8194 => x"C0C0C0BF80F99099",
 -8193 => x"C0C0C0BF80F990B0",
 -8192 => x"C0C0C0BF80F990A4",
 -8191 => x"C0C0C0BF80F990F9",
 -8190 => x"C0C0C0BF80F990C0",
 -8189 => x"C0C0C0BF80F98090",
 -8188 => x"C0C0C0BF80F98080",
 -8187 => x"C0C0C0BF80F980F8",
 -8186 => x"C0C0C0BF80F98082",
 -8185 => x"C0C0C0BF80F98092",
 -8184 => x"C0C0C0BF80F98099",
 -8183 => x"C0C0C0BF80F980B0",
 -8182 => x"C0C0C0BF80F980A4",
 -8181 => x"C0C0C0BF80F980F9",
 -8180 => x"C0C0C0BF80F980C0",
 -8179 => x"C0C0C0BF80F9F890",
 -8178 => x"C0C0C0BF80F9F880",
 -8177 => x"C0C0C0BF80F9F8F8",
 -8176 => x"C0C0C0BF80F9F882",
 -8175 => x"C0C0C0BF80F9F892",
 -8174 => x"C0C0C0BF80F9F899",
 -8173 => x"C0C0C0BF80F9F8B0",
 -8172 => x"C0C0C0BF80F9F8A4",
 -8171 => x"C0C0C0BF80F9F8F9",
 -8170 => x"C0C0C0BF80F9F8C0",
 -8169 => x"C0C0C0BF80F98290",
 -8168 => x"C0C0C0BF80F98280",
 -8167 => x"C0C0C0BF80F982F8",
 -8166 => x"C0C0C0BF80F98282",
 -8165 => x"C0C0C0BF80F98292",
 -8164 => x"C0C0C0BF80F98299",
 -8163 => x"C0C0C0BF80F982B0",
 -8162 => x"C0C0C0BF80F982A4",
 -8161 => x"C0C0C0BF80F982F9",
 -8160 => x"C0C0C0BF80F982C0",
 -8159 => x"C0C0C0BF80F99290",
 -8158 => x"C0C0C0BF80F99280",
 -8157 => x"C0C0C0BF80F992F8",
 -8156 => x"C0C0C0BF80F99282",
 -8155 => x"C0C0C0BF80F99292",
 -8154 => x"C0C0C0BF80F99299",
 -8153 => x"C0C0C0BF80F992B0",
 -8152 => x"C0C0C0BF80F992A4",
 -8151 => x"C0C0C0BF80F992F9",
 -8150 => x"C0C0C0BF80F992C0",
 -8149 => x"C0C0C0BF80F99990",
 -8148 => x"C0C0C0BF80F99980",
 -8147 => x"C0C0C0BF80F999F8",
 -8146 => x"C0C0C0BF80F99982",
 -8145 => x"C0C0C0BF80F99992",
 -8144 => x"C0C0C0BF80F99999",
 -8143 => x"C0C0C0BF80F999B0",
 -8142 => x"C0C0C0BF80F999A4",
 -8141 => x"C0C0C0BF80F999F9",
 -8140 => x"C0C0C0BF80F999C0",
 -8139 => x"C0C0C0BF80F9B090",
 -8138 => x"C0C0C0BF80F9B080",
 -8137 => x"C0C0C0BF80F9B0F8",
 -8136 => x"C0C0C0BF80F9B082",
 -8135 => x"C0C0C0BF80F9B092",
 -8134 => x"C0C0C0BF80F9B099",
 -8133 => x"C0C0C0BF80F9B0B0",
 -8132 => x"C0C0C0BF80F9B0A4",
 -8131 => x"C0C0C0BF80F9B0F9",
 -8130 => x"C0C0C0BF80F9B0C0",
 -8129 => x"C0C0C0BF80F9A490",
 -8128 => x"C0C0C0BF80F9A480",
 -8127 => x"C0C0C0BF80F9A4F8",
 -8126 => x"C0C0C0BF80F9A482",
 -8125 => x"C0C0C0BF80F9A492",
 -8124 => x"C0C0C0BF80F9A499",
 -8123 => x"C0C0C0BF80F9A4B0",
 -8122 => x"C0C0C0BF80F9A4A4",
 -8121 => x"C0C0C0BF80F9A4F9",
 -8120 => x"C0C0C0BF80F9A4C0",
 -8119 => x"C0C0C0BF80F9F990",
 -8118 => x"C0C0C0BF80F9F980",
 -8117 => x"C0C0C0BF80F9F9F8",
 -8116 => x"C0C0C0BF80F9F982",
 -8115 => x"C0C0C0BF80F9F992",
 -8114 => x"C0C0C0BF80F9F999",
 -8113 => x"C0C0C0BF80F9F9B0",
 -8112 => x"C0C0C0BF80F9F9A4",
 -8111 => x"C0C0C0BF80F9F9F9",
 -8110 => x"C0C0C0BF80F9F9C0",
 -8109 => x"C0C0C0BF80F9C090",
 -8108 => x"C0C0C0BF80F9C080",
 -8107 => x"C0C0C0BF80F9C0F8",
 -8106 => x"C0C0C0BF80F9C082",
 -8105 => x"C0C0C0BF80F9C092",
 -8104 => x"C0C0C0BF80F9C099",
 -8103 => x"C0C0C0BF80F9C0B0",
 -8102 => x"C0C0C0BF80F9C0A4",
 -8101 => x"C0C0C0BF80F9C0F9",
 -8100 => x"C0C0C0BF80F9C0C0",
 -8099 => x"C0C0C0BF80C09090",
 -8098 => x"C0C0C0BF80C09080",
 -8097 => x"C0C0C0BF80C090F8",
 -8096 => x"C0C0C0BF80C09082",
 -8095 => x"C0C0C0BF80C09092",
 -8094 => x"C0C0C0BF80C09099",
 -8093 => x"C0C0C0BF80C090B0",
 -8092 => x"C0C0C0BF80C090A4",
 -8091 => x"C0C0C0BF80C090F9",
 -8090 => x"C0C0C0BF80C090C0",
 -8089 => x"C0C0C0BF80C08090",
 -8088 => x"C0C0C0BF80C08080",
 -8087 => x"C0C0C0BF80C080F8",
 -8086 => x"C0C0C0BF80C08082",
 -8085 => x"C0C0C0BF80C08092",
 -8084 => x"C0C0C0BF80C08099",
 -8083 => x"C0C0C0BF80C080B0",
 -8082 => x"C0C0C0BF80C080A4",
 -8081 => x"C0C0C0BF80C080F9",
 -8080 => x"C0C0C0BF80C080C0",
 -8079 => x"C0C0C0BF80C0F890",
 -8078 => x"C0C0C0BF80C0F880",
 -8077 => x"C0C0C0BF80C0F8F8",
 -8076 => x"C0C0C0BF80C0F882",
 -8075 => x"C0C0C0BF80C0F892",
 -8074 => x"C0C0C0BF80C0F899",
 -8073 => x"C0C0C0BF80C0F8B0",
 -8072 => x"C0C0C0BF80C0F8A4",
 -8071 => x"C0C0C0BF80C0F8F9",
 -8070 => x"C0C0C0BF80C0F8C0",
 -8069 => x"C0C0C0BF80C08290",
 -8068 => x"C0C0C0BF80C08280",
 -8067 => x"C0C0C0BF80C082F8",
 -8066 => x"C0C0C0BF80C08282",
 -8065 => x"C0C0C0BF80C08292",
 -8064 => x"C0C0C0BF80C08299",
 -8063 => x"C0C0C0BF80C082B0",
 -8062 => x"C0C0C0BF80C082A4",
 -8061 => x"C0C0C0BF80C082F9",
 -8060 => x"C0C0C0BF80C082C0",
 -8059 => x"C0C0C0BF80C09290",
 -8058 => x"C0C0C0BF80C09280",
 -8057 => x"C0C0C0BF80C092F8",
 -8056 => x"C0C0C0BF80C09282",
 -8055 => x"C0C0C0BF80C09292",
 -8054 => x"C0C0C0BF80C09299",
 -8053 => x"C0C0C0BF80C092B0",
 -8052 => x"C0C0C0BF80C092A4",
 -8051 => x"C0C0C0BF80C092F9",
 -8050 => x"C0C0C0BF80C092C0",
 -8049 => x"C0C0C0BF80C09990",
 -8048 => x"C0C0C0BF80C09980",
 -8047 => x"C0C0C0BF80C099F8",
 -8046 => x"C0C0C0BF80C09982",
 -8045 => x"C0C0C0BF80C09992",
 -8044 => x"C0C0C0BF80C09999",
 -8043 => x"C0C0C0BF80C099B0",
 -8042 => x"C0C0C0BF80C099A4",
 -8041 => x"C0C0C0BF80C099F9",
 -8040 => x"C0C0C0BF80C099C0",
 -8039 => x"C0C0C0BF80C0B090",
 -8038 => x"C0C0C0BF80C0B080",
 -8037 => x"C0C0C0BF80C0B0F8",
 -8036 => x"C0C0C0BF80C0B082",
 -8035 => x"C0C0C0BF80C0B092",
 -8034 => x"C0C0C0BF80C0B099",
 -8033 => x"C0C0C0BF80C0B0B0",
 -8032 => x"C0C0C0BF80C0B0A4",
 -8031 => x"C0C0C0BF80C0B0F9",
 -8030 => x"C0C0C0BF80C0B0C0",
 -8029 => x"C0C0C0BF80C0A490",
 -8028 => x"C0C0C0BF80C0A480",
 -8027 => x"C0C0C0BF80C0A4F8",
 -8026 => x"C0C0C0BF80C0A482",
 -8025 => x"C0C0C0BF80C0A492",
 -8024 => x"C0C0C0BF80C0A499",
 -8023 => x"C0C0C0BF80C0A4B0",
 -8022 => x"C0C0C0BF80C0A4A4",
 -8021 => x"C0C0C0BF80C0A4F9",
 -8020 => x"C0C0C0BF80C0A4C0",
 -8019 => x"C0C0C0BF80C0F990",
 -8018 => x"C0C0C0BF80C0F980",
 -8017 => x"C0C0C0BF80C0F9F8",
 -8016 => x"C0C0C0BF80C0F982",
 -8015 => x"C0C0C0BF80C0F992",
 -8014 => x"C0C0C0BF80C0F999",
 -8013 => x"C0C0C0BF80C0F9B0",
 -8012 => x"C0C0C0BF80C0F9A4",
 -8011 => x"C0C0C0BF80C0F9F9",
 -8010 => x"C0C0C0BF80C0F9C0",
 -8009 => x"C0C0C0BF80C0C090",
 -8008 => x"C0C0C0BF80C0C080",
 -8007 => x"C0C0C0BF80C0C0F8",
 -8006 => x"C0C0C0BF80C0C082",
 -8005 => x"C0C0C0BF80C0C092",
 -8004 => x"C0C0C0BF80C0C099",
 -8003 => x"C0C0C0BF80C0C0B0",
 -8002 => x"C0C0C0BF80C0C0A4",
 -8001 => x"C0C0C0BF80C0C0F9",
 -8000 => x"C0C0C0BF80C0C0C0",
 -7999 => x"C0C0C0BFF8909090",
 -7998 => x"C0C0C0BFF8909080",
 -7997 => x"C0C0C0BFF89090F8",
 -7996 => x"C0C0C0BFF8909082",
 -7995 => x"C0C0C0BFF8909092",
 -7994 => x"C0C0C0BFF8909099",
 -7993 => x"C0C0C0BFF89090B0",
 -7992 => x"C0C0C0BFF89090A4",
 -7991 => x"C0C0C0BFF89090F9",
 -7990 => x"C0C0C0BFF89090C0",
 -7989 => x"C0C0C0BFF8908090",
 -7988 => x"C0C0C0BFF8908080",
 -7987 => x"C0C0C0BFF89080F8",
 -7986 => x"C0C0C0BFF8908082",
 -7985 => x"C0C0C0BFF8908092",
 -7984 => x"C0C0C0BFF8908099",
 -7983 => x"C0C0C0BFF89080B0",
 -7982 => x"C0C0C0BFF89080A4",
 -7981 => x"C0C0C0BFF89080F9",
 -7980 => x"C0C0C0BFF89080C0",
 -7979 => x"C0C0C0BFF890F890",
 -7978 => x"C0C0C0BFF890F880",
 -7977 => x"C0C0C0BFF890F8F8",
 -7976 => x"C0C0C0BFF890F882",
 -7975 => x"C0C0C0BFF890F892",
 -7974 => x"C0C0C0BFF890F899",
 -7973 => x"C0C0C0BFF890F8B0",
 -7972 => x"C0C0C0BFF890F8A4",
 -7971 => x"C0C0C0BFF890F8F9",
 -7970 => x"C0C0C0BFF890F8C0",
 -7969 => x"C0C0C0BFF8908290",
 -7968 => x"C0C0C0BFF8908280",
 -7967 => x"C0C0C0BFF89082F8",
 -7966 => x"C0C0C0BFF8908282",
 -7965 => x"C0C0C0BFF8908292",
 -7964 => x"C0C0C0BFF8908299",
 -7963 => x"C0C0C0BFF89082B0",
 -7962 => x"C0C0C0BFF89082A4",
 -7961 => x"C0C0C0BFF89082F9",
 -7960 => x"C0C0C0BFF89082C0",
 -7959 => x"C0C0C0BFF8909290",
 -7958 => x"C0C0C0BFF8909280",
 -7957 => x"C0C0C0BFF89092F8",
 -7956 => x"C0C0C0BFF8909282",
 -7955 => x"C0C0C0BFF8909292",
 -7954 => x"C0C0C0BFF8909299",
 -7953 => x"C0C0C0BFF89092B0",
 -7952 => x"C0C0C0BFF89092A4",
 -7951 => x"C0C0C0BFF89092F9",
 -7950 => x"C0C0C0BFF89092C0",
 -7949 => x"C0C0C0BFF8909990",
 -7948 => x"C0C0C0BFF8909980",
 -7947 => x"C0C0C0BFF89099F8",
 -7946 => x"C0C0C0BFF8909982",
 -7945 => x"C0C0C0BFF8909992",
 -7944 => x"C0C0C0BFF8909999",
 -7943 => x"C0C0C0BFF89099B0",
 -7942 => x"C0C0C0BFF89099A4",
 -7941 => x"C0C0C0BFF89099F9",
 -7940 => x"C0C0C0BFF89099C0",
 -7939 => x"C0C0C0BFF890B090",
 -7938 => x"C0C0C0BFF890B080",
 -7937 => x"C0C0C0BFF890B0F8",
 -7936 => x"C0C0C0BFF890B082",
 -7935 => x"C0C0C0BFF890B092",
 -7934 => x"C0C0C0BFF890B099",
 -7933 => x"C0C0C0BFF890B0B0",
 -7932 => x"C0C0C0BFF890B0A4",
 -7931 => x"C0C0C0BFF890B0F9",
 -7930 => x"C0C0C0BFF890B0C0",
 -7929 => x"C0C0C0BFF890A490",
 -7928 => x"C0C0C0BFF890A480",
 -7927 => x"C0C0C0BFF890A4F8",
 -7926 => x"C0C0C0BFF890A482",
 -7925 => x"C0C0C0BFF890A492",
 -7924 => x"C0C0C0BFF890A499",
 -7923 => x"C0C0C0BFF890A4B0",
 -7922 => x"C0C0C0BFF890A4A4",
 -7921 => x"C0C0C0BFF890A4F9",
 -7920 => x"C0C0C0BFF890A4C0",
 -7919 => x"C0C0C0BFF890F990",
 -7918 => x"C0C0C0BFF890F980",
 -7917 => x"C0C0C0BFF890F9F8",
 -7916 => x"C0C0C0BFF890F982",
 -7915 => x"C0C0C0BFF890F992",
 -7914 => x"C0C0C0BFF890F999",
 -7913 => x"C0C0C0BFF890F9B0",
 -7912 => x"C0C0C0BFF890F9A4",
 -7911 => x"C0C0C0BFF890F9F9",
 -7910 => x"C0C0C0BFF890F9C0",
 -7909 => x"C0C0C0BFF890C090",
 -7908 => x"C0C0C0BFF890C080",
 -7907 => x"C0C0C0BFF890C0F8",
 -7906 => x"C0C0C0BFF890C082",
 -7905 => x"C0C0C0BFF890C092",
 -7904 => x"C0C0C0BFF890C099",
 -7903 => x"C0C0C0BFF890C0B0",
 -7902 => x"C0C0C0BFF890C0A4",
 -7901 => x"C0C0C0BFF890C0F9",
 -7900 => x"C0C0C0BFF890C0C0",
 -7899 => x"C0C0C0BFF8809090",
 -7898 => x"C0C0C0BFF8809080",
 -7897 => x"C0C0C0BFF88090F8",
 -7896 => x"C0C0C0BFF8809082",
 -7895 => x"C0C0C0BFF8809092",
 -7894 => x"C0C0C0BFF8809099",
 -7893 => x"C0C0C0BFF88090B0",
 -7892 => x"C0C0C0BFF88090A4",
 -7891 => x"C0C0C0BFF88090F9",
 -7890 => x"C0C0C0BFF88090C0",
 -7889 => x"C0C0C0BFF8808090",
 -7888 => x"C0C0C0BFF8808080",
 -7887 => x"C0C0C0BFF88080F8",
 -7886 => x"C0C0C0BFF8808082",
 -7885 => x"C0C0C0BFF8808092",
 -7884 => x"C0C0C0BFF8808099",
 -7883 => x"C0C0C0BFF88080B0",
 -7882 => x"C0C0C0BFF88080A4",
 -7881 => x"C0C0C0BFF88080F9",
 -7880 => x"C0C0C0BFF88080C0",
 -7879 => x"C0C0C0BFF880F890",
 -7878 => x"C0C0C0BFF880F880",
 -7877 => x"C0C0C0BFF880F8F8",
 -7876 => x"C0C0C0BFF880F882",
 -7875 => x"C0C0C0BFF880F892",
 -7874 => x"C0C0C0BFF880F899",
 -7873 => x"C0C0C0BFF880F8B0",
 -7872 => x"C0C0C0BFF880F8A4",
 -7871 => x"C0C0C0BFF880F8F9",
 -7870 => x"C0C0C0BFF880F8C0",
 -7869 => x"C0C0C0BFF8808290",
 -7868 => x"C0C0C0BFF8808280",
 -7867 => x"C0C0C0BFF88082F8",
 -7866 => x"C0C0C0BFF8808282",
 -7865 => x"C0C0C0BFF8808292",
 -7864 => x"C0C0C0BFF8808299",
 -7863 => x"C0C0C0BFF88082B0",
 -7862 => x"C0C0C0BFF88082A4",
 -7861 => x"C0C0C0BFF88082F9",
 -7860 => x"C0C0C0BFF88082C0",
 -7859 => x"C0C0C0BFF8809290",
 -7858 => x"C0C0C0BFF8809280",
 -7857 => x"C0C0C0BFF88092F8",
 -7856 => x"C0C0C0BFF8809282",
 -7855 => x"C0C0C0BFF8809292",
 -7854 => x"C0C0C0BFF8809299",
 -7853 => x"C0C0C0BFF88092B0",
 -7852 => x"C0C0C0BFF88092A4",
 -7851 => x"C0C0C0BFF88092F9",
 -7850 => x"C0C0C0BFF88092C0",
 -7849 => x"C0C0C0BFF8809990",
 -7848 => x"C0C0C0BFF8809980",
 -7847 => x"C0C0C0BFF88099F8",
 -7846 => x"C0C0C0BFF8809982",
 -7845 => x"C0C0C0BFF8809992",
 -7844 => x"C0C0C0BFF8809999",
 -7843 => x"C0C0C0BFF88099B0",
 -7842 => x"C0C0C0BFF88099A4",
 -7841 => x"C0C0C0BFF88099F9",
 -7840 => x"C0C0C0BFF88099C0",
 -7839 => x"C0C0C0BFF880B090",
 -7838 => x"C0C0C0BFF880B080",
 -7837 => x"C0C0C0BFF880B0F8",
 -7836 => x"C0C0C0BFF880B082",
 -7835 => x"C0C0C0BFF880B092",
 -7834 => x"C0C0C0BFF880B099",
 -7833 => x"C0C0C0BFF880B0B0",
 -7832 => x"C0C0C0BFF880B0A4",
 -7831 => x"C0C0C0BFF880B0F9",
 -7830 => x"C0C0C0BFF880B0C0",
 -7829 => x"C0C0C0BFF880A490",
 -7828 => x"C0C0C0BFF880A480",
 -7827 => x"C0C0C0BFF880A4F8",
 -7826 => x"C0C0C0BFF880A482",
 -7825 => x"C0C0C0BFF880A492",
 -7824 => x"C0C0C0BFF880A499",
 -7823 => x"C0C0C0BFF880A4B0",
 -7822 => x"C0C0C0BFF880A4A4",
 -7821 => x"C0C0C0BFF880A4F9",
 -7820 => x"C0C0C0BFF880A4C0",
 -7819 => x"C0C0C0BFF880F990",
 -7818 => x"C0C0C0BFF880F980",
 -7817 => x"C0C0C0BFF880F9F8",
 -7816 => x"C0C0C0BFF880F982",
 -7815 => x"C0C0C0BFF880F992",
 -7814 => x"C0C0C0BFF880F999",
 -7813 => x"C0C0C0BFF880F9B0",
 -7812 => x"C0C0C0BFF880F9A4",
 -7811 => x"C0C0C0BFF880F9F9",
 -7810 => x"C0C0C0BFF880F9C0",
 -7809 => x"C0C0C0BFF880C090",
 -7808 => x"C0C0C0BFF880C080",
 -7807 => x"C0C0C0BFF880C0F8",
 -7806 => x"C0C0C0BFF880C082",
 -7805 => x"C0C0C0BFF880C092",
 -7804 => x"C0C0C0BFF880C099",
 -7803 => x"C0C0C0BFF880C0B0",
 -7802 => x"C0C0C0BFF880C0A4",
 -7801 => x"C0C0C0BFF880C0F9",
 -7800 => x"C0C0C0BFF880C0C0",
 -7799 => x"C0C0C0BFF8F89090",
 -7798 => x"C0C0C0BFF8F89080",
 -7797 => x"C0C0C0BFF8F890F8",
 -7796 => x"C0C0C0BFF8F89082",
 -7795 => x"C0C0C0BFF8F89092",
 -7794 => x"C0C0C0BFF8F89099",
 -7793 => x"C0C0C0BFF8F890B0",
 -7792 => x"C0C0C0BFF8F890A4",
 -7791 => x"C0C0C0BFF8F890F9",
 -7790 => x"C0C0C0BFF8F890C0",
 -7789 => x"C0C0C0BFF8F88090",
 -7788 => x"C0C0C0BFF8F88080",
 -7787 => x"C0C0C0BFF8F880F8",
 -7786 => x"C0C0C0BFF8F88082",
 -7785 => x"C0C0C0BFF8F88092",
 -7784 => x"C0C0C0BFF8F88099",
 -7783 => x"C0C0C0BFF8F880B0",
 -7782 => x"C0C0C0BFF8F880A4",
 -7781 => x"C0C0C0BFF8F880F9",
 -7780 => x"C0C0C0BFF8F880C0",
 -7779 => x"C0C0C0BFF8F8F890",
 -7778 => x"C0C0C0BFF8F8F880",
 -7777 => x"C0C0C0BFF8F8F8F8",
 -7776 => x"C0C0C0BFF8F8F882",
 -7775 => x"C0C0C0BFF8F8F892",
 -7774 => x"C0C0C0BFF8F8F899",
 -7773 => x"C0C0C0BFF8F8F8B0",
 -7772 => x"C0C0C0BFF8F8F8A4",
 -7771 => x"C0C0C0BFF8F8F8F9",
 -7770 => x"C0C0C0BFF8F8F8C0",
 -7769 => x"C0C0C0BFF8F88290",
 -7768 => x"C0C0C0BFF8F88280",
 -7767 => x"C0C0C0BFF8F882F8",
 -7766 => x"C0C0C0BFF8F88282",
 -7765 => x"C0C0C0BFF8F88292",
 -7764 => x"C0C0C0BFF8F88299",
 -7763 => x"C0C0C0BFF8F882B0",
 -7762 => x"C0C0C0BFF8F882A4",
 -7761 => x"C0C0C0BFF8F882F9",
 -7760 => x"C0C0C0BFF8F882C0",
 -7759 => x"C0C0C0BFF8F89290",
 -7758 => x"C0C0C0BFF8F89280",
 -7757 => x"C0C0C0BFF8F892F8",
 -7756 => x"C0C0C0BFF8F89282",
 -7755 => x"C0C0C0BFF8F89292",
 -7754 => x"C0C0C0BFF8F89299",
 -7753 => x"C0C0C0BFF8F892B0",
 -7752 => x"C0C0C0BFF8F892A4",
 -7751 => x"C0C0C0BFF8F892F9",
 -7750 => x"C0C0C0BFF8F892C0",
 -7749 => x"C0C0C0BFF8F89990",
 -7748 => x"C0C0C0BFF8F89980",
 -7747 => x"C0C0C0BFF8F899F8",
 -7746 => x"C0C0C0BFF8F89982",
 -7745 => x"C0C0C0BFF8F89992",
 -7744 => x"C0C0C0BFF8F89999",
 -7743 => x"C0C0C0BFF8F899B0",
 -7742 => x"C0C0C0BFF8F899A4",
 -7741 => x"C0C0C0BFF8F899F9",
 -7740 => x"C0C0C0BFF8F899C0",
 -7739 => x"C0C0C0BFF8F8B090",
 -7738 => x"C0C0C0BFF8F8B080",
 -7737 => x"C0C0C0BFF8F8B0F8",
 -7736 => x"C0C0C0BFF8F8B082",
 -7735 => x"C0C0C0BFF8F8B092",
 -7734 => x"C0C0C0BFF8F8B099",
 -7733 => x"C0C0C0BFF8F8B0B0",
 -7732 => x"C0C0C0BFF8F8B0A4",
 -7731 => x"C0C0C0BFF8F8B0F9",
 -7730 => x"C0C0C0BFF8F8B0C0",
 -7729 => x"C0C0C0BFF8F8A490",
 -7728 => x"C0C0C0BFF8F8A480",
 -7727 => x"C0C0C0BFF8F8A4F8",
 -7726 => x"C0C0C0BFF8F8A482",
 -7725 => x"C0C0C0BFF8F8A492",
 -7724 => x"C0C0C0BFF8F8A499",
 -7723 => x"C0C0C0BFF8F8A4B0",
 -7722 => x"C0C0C0BFF8F8A4A4",
 -7721 => x"C0C0C0BFF8F8A4F9",
 -7720 => x"C0C0C0BFF8F8A4C0",
 -7719 => x"C0C0C0BFF8F8F990",
 -7718 => x"C0C0C0BFF8F8F980",
 -7717 => x"C0C0C0BFF8F8F9F8",
 -7716 => x"C0C0C0BFF8F8F982",
 -7715 => x"C0C0C0BFF8F8F992",
 -7714 => x"C0C0C0BFF8F8F999",
 -7713 => x"C0C0C0BFF8F8F9B0",
 -7712 => x"C0C0C0BFF8F8F9A4",
 -7711 => x"C0C0C0BFF8F8F9F9",
 -7710 => x"C0C0C0BFF8F8F9C0",
 -7709 => x"C0C0C0BFF8F8C090",
 -7708 => x"C0C0C0BFF8F8C080",
 -7707 => x"C0C0C0BFF8F8C0F8",
 -7706 => x"C0C0C0BFF8F8C082",
 -7705 => x"C0C0C0BFF8F8C092",
 -7704 => x"C0C0C0BFF8F8C099",
 -7703 => x"C0C0C0BFF8F8C0B0",
 -7702 => x"C0C0C0BFF8F8C0A4",
 -7701 => x"C0C0C0BFF8F8C0F9",
 -7700 => x"C0C0C0BFF8F8C0C0",
 -7699 => x"C0C0C0BFF8829090",
 -7698 => x"C0C0C0BFF8829080",
 -7697 => x"C0C0C0BFF88290F8",
 -7696 => x"C0C0C0BFF8829082",
 -7695 => x"C0C0C0BFF8829092",
 -7694 => x"C0C0C0BFF8829099",
 -7693 => x"C0C0C0BFF88290B0",
 -7692 => x"C0C0C0BFF88290A4",
 -7691 => x"C0C0C0BFF88290F9",
 -7690 => x"C0C0C0BFF88290C0",
 -7689 => x"C0C0C0BFF8828090",
 -7688 => x"C0C0C0BFF8828080",
 -7687 => x"C0C0C0BFF88280F8",
 -7686 => x"C0C0C0BFF8828082",
 -7685 => x"C0C0C0BFF8828092",
 -7684 => x"C0C0C0BFF8828099",
 -7683 => x"C0C0C0BFF88280B0",
 -7682 => x"C0C0C0BFF88280A4",
 -7681 => x"C0C0C0BFF88280F9",
 -7680 => x"C0C0C0BFF88280C0",
 -7679 => x"C0C0C0BFF882F890",
 -7678 => x"C0C0C0BFF882F880",
 -7677 => x"C0C0C0BFF882F8F8",
 -7676 => x"C0C0C0BFF882F882",
 -7675 => x"C0C0C0BFF882F892",
 -7674 => x"C0C0C0BFF882F899",
 -7673 => x"C0C0C0BFF882F8B0",
 -7672 => x"C0C0C0BFF882F8A4",
 -7671 => x"C0C0C0BFF882F8F9",
 -7670 => x"C0C0C0BFF882F8C0",
 -7669 => x"C0C0C0BFF8828290",
 -7668 => x"C0C0C0BFF8828280",
 -7667 => x"C0C0C0BFF88282F8",
 -7666 => x"C0C0C0BFF8828282",
 -7665 => x"C0C0C0BFF8828292",
 -7664 => x"C0C0C0BFF8828299",
 -7663 => x"C0C0C0BFF88282B0",
 -7662 => x"C0C0C0BFF88282A4",
 -7661 => x"C0C0C0BFF88282F9",
 -7660 => x"C0C0C0BFF88282C0",
 -7659 => x"C0C0C0BFF8829290",
 -7658 => x"C0C0C0BFF8829280",
 -7657 => x"C0C0C0BFF88292F8",
 -7656 => x"C0C0C0BFF8829282",
 -7655 => x"C0C0C0BFF8829292",
 -7654 => x"C0C0C0BFF8829299",
 -7653 => x"C0C0C0BFF88292B0",
 -7652 => x"C0C0C0BFF88292A4",
 -7651 => x"C0C0C0BFF88292F9",
 -7650 => x"C0C0C0BFF88292C0",
 -7649 => x"C0C0C0BFF8829990",
 -7648 => x"C0C0C0BFF8829980",
 -7647 => x"C0C0C0BFF88299F8",
 -7646 => x"C0C0C0BFF8829982",
 -7645 => x"C0C0C0BFF8829992",
 -7644 => x"C0C0C0BFF8829999",
 -7643 => x"C0C0C0BFF88299B0",
 -7642 => x"C0C0C0BFF88299A4",
 -7641 => x"C0C0C0BFF88299F9",
 -7640 => x"C0C0C0BFF88299C0",
 -7639 => x"C0C0C0BFF882B090",
 -7638 => x"C0C0C0BFF882B080",
 -7637 => x"C0C0C0BFF882B0F8",
 -7636 => x"C0C0C0BFF882B082",
 -7635 => x"C0C0C0BFF882B092",
 -7634 => x"C0C0C0BFF882B099",
 -7633 => x"C0C0C0BFF882B0B0",
 -7632 => x"C0C0C0BFF882B0A4",
 -7631 => x"C0C0C0BFF882B0F9",
 -7630 => x"C0C0C0BFF882B0C0",
 -7629 => x"C0C0C0BFF882A490",
 -7628 => x"C0C0C0BFF882A480",
 -7627 => x"C0C0C0BFF882A4F8",
 -7626 => x"C0C0C0BFF882A482",
 -7625 => x"C0C0C0BFF882A492",
 -7624 => x"C0C0C0BFF882A499",
 -7623 => x"C0C0C0BFF882A4B0",
 -7622 => x"C0C0C0BFF882A4A4",
 -7621 => x"C0C0C0BFF882A4F9",
 -7620 => x"C0C0C0BFF882A4C0",
 -7619 => x"C0C0C0BFF882F990",
 -7618 => x"C0C0C0BFF882F980",
 -7617 => x"C0C0C0BFF882F9F8",
 -7616 => x"C0C0C0BFF882F982",
 -7615 => x"C0C0C0BFF882F992",
 -7614 => x"C0C0C0BFF882F999",
 -7613 => x"C0C0C0BFF882F9B0",
 -7612 => x"C0C0C0BFF882F9A4",
 -7611 => x"C0C0C0BFF882F9F9",
 -7610 => x"C0C0C0BFF882F9C0",
 -7609 => x"C0C0C0BFF882C090",
 -7608 => x"C0C0C0BFF882C080",
 -7607 => x"C0C0C0BFF882C0F8",
 -7606 => x"C0C0C0BFF882C082",
 -7605 => x"C0C0C0BFF882C092",
 -7604 => x"C0C0C0BFF882C099",
 -7603 => x"C0C0C0BFF882C0B0",
 -7602 => x"C0C0C0BFF882C0A4",
 -7601 => x"C0C0C0BFF882C0F9",
 -7600 => x"C0C0C0BFF882C0C0",
 -7599 => x"C0C0C0BFF8929090",
 -7598 => x"C0C0C0BFF8929080",
 -7597 => x"C0C0C0BFF89290F8",
 -7596 => x"C0C0C0BFF8929082",
 -7595 => x"C0C0C0BFF8929092",
 -7594 => x"C0C0C0BFF8929099",
 -7593 => x"C0C0C0BFF89290B0",
 -7592 => x"C0C0C0BFF89290A4",
 -7591 => x"C0C0C0BFF89290F9",
 -7590 => x"C0C0C0BFF89290C0",
 -7589 => x"C0C0C0BFF8928090",
 -7588 => x"C0C0C0BFF8928080",
 -7587 => x"C0C0C0BFF89280F8",
 -7586 => x"C0C0C0BFF8928082",
 -7585 => x"C0C0C0BFF8928092",
 -7584 => x"C0C0C0BFF8928099",
 -7583 => x"C0C0C0BFF89280B0",
 -7582 => x"C0C0C0BFF89280A4",
 -7581 => x"C0C0C0BFF89280F9",
 -7580 => x"C0C0C0BFF89280C0",
 -7579 => x"C0C0C0BFF892F890",
 -7578 => x"C0C0C0BFF892F880",
 -7577 => x"C0C0C0BFF892F8F8",
 -7576 => x"C0C0C0BFF892F882",
 -7575 => x"C0C0C0BFF892F892",
 -7574 => x"C0C0C0BFF892F899",
 -7573 => x"C0C0C0BFF892F8B0",
 -7572 => x"C0C0C0BFF892F8A4",
 -7571 => x"C0C0C0BFF892F8F9",
 -7570 => x"C0C0C0BFF892F8C0",
 -7569 => x"C0C0C0BFF8928290",
 -7568 => x"C0C0C0BFF8928280",
 -7567 => x"C0C0C0BFF89282F8",
 -7566 => x"C0C0C0BFF8928282",
 -7565 => x"C0C0C0BFF8928292",
 -7564 => x"C0C0C0BFF8928299",
 -7563 => x"C0C0C0BFF89282B0",
 -7562 => x"C0C0C0BFF89282A4",
 -7561 => x"C0C0C0BFF89282F9",
 -7560 => x"C0C0C0BFF89282C0",
 -7559 => x"C0C0C0BFF8929290",
 -7558 => x"C0C0C0BFF8929280",
 -7557 => x"C0C0C0BFF89292F8",
 -7556 => x"C0C0C0BFF8929282",
 -7555 => x"C0C0C0BFF8929292",
 -7554 => x"C0C0C0BFF8929299",
 -7553 => x"C0C0C0BFF89292B0",
 -7552 => x"C0C0C0BFF89292A4",
 -7551 => x"C0C0C0BFF89292F9",
 -7550 => x"C0C0C0BFF89292C0",
 -7549 => x"C0C0C0BFF8929990",
 -7548 => x"C0C0C0BFF8929980",
 -7547 => x"C0C0C0BFF89299F8",
 -7546 => x"C0C0C0BFF8929982",
 -7545 => x"C0C0C0BFF8929992",
 -7544 => x"C0C0C0BFF8929999",
 -7543 => x"C0C0C0BFF89299B0",
 -7542 => x"C0C0C0BFF89299A4",
 -7541 => x"C0C0C0BFF89299F9",
 -7540 => x"C0C0C0BFF89299C0",
 -7539 => x"C0C0C0BFF892B090",
 -7538 => x"C0C0C0BFF892B080",
 -7537 => x"C0C0C0BFF892B0F8",
 -7536 => x"C0C0C0BFF892B082",
 -7535 => x"C0C0C0BFF892B092",
 -7534 => x"C0C0C0BFF892B099",
 -7533 => x"C0C0C0BFF892B0B0",
 -7532 => x"C0C0C0BFF892B0A4",
 -7531 => x"C0C0C0BFF892B0F9",
 -7530 => x"C0C0C0BFF892B0C0",
 -7529 => x"C0C0C0BFF892A490",
 -7528 => x"C0C0C0BFF892A480",
 -7527 => x"C0C0C0BFF892A4F8",
 -7526 => x"C0C0C0BFF892A482",
 -7525 => x"C0C0C0BFF892A492",
 -7524 => x"C0C0C0BFF892A499",
 -7523 => x"C0C0C0BFF892A4B0",
 -7522 => x"C0C0C0BFF892A4A4",
 -7521 => x"C0C0C0BFF892A4F9",
 -7520 => x"C0C0C0BFF892A4C0",
 -7519 => x"C0C0C0BFF892F990",
 -7518 => x"C0C0C0BFF892F980",
 -7517 => x"C0C0C0BFF892F9F8",
 -7516 => x"C0C0C0BFF892F982",
 -7515 => x"C0C0C0BFF892F992",
 -7514 => x"C0C0C0BFF892F999",
 -7513 => x"C0C0C0BFF892F9B0",
 -7512 => x"C0C0C0BFF892F9A4",
 -7511 => x"C0C0C0BFF892F9F9",
 -7510 => x"C0C0C0BFF892F9C0",
 -7509 => x"C0C0C0BFF892C090",
 -7508 => x"C0C0C0BFF892C080",
 -7507 => x"C0C0C0BFF892C0F8",
 -7506 => x"C0C0C0BFF892C082",
 -7505 => x"C0C0C0BFF892C092",
 -7504 => x"C0C0C0BFF892C099",
 -7503 => x"C0C0C0BFF892C0B0",
 -7502 => x"C0C0C0BFF892C0A4",
 -7501 => x"C0C0C0BFF892C0F9",
 -7500 => x"C0C0C0BFF892C0C0",
 -7499 => x"C0C0C0BFF8999090",
 -7498 => x"C0C0C0BFF8999080",
 -7497 => x"C0C0C0BFF89990F8",
 -7496 => x"C0C0C0BFF8999082",
 -7495 => x"C0C0C0BFF8999092",
 -7494 => x"C0C0C0BFF8999099",
 -7493 => x"C0C0C0BFF89990B0",
 -7492 => x"C0C0C0BFF89990A4",
 -7491 => x"C0C0C0BFF89990F9",
 -7490 => x"C0C0C0BFF89990C0",
 -7489 => x"C0C0C0BFF8998090",
 -7488 => x"C0C0C0BFF8998080",
 -7487 => x"C0C0C0BFF89980F8",
 -7486 => x"C0C0C0BFF8998082",
 -7485 => x"C0C0C0BFF8998092",
 -7484 => x"C0C0C0BFF8998099",
 -7483 => x"C0C0C0BFF89980B0",
 -7482 => x"C0C0C0BFF89980A4",
 -7481 => x"C0C0C0BFF89980F9",
 -7480 => x"C0C0C0BFF89980C0",
 -7479 => x"C0C0C0BFF899F890",
 -7478 => x"C0C0C0BFF899F880",
 -7477 => x"C0C0C0BFF899F8F8",
 -7476 => x"C0C0C0BFF899F882",
 -7475 => x"C0C0C0BFF899F892",
 -7474 => x"C0C0C0BFF899F899",
 -7473 => x"C0C0C0BFF899F8B0",
 -7472 => x"C0C0C0BFF899F8A4",
 -7471 => x"C0C0C0BFF899F8F9",
 -7470 => x"C0C0C0BFF899F8C0",
 -7469 => x"C0C0C0BFF8998290",
 -7468 => x"C0C0C0BFF8998280",
 -7467 => x"C0C0C0BFF89982F8",
 -7466 => x"C0C0C0BFF8998282",
 -7465 => x"C0C0C0BFF8998292",
 -7464 => x"C0C0C0BFF8998299",
 -7463 => x"C0C0C0BFF89982B0",
 -7462 => x"C0C0C0BFF89982A4",
 -7461 => x"C0C0C0BFF89982F9",
 -7460 => x"C0C0C0BFF89982C0",
 -7459 => x"C0C0C0BFF8999290",
 -7458 => x"C0C0C0BFF8999280",
 -7457 => x"C0C0C0BFF89992F8",
 -7456 => x"C0C0C0BFF8999282",
 -7455 => x"C0C0C0BFF8999292",
 -7454 => x"C0C0C0BFF8999299",
 -7453 => x"C0C0C0BFF89992B0",
 -7452 => x"C0C0C0BFF89992A4",
 -7451 => x"C0C0C0BFF89992F9",
 -7450 => x"C0C0C0BFF89992C0",
 -7449 => x"C0C0C0BFF8999990",
 -7448 => x"C0C0C0BFF8999980",
 -7447 => x"C0C0C0BFF89999F8",
 -7446 => x"C0C0C0BFF8999982",
 -7445 => x"C0C0C0BFF8999992",
 -7444 => x"C0C0C0BFF8999999",
 -7443 => x"C0C0C0BFF89999B0",
 -7442 => x"C0C0C0BFF89999A4",
 -7441 => x"C0C0C0BFF89999F9",
 -7440 => x"C0C0C0BFF89999C0",
 -7439 => x"C0C0C0BFF899B090",
 -7438 => x"C0C0C0BFF899B080",
 -7437 => x"C0C0C0BFF899B0F8",
 -7436 => x"C0C0C0BFF899B082",
 -7435 => x"C0C0C0BFF899B092",
 -7434 => x"C0C0C0BFF899B099",
 -7433 => x"C0C0C0BFF899B0B0",
 -7432 => x"C0C0C0BFF899B0A4",
 -7431 => x"C0C0C0BFF899B0F9",
 -7430 => x"C0C0C0BFF899B0C0",
 -7429 => x"C0C0C0BFF899A490",
 -7428 => x"C0C0C0BFF899A480",
 -7427 => x"C0C0C0BFF899A4F8",
 -7426 => x"C0C0C0BFF899A482",
 -7425 => x"C0C0C0BFF899A492",
 -7424 => x"C0C0C0BFF899A499",
 -7423 => x"C0C0C0BFF899A4B0",
 -7422 => x"C0C0C0BFF899A4A4",
 -7421 => x"C0C0C0BFF899A4F9",
 -7420 => x"C0C0C0BFF899A4C0",
 -7419 => x"C0C0C0BFF899F990",
 -7418 => x"C0C0C0BFF899F980",
 -7417 => x"C0C0C0BFF899F9F8",
 -7416 => x"C0C0C0BFF899F982",
 -7415 => x"C0C0C0BFF899F992",
 -7414 => x"C0C0C0BFF899F999",
 -7413 => x"C0C0C0BFF899F9B0",
 -7412 => x"C0C0C0BFF899F9A4",
 -7411 => x"C0C0C0BFF899F9F9",
 -7410 => x"C0C0C0BFF899F9C0",
 -7409 => x"C0C0C0BFF899C090",
 -7408 => x"C0C0C0BFF899C080",
 -7407 => x"C0C0C0BFF899C0F8",
 -7406 => x"C0C0C0BFF899C082",
 -7405 => x"C0C0C0BFF899C092",
 -7404 => x"C0C0C0BFF899C099",
 -7403 => x"C0C0C0BFF899C0B0",
 -7402 => x"C0C0C0BFF899C0A4",
 -7401 => x"C0C0C0BFF899C0F9",
 -7400 => x"C0C0C0BFF899C0C0",
 -7399 => x"C0C0C0BFF8B09090",
 -7398 => x"C0C0C0BFF8B09080",
 -7397 => x"C0C0C0BFF8B090F8",
 -7396 => x"C0C0C0BFF8B09082",
 -7395 => x"C0C0C0BFF8B09092",
 -7394 => x"C0C0C0BFF8B09099",
 -7393 => x"C0C0C0BFF8B090B0",
 -7392 => x"C0C0C0BFF8B090A4",
 -7391 => x"C0C0C0BFF8B090F9",
 -7390 => x"C0C0C0BFF8B090C0",
 -7389 => x"C0C0C0BFF8B08090",
 -7388 => x"C0C0C0BFF8B08080",
 -7387 => x"C0C0C0BFF8B080F8",
 -7386 => x"C0C0C0BFF8B08082",
 -7385 => x"C0C0C0BFF8B08092",
 -7384 => x"C0C0C0BFF8B08099",
 -7383 => x"C0C0C0BFF8B080B0",
 -7382 => x"C0C0C0BFF8B080A4",
 -7381 => x"C0C0C0BFF8B080F9",
 -7380 => x"C0C0C0BFF8B080C0",
 -7379 => x"C0C0C0BFF8B0F890",
 -7378 => x"C0C0C0BFF8B0F880",
 -7377 => x"C0C0C0BFF8B0F8F8",
 -7376 => x"C0C0C0BFF8B0F882",
 -7375 => x"C0C0C0BFF8B0F892",
 -7374 => x"C0C0C0BFF8B0F899",
 -7373 => x"C0C0C0BFF8B0F8B0",
 -7372 => x"C0C0C0BFF8B0F8A4",
 -7371 => x"C0C0C0BFF8B0F8F9",
 -7370 => x"C0C0C0BFF8B0F8C0",
 -7369 => x"C0C0C0BFF8B08290",
 -7368 => x"C0C0C0BFF8B08280",
 -7367 => x"C0C0C0BFF8B082F8",
 -7366 => x"C0C0C0BFF8B08282",
 -7365 => x"C0C0C0BFF8B08292",
 -7364 => x"C0C0C0BFF8B08299",
 -7363 => x"C0C0C0BFF8B082B0",
 -7362 => x"C0C0C0BFF8B082A4",
 -7361 => x"C0C0C0BFF8B082F9",
 -7360 => x"C0C0C0BFF8B082C0",
 -7359 => x"C0C0C0BFF8B09290",
 -7358 => x"C0C0C0BFF8B09280",
 -7357 => x"C0C0C0BFF8B092F8",
 -7356 => x"C0C0C0BFF8B09282",
 -7355 => x"C0C0C0BFF8B09292",
 -7354 => x"C0C0C0BFF8B09299",
 -7353 => x"C0C0C0BFF8B092B0",
 -7352 => x"C0C0C0BFF8B092A4",
 -7351 => x"C0C0C0BFF8B092F9",
 -7350 => x"C0C0C0BFF8B092C0",
 -7349 => x"C0C0C0BFF8B09990",
 -7348 => x"C0C0C0BFF8B09980",
 -7347 => x"C0C0C0BFF8B099F8",
 -7346 => x"C0C0C0BFF8B09982",
 -7345 => x"C0C0C0BFF8B09992",
 -7344 => x"C0C0C0BFF8B09999",
 -7343 => x"C0C0C0BFF8B099B0",
 -7342 => x"C0C0C0BFF8B099A4",
 -7341 => x"C0C0C0BFF8B099F9",
 -7340 => x"C0C0C0BFF8B099C0",
 -7339 => x"C0C0C0BFF8B0B090",
 -7338 => x"C0C0C0BFF8B0B080",
 -7337 => x"C0C0C0BFF8B0B0F8",
 -7336 => x"C0C0C0BFF8B0B082",
 -7335 => x"C0C0C0BFF8B0B092",
 -7334 => x"C0C0C0BFF8B0B099",
 -7333 => x"C0C0C0BFF8B0B0B0",
 -7332 => x"C0C0C0BFF8B0B0A4",
 -7331 => x"C0C0C0BFF8B0B0F9",
 -7330 => x"C0C0C0BFF8B0B0C0",
 -7329 => x"C0C0C0BFF8B0A490",
 -7328 => x"C0C0C0BFF8B0A480",
 -7327 => x"C0C0C0BFF8B0A4F8",
 -7326 => x"C0C0C0BFF8B0A482",
 -7325 => x"C0C0C0BFF8B0A492",
 -7324 => x"C0C0C0BFF8B0A499",
 -7323 => x"C0C0C0BFF8B0A4B0",
 -7322 => x"C0C0C0BFF8B0A4A4",
 -7321 => x"C0C0C0BFF8B0A4F9",
 -7320 => x"C0C0C0BFF8B0A4C0",
 -7319 => x"C0C0C0BFF8B0F990",
 -7318 => x"C0C0C0BFF8B0F980",
 -7317 => x"C0C0C0BFF8B0F9F8",
 -7316 => x"C0C0C0BFF8B0F982",
 -7315 => x"C0C0C0BFF8B0F992",
 -7314 => x"C0C0C0BFF8B0F999",
 -7313 => x"C0C0C0BFF8B0F9B0",
 -7312 => x"C0C0C0BFF8B0F9A4",
 -7311 => x"C0C0C0BFF8B0F9F9",
 -7310 => x"C0C0C0BFF8B0F9C0",
 -7309 => x"C0C0C0BFF8B0C090",
 -7308 => x"C0C0C0BFF8B0C080",
 -7307 => x"C0C0C0BFF8B0C0F8",
 -7306 => x"C0C0C0BFF8B0C082",
 -7305 => x"C0C0C0BFF8B0C092",
 -7304 => x"C0C0C0BFF8B0C099",
 -7303 => x"C0C0C0BFF8B0C0B0",
 -7302 => x"C0C0C0BFF8B0C0A4",
 -7301 => x"C0C0C0BFF8B0C0F9",
 -7300 => x"C0C0C0BFF8B0C0C0",
 -7299 => x"C0C0C0BFF8A49090",
 -7298 => x"C0C0C0BFF8A49080",
 -7297 => x"C0C0C0BFF8A490F8",
 -7296 => x"C0C0C0BFF8A49082",
 -7295 => x"C0C0C0BFF8A49092",
 -7294 => x"C0C0C0BFF8A49099",
 -7293 => x"C0C0C0BFF8A490B0",
 -7292 => x"C0C0C0BFF8A490A4",
 -7291 => x"C0C0C0BFF8A490F9",
 -7290 => x"C0C0C0BFF8A490C0",
 -7289 => x"C0C0C0BFF8A48090",
 -7288 => x"C0C0C0BFF8A48080",
 -7287 => x"C0C0C0BFF8A480F8",
 -7286 => x"C0C0C0BFF8A48082",
 -7285 => x"C0C0C0BFF8A48092",
 -7284 => x"C0C0C0BFF8A48099",
 -7283 => x"C0C0C0BFF8A480B0",
 -7282 => x"C0C0C0BFF8A480A4",
 -7281 => x"C0C0C0BFF8A480F9",
 -7280 => x"C0C0C0BFF8A480C0",
 -7279 => x"C0C0C0BFF8A4F890",
 -7278 => x"C0C0C0BFF8A4F880",
 -7277 => x"C0C0C0BFF8A4F8F8",
 -7276 => x"C0C0C0BFF8A4F882",
 -7275 => x"C0C0C0BFF8A4F892",
 -7274 => x"C0C0C0BFF8A4F899",
 -7273 => x"C0C0C0BFF8A4F8B0",
 -7272 => x"C0C0C0BFF8A4F8A4",
 -7271 => x"C0C0C0BFF8A4F8F9",
 -7270 => x"C0C0C0BFF8A4F8C0",
 -7269 => x"C0C0C0BFF8A48290",
 -7268 => x"C0C0C0BFF8A48280",
 -7267 => x"C0C0C0BFF8A482F8",
 -7266 => x"C0C0C0BFF8A48282",
 -7265 => x"C0C0C0BFF8A48292",
 -7264 => x"C0C0C0BFF8A48299",
 -7263 => x"C0C0C0BFF8A482B0",
 -7262 => x"C0C0C0BFF8A482A4",
 -7261 => x"C0C0C0BFF8A482F9",
 -7260 => x"C0C0C0BFF8A482C0",
 -7259 => x"C0C0C0BFF8A49290",
 -7258 => x"C0C0C0BFF8A49280",
 -7257 => x"C0C0C0BFF8A492F8",
 -7256 => x"C0C0C0BFF8A49282",
 -7255 => x"C0C0C0BFF8A49292",
 -7254 => x"C0C0C0BFF8A49299",
 -7253 => x"C0C0C0BFF8A492B0",
 -7252 => x"C0C0C0BFF8A492A4",
 -7251 => x"C0C0C0BFF8A492F9",
 -7250 => x"C0C0C0BFF8A492C0",
 -7249 => x"C0C0C0BFF8A49990",
 -7248 => x"C0C0C0BFF8A49980",
 -7247 => x"C0C0C0BFF8A499F8",
 -7246 => x"C0C0C0BFF8A49982",
 -7245 => x"C0C0C0BFF8A49992",
 -7244 => x"C0C0C0BFF8A49999",
 -7243 => x"C0C0C0BFF8A499B0",
 -7242 => x"C0C0C0BFF8A499A4",
 -7241 => x"C0C0C0BFF8A499F9",
 -7240 => x"C0C0C0BFF8A499C0",
 -7239 => x"C0C0C0BFF8A4B090",
 -7238 => x"C0C0C0BFF8A4B080",
 -7237 => x"C0C0C0BFF8A4B0F8",
 -7236 => x"C0C0C0BFF8A4B082",
 -7235 => x"C0C0C0BFF8A4B092",
 -7234 => x"C0C0C0BFF8A4B099",
 -7233 => x"C0C0C0BFF8A4B0B0",
 -7232 => x"C0C0C0BFF8A4B0A4",
 -7231 => x"C0C0C0BFF8A4B0F9",
 -7230 => x"C0C0C0BFF8A4B0C0",
 -7229 => x"C0C0C0BFF8A4A490",
 -7228 => x"C0C0C0BFF8A4A480",
 -7227 => x"C0C0C0BFF8A4A4F8",
 -7226 => x"C0C0C0BFF8A4A482",
 -7225 => x"C0C0C0BFF8A4A492",
 -7224 => x"C0C0C0BFF8A4A499",
 -7223 => x"C0C0C0BFF8A4A4B0",
 -7222 => x"C0C0C0BFF8A4A4A4",
 -7221 => x"C0C0C0BFF8A4A4F9",
 -7220 => x"C0C0C0BFF8A4A4C0",
 -7219 => x"C0C0C0BFF8A4F990",
 -7218 => x"C0C0C0BFF8A4F980",
 -7217 => x"C0C0C0BFF8A4F9F8",
 -7216 => x"C0C0C0BFF8A4F982",
 -7215 => x"C0C0C0BFF8A4F992",
 -7214 => x"C0C0C0BFF8A4F999",
 -7213 => x"C0C0C0BFF8A4F9B0",
 -7212 => x"C0C0C0BFF8A4F9A4",
 -7211 => x"C0C0C0BFF8A4F9F9",
 -7210 => x"C0C0C0BFF8A4F9C0",
 -7209 => x"C0C0C0BFF8A4C090",
 -7208 => x"C0C0C0BFF8A4C080",
 -7207 => x"C0C0C0BFF8A4C0F8",
 -7206 => x"C0C0C0BFF8A4C082",
 -7205 => x"C0C0C0BFF8A4C092",
 -7204 => x"C0C0C0BFF8A4C099",
 -7203 => x"C0C0C0BFF8A4C0B0",
 -7202 => x"C0C0C0BFF8A4C0A4",
 -7201 => x"C0C0C0BFF8A4C0F9",
 -7200 => x"C0C0C0BFF8A4C0C0",
 -7199 => x"C0C0C0BFF8F99090",
 -7198 => x"C0C0C0BFF8F99080",
 -7197 => x"C0C0C0BFF8F990F8",
 -7196 => x"C0C0C0BFF8F99082",
 -7195 => x"C0C0C0BFF8F99092",
 -7194 => x"C0C0C0BFF8F99099",
 -7193 => x"C0C0C0BFF8F990B0",
 -7192 => x"C0C0C0BFF8F990A4",
 -7191 => x"C0C0C0BFF8F990F9",
 -7190 => x"C0C0C0BFF8F990C0",
 -7189 => x"C0C0C0BFF8F98090",
 -7188 => x"C0C0C0BFF8F98080",
 -7187 => x"C0C0C0BFF8F980F8",
 -7186 => x"C0C0C0BFF8F98082",
 -7185 => x"C0C0C0BFF8F98092",
 -7184 => x"C0C0C0BFF8F98099",
 -7183 => x"C0C0C0BFF8F980B0",
 -7182 => x"C0C0C0BFF8F980A4",
 -7181 => x"C0C0C0BFF8F980F9",
 -7180 => x"C0C0C0BFF8F980C0",
 -7179 => x"C0C0C0BFF8F9F890",
 -7178 => x"C0C0C0BFF8F9F880",
 -7177 => x"C0C0C0BFF8F9F8F8",
 -7176 => x"C0C0C0BFF8F9F882",
 -7175 => x"C0C0C0BFF8F9F892",
 -7174 => x"C0C0C0BFF8F9F899",
 -7173 => x"C0C0C0BFF8F9F8B0",
 -7172 => x"C0C0C0BFF8F9F8A4",
 -7171 => x"C0C0C0BFF8F9F8F9",
 -7170 => x"C0C0C0BFF8F9F8C0",
 -7169 => x"C0C0C0BFF8F98290",
 -7168 => x"C0C0C0BFF8F98280",
 -7167 => x"C0C0C0BFF8F982F8",
 -7166 => x"C0C0C0BFF8F98282",
 -7165 => x"C0C0C0BFF8F98292",
 -7164 => x"C0C0C0BFF8F98299",
 -7163 => x"C0C0C0BFF8F982B0",
 -7162 => x"C0C0C0BFF8F982A4",
 -7161 => x"C0C0C0BFF8F982F9",
 -7160 => x"C0C0C0BFF8F982C0",
 -7159 => x"C0C0C0BFF8F99290",
 -7158 => x"C0C0C0BFF8F99280",
 -7157 => x"C0C0C0BFF8F992F8",
 -7156 => x"C0C0C0BFF8F99282",
 -7155 => x"C0C0C0BFF8F99292",
 -7154 => x"C0C0C0BFF8F99299",
 -7153 => x"C0C0C0BFF8F992B0",
 -7152 => x"C0C0C0BFF8F992A4",
 -7151 => x"C0C0C0BFF8F992F9",
 -7150 => x"C0C0C0BFF8F992C0",
 -7149 => x"C0C0C0BFF8F99990",
 -7148 => x"C0C0C0BFF8F99980",
 -7147 => x"C0C0C0BFF8F999F8",
 -7146 => x"C0C0C0BFF8F99982",
 -7145 => x"C0C0C0BFF8F99992",
 -7144 => x"C0C0C0BFF8F99999",
 -7143 => x"C0C0C0BFF8F999B0",
 -7142 => x"C0C0C0BFF8F999A4",
 -7141 => x"C0C0C0BFF8F999F9",
 -7140 => x"C0C0C0BFF8F999C0",
 -7139 => x"C0C0C0BFF8F9B090",
 -7138 => x"C0C0C0BFF8F9B080",
 -7137 => x"C0C0C0BFF8F9B0F8",
 -7136 => x"C0C0C0BFF8F9B082",
 -7135 => x"C0C0C0BFF8F9B092",
 -7134 => x"C0C0C0BFF8F9B099",
 -7133 => x"C0C0C0BFF8F9B0B0",
 -7132 => x"C0C0C0BFF8F9B0A4",
 -7131 => x"C0C0C0BFF8F9B0F9",
 -7130 => x"C0C0C0BFF8F9B0C0",
 -7129 => x"C0C0C0BFF8F9A490",
 -7128 => x"C0C0C0BFF8F9A480",
 -7127 => x"C0C0C0BFF8F9A4F8",
 -7126 => x"C0C0C0BFF8F9A482",
 -7125 => x"C0C0C0BFF8F9A492",
 -7124 => x"C0C0C0BFF8F9A499",
 -7123 => x"C0C0C0BFF8F9A4B0",
 -7122 => x"C0C0C0BFF8F9A4A4",
 -7121 => x"C0C0C0BFF8F9A4F9",
 -7120 => x"C0C0C0BFF8F9A4C0",
 -7119 => x"C0C0C0BFF8F9F990",
 -7118 => x"C0C0C0BFF8F9F980",
 -7117 => x"C0C0C0BFF8F9F9F8",
 -7116 => x"C0C0C0BFF8F9F982",
 -7115 => x"C0C0C0BFF8F9F992",
 -7114 => x"C0C0C0BFF8F9F999",
 -7113 => x"C0C0C0BFF8F9F9B0",
 -7112 => x"C0C0C0BFF8F9F9A4",
 -7111 => x"C0C0C0BFF8F9F9F9",
 -7110 => x"C0C0C0BFF8F9F9C0",
 -7109 => x"C0C0C0BFF8F9C090",
 -7108 => x"C0C0C0BFF8F9C080",
 -7107 => x"C0C0C0BFF8F9C0F8",
 -7106 => x"C0C0C0BFF8F9C082",
 -7105 => x"C0C0C0BFF8F9C092",
 -7104 => x"C0C0C0BFF8F9C099",
 -7103 => x"C0C0C0BFF8F9C0B0",
 -7102 => x"C0C0C0BFF8F9C0A4",
 -7101 => x"C0C0C0BFF8F9C0F9",
 -7100 => x"C0C0C0BFF8F9C0C0",
 -7099 => x"C0C0C0BFF8C09090",
 -7098 => x"C0C0C0BFF8C09080",
 -7097 => x"C0C0C0BFF8C090F8",
 -7096 => x"C0C0C0BFF8C09082",
 -7095 => x"C0C0C0BFF8C09092",
 -7094 => x"C0C0C0BFF8C09099",
 -7093 => x"C0C0C0BFF8C090B0",
 -7092 => x"C0C0C0BFF8C090A4",
 -7091 => x"C0C0C0BFF8C090F9",
 -7090 => x"C0C0C0BFF8C090C0",
 -7089 => x"C0C0C0BFF8C08090",
 -7088 => x"C0C0C0BFF8C08080",
 -7087 => x"C0C0C0BFF8C080F8",
 -7086 => x"C0C0C0BFF8C08082",
 -7085 => x"C0C0C0BFF8C08092",
 -7084 => x"C0C0C0BFF8C08099",
 -7083 => x"C0C0C0BFF8C080B0",
 -7082 => x"C0C0C0BFF8C080A4",
 -7081 => x"C0C0C0BFF8C080F9",
 -7080 => x"C0C0C0BFF8C080C0",
 -7079 => x"C0C0C0BFF8C0F890",
 -7078 => x"C0C0C0BFF8C0F880",
 -7077 => x"C0C0C0BFF8C0F8F8",
 -7076 => x"C0C0C0BFF8C0F882",
 -7075 => x"C0C0C0BFF8C0F892",
 -7074 => x"C0C0C0BFF8C0F899",
 -7073 => x"C0C0C0BFF8C0F8B0",
 -7072 => x"C0C0C0BFF8C0F8A4",
 -7071 => x"C0C0C0BFF8C0F8F9",
 -7070 => x"C0C0C0BFF8C0F8C0",
 -7069 => x"C0C0C0BFF8C08290",
 -7068 => x"C0C0C0BFF8C08280",
 -7067 => x"C0C0C0BFF8C082F8",
 -7066 => x"C0C0C0BFF8C08282",
 -7065 => x"C0C0C0BFF8C08292",
 -7064 => x"C0C0C0BFF8C08299",
 -7063 => x"C0C0C0BFF8C082B0",
 -7062 => x"C0C0C0BFF8C082A4",
 -7061 => x"C0C0C0BFF8C082F9",
 -7060 => x"C0C0C0BFF8C082C0",
 -7059 => x"C0C0C0BFF8C09290",
 -7058 => x"C0C0C0BFF8C09280",
 -7057 => x"C0C0C0BFF8C092F8",
 -7056 => x"C0C0C0BFF8C09282",
 -7055 => x"C0C0C0BFF8C09292",
 -7054 => x"C0C0C0BFF8C09299",
 -7053 => x"C0C0C0BFF8C092B0",
 -7052 => x"C0C0C0BFF8C092A4",
 -7051 => x"C0C0C0BFF8C092F9",
 -7050 => x"C0C0C0BFF8C092C0",
 -7049 => x"C0C0C0BFF8C09990",
 -7048 => x"C0C0C0BFF8C09980",
 -7047 => x"C0C0C0BFF8C099F8",
 -7046 => x"C0C0C0BFF8C09982",
 -7045 => x"C0C0C0BFF8C09992",
 -7044 => x"C0C0C0BFF8C09999",
 -7043 => x"C0C0C0BFF8C099B0",
 -7042 => x"C0C0C0BFF8C099A4",
 -7041 => x"C0C0C0BFF8C099F9",
 -7040 => x"C0C0C0BFF8C099C0",
 -7039 => x"C0C0C0BFF8C0B090",
 -7038 => x"C0C0C0BFF8C0B080",
 -7037 => x"C0C0C0BFF8C0B0F8",
 -7036 => x"C0C0C0BFF8C0B082",
 -7035 => x"C0C0C0BFF8C0B092",
 -7034 => x"C0C0C0BFF8C0B099",
 -7033 => x"C0C0C0BFF8C0B0B0",
 -7032 => x"C0C0C0BFF8C0B0A4",
 -7031 => x"C0C0C0BFF8C0B0F9",
 -7030 => x"C0C0C0BFF8C0B0C0",
 -7029 => x"C0C0C0BFF8C0A490",
 -7028 => x"C0C0C0BFF8C0A480",
 -7027 => x"C0C0C0BFF8C0A4F8",
 -7026 => x"C0C0C0BFF8C0A482",
 -7025 => x"C0C0C0BFF8C0A492",
 -7024 => x"C0C0C0BFF8C0A499",
 -7023 => x"C0C0C0BFF8C0A4B0",
 -7022 => x"C0C0C0BFF8C0A4A4",
 -7021 => x"C0C0C0BFF8C0A4F9",
 -7020 => x"C0C0C0BFF8C0A4C0",
 -7019 => x"C0C0C0BFF8C0F990",
 -7018 => x"C0C0C0BFF8C0F980",
 -7017 => x"C0C0C0BFF8C0F9F8",
 -7016 => x"C0C0C0BFF8C0F982",
 -7015 => x"C0C0C0BFF8C0F992",
 -7014 => x"C0C0C0BFF8C0F999",
 -7013 => x"C0C0C0BFF8C0F9B0",
 -7012 => x"C0C0C0BFF8C0F9A4",
 -7011 => x"C0C0C0BFF8C0F9F9",
 -7010 => x"C0C0C0BFF8C0F9C0",
 -7009 => x"C0C0C0BFF8C0C090",
 -7008 => x"C0C0C0BFF8C0C080",
 -7007 => x"C0C0C0BFF8C0C0F8",
 -7006 => x"C0C0C0BFF8C0C082",
 -7005 => x"C0C0C0BFF8C0C092",
 -7004 => x"C0C0C0BFF8C0C099",
 -7003 => x"C0C0C0BFF8C0C0B0",
 -7002 => x"C0C0C0BFF8C0C0A4",
 -7001 => x"C0C0C0BFF8C0C0F9",
 -7000 => x"C0C0C0BFF8C0C0C0",
 -6999 => x"C0C0C0BF82909090",
 -6998 => x"C0C0C0BF82909080",
 -6997 => x"C0C0C0BF829090F8",
 -6996 => x"C0C0C0BF82909082",
 -6995 => x"C0C0C0BF82909092",
 -6994 => x"C0C0C0BF82909099",
 -6993 => x"C0C0C0BF829090B0",
 -6992 => x"C0C0C0BF829090A4",
 -6991 => x"C0C0C0BF829090F9",
 -6990 => x"C0C0C0BF829090C0",
 -6989 => x"C0C0C0BF82908090",
 -6988 => x"C0C0C0BF82908080",
 -6987 => x"C0C0C0BF829080F8",
 -6986 => x"C0C0C0BF82908082",
 -6985 => x"C0C0C0BF82908092",
 -6984 => x"C0C0C0BF82908099",
 -6983 => x"C0C0C0BF829080B0",
 -6982 => x"C0C0C0BF829080A4",
 -6981 => x"C0C0C0BF829080F9",
 -6980 => x"C0C0C0BF829080C0",
 -6979 => x"C0C0C0BF8290F890",
 -6978 => x"C0C0C0BF8290F880",
 -6977 => x"C0C0C0BF8290F8F8",
 -6976 => x"C0C0C0BF8290F882",
 -6975 => x"C0C0C0BF8290F892",
 -6974 => x"C0C0C0BF8290F899",
 -6973 => x"C0C0C0BF8290F8B0",
 -6972 => x"C0C0C0BF8290F8A4",
 -6971 => x"C0C0C0BF8290F8F9",
 -6970 => x"C0C0C0BF8290F8C0",
 -6969 => x"C0C0C0BF82908290",
 -6968 => x"C0C0C0BF82908280",
 -6967 => x"C0C0C0BF829082F8",
 -6966 => x"C0C0C0BF82908282",
 -6965 => x"C0C0C0BF82908292",
 -6964 => x"C0C0C0BF82908299",
 -6963 => x"C0C0C0BF829082B0",
 -6962 => x"C0C0C0BF829082A4",
 -6961 => x"C0C0C0BF829082F9",
 -6960 => x"C0C0C0BF829082C0",
 -6959 => x"C0C0C0BF82909290",
 -6958 => x"C0C0C0BF82909280",
 -6957 => x"C0C0C0BF829092F8",
 -6956 => x"C0C0C0BF82909282",
 -6955 => x"C0C0C0BF82909292",
 -6954 => x"C0C0C0BF82909299",
 -6953 => x"C0C0C0BF829092B0",
 -6952 => x"C0C0C0BF829092A4",
 -6951 => x"C0C0C0BF829092F9",
 -6950 => x"C0C0C0BF829092C0",
 -6949 => x"C0C0C0BF82909990",
 -6948 => x"C0C0C0BF82909980",
 -6947 => x"C0C0C0BF829099F8",
 -6946 => x"C0C0C0BF82909982",
 -6945 => x"C0C0C0BF82909992",
 -6944 => x"C0C0C0BF82909999",
 -6943 => x"C0C0C0BF829099B0",
 -6942 => x"C0C0C0BF829099A4",
 -6941 => x"C0C0C0BF829099F9",
 -6940 => x"C0C0C0BF829099C0",
 -6939 => x"C0C0C0BF8290B090",
 -6938 => x"C0C0C0BF8290B080",
 -6937 => x"C0C0C0BF8290B0F8",
 -6936 => x"C0C0C0BF8290B082",
 -6935 => x"C0C0C0BF8290B092",
 -6934 => x"C0C0C0BF8290B099",
 -6933 => x"C0C0C0BF8290B0B0",
 -6932 => x"C0C0C0BF8290B0A4",
 -6931 => x"C0C0C0BF8290B0F9",
 -6930 => x"C0C0C0BF8290B0C0",
 -6929 => x"C0C0C0BF8290A490",
 -6928 => x"C0C0C0BF8290A480",
 -6927 => x"C0C0C0BF8290A4F8",
 -6926 => x"C0C0C0BF8290A482",
 -6925 => x"C0C0C0BF8290A492",
 -6924 => x"C0C0C0BF8290A499",
 -6923 => x"C0C0C0BF8290A4B0",
 -6922 => x"C0C0C0BF8290A4A4",
 -6921 => x"C0C0C0BF8290A4F9",
 -6920 => x"C0C0C0BF8290A4C0",
 -6919 => x"C0C0C0BF8290F990",
 -6918 => x"C0C0C0BF8290F980",
 -6917 => x"C0C0C0BF8290F9F8",
 -6916 => x"C0C0C0BF8290F982",
 -6915 => x"C0C0C0BF8290F992",
 -6914 => x"C0C0C0BF8290F999",
 -6913 => x"C0C0C0BF8290F9B0",
 -6912 => x"C0C0C0BF8290F9A4",
 -6911 => x"C0C0C0BF8290F9F9",
 -6910 => x"C0C0C0BF8290F9C0",
 -6909 => x"C0C0C0BF8290C090",
 -6908 => x"C0C0C0BF8290C080",
 -6907 => x"C0C0C0BF8290C0F8",
 -6906 => x"C0C0C0BF8290C082",
 -6905 => x"C0C0C0BF8290C092",
 -6904 => x"C0C0C0BF8290C099",
 -6903 => x"C0C0C0BF8290C0B0",
 -6902 => x"C0C0C0BF8290C0A4",
 -6901 => x"C0C0C0BF8290C0F9",
 -6900 => x"C0C0C0BF8290C0C0",
 -6899 => x"C0C0C0BF82809090",
 -6898 => x"C0C0C0BF82809080",
 -6897 => x"C0C0C0BF828090F8",
 -6896 => x"C0C0C0BF82809082",
 -6895 => x"C0C0C0BF82809092",
 -6894 => x"C0C0C0BF82809099",
 -6893 => x"C0C0C0BF828090B0",
 -6892 => x"C0C0C0BF828090A4",
 -6891 => x"C0C0C0BF828090F9",
 -6890 => x"C0C0C0BF828090C0",
 -6889 => x"C0C0C0BF82808090",
 -6888 => x"C0C0C0BF82808080",
 -6887 => x"C0C0C0BF828080F8",
 -6886 => x"C0C0C0BF82808082",
 -6885 => x"C0C0C0BF82808092",
 -6884 => x"C0C0C0BF82808099",
 -6883 => x"C0C0C0BF828080B0",
 -6882 => x"C0C0C0BF828080A4",
 -6881 => x"C0C0C0BF828080F9",
 -6880 => x"C0C0C0BF828080C0",
 -6879 => x"C0C0C0BF8280F890",
 -6878 => x"C0C0C0BF8280F880",
 -6877 => x"C0C0C0BF8280F8F8",
 -6876 => x"C0C0C0BF8280F882",
 -6875 => x"C0C0C0BF8280F892",
 -6874 => x"C0C0C0BF8280F899",
 -6873 => x"C0C0C0BF8280F8B0",
 -6872 => x"C0C0C0BF8280F8A4",
 -6871 => x"C0C0C0BF8280F8F9",
 -6870 => x"C0C0C0BF8280F8C0",
 -6869 => x"C0C0C0BF82808290",
 -6868 => x"C0C0C0BF82808280",
 -6867 => x"C0C0C0BF828082F8",
 -6866 => x"C0C0C0BF82808282",
 -6865 => x"C0C0C0BF82808292",
 -6864 => x"C0C0C0BF82808299",
 -6863 => x"C0C0C0BF828082B0",
 -6862 => x"C0C0C0BF828082A4",
 -6861 => x"C0C0C0BF828082F9",
 -6860 => x"C0C0C0BF828082C0",
 -6859 => x"C0C0C0BF82809290",
 -6858 => x"C0C0C0BF82809280",
 -6857 => x"C0C0C0BF828092F8",
 -6856 => x"C0C0C0BF82809282",
 -6855 => x"C0C0C0BF82809292",
 -6854 => x"C0C0C0BF82809299",
 -6853 => x"C0C0C0BF828092B0",
 -6852 => x"C0C0C0BF828092A4",
 -6851 => x"C0C0C0BF828092F9",
 -6850 => x"C0C0C0BF828092C0",
 -6849 => x"C0C0C0BF82809990",
 -6848 => x"C0C0C0BF82809980",
 -6847 => x"C0C0C0BF828099F8",
 -6846 => x"C0C0C0BF82809982",
 -6845 => x"C0C0C0BF82809992",
 -6844 => x"C0C0C0BF82809999",
 -6843 => x"C0C0C0BF828099B0",
 -6842 => x"C0C0C0BF828099A4",
 -6841 => x"C0C0C0BF828099F9",
 -6840 => x"C0C0C0BF828099C0",
 -6839 => x"C0C0C0BF8280B090",
 -6838 => x"C0C0C0BF8280B080",
 -6837 => x"C0C0C0BF8280B0F8",
 -6836 => x"C0C0C0BF8280B082",
 -6835 => x"C0C0C0BF8280B092",
 -6834 => x"C0C0C0BF8280B099",
 -6833 => x"C0C0C0BF8280B0B0",
 -6832 => x"C0C0C0BF8280B0A4",
 -6831 => x"C0C0C0BF8280B0F9",
 -6830 => x"C0C0C0BF8280B0C0",
 -6829 => x"C0C0C0BF8280A490",
 -6828 => x"C0C0C0BF8280A480",
 -6827 => x"C0C0C0BF8280A4F8",
 -6826 => x"C0C0C0BF8280A482",
 -6825 => x"C0C0C0BF8280A492",
 -6824 => x"C0C0C0BF8280A499",
 -6823 => x"C0C0C0BF8280A4B0",
 -6822 => x"C0C0C0BF8280A4A4",
 -6821 => x"C0C0C0BF8280A4F9",
 -6820 => x"C0C0C0BF8280A4C0",
 -6819 => x"C0C0C0BF8280F990",
 -6818 => x"C0C0C0BF8280F980",
 -6817 => x"C0C0C0BF8280F9F8",
 -6816 => x"C0C0C0BF8280F982",
 -6815 => x"C0C0C0BF8280F992",
 -6814 => x"C0C0C0BF8280F999",
 -6813 => x"C0C0C0BF8280F9B0",
 -6812 => x"C0C0C0BF8280F9A4",
 -6811 => x"C0C0C0BF8280F9F9",
 -6810 => x"C0C0C0BF8280F9C0",
 -6809 => x"C0C0C0BF8280C090",
 -6808 => x"C0C0C0BF8280C080",
 -6807 => x"C0C0C0BF8280C0F8",
 -6806 => x"C0C0C0BF8280C082",
 -6805 => x"C0C0C0BF8280C092",
 -6804 => x"C0C0C0BF8280C099",
 -6803 => x"C0C0C0BF8280C0B0",
 -6802 => x"C0C0C0BF8280C0A4",
 -6801 => x"C0C0C0BF8280C0F9",
 -6800 => x"C0C0C0BF8280C0C0",
 -6799 => x"C0C0C0BF82F89090",
 -6798 => x"C0C0C0BF82F89080",
 -6797 => x"C0C0C0BF82F890F8",
 -6796 => x"C0C0C0BF82F89082",
 -6795 => x"C0C0C0BF82F89092",
 -6794 => x"C0C0C0BF82F89099",
 -6793 => x"C0C0C0BF82F890B0",
 -6792 => x"C0C0C0BF82F890A4",
 -6791 => x"C0C0C0BF82F890F9",
 -6790 => x"C0C0C0BF82F890C0",
 -6789 => x"C0C0C0BF82F88090",
 -6788 => x"C0C0C0BF82F88080",
 -6787 => x"C0C0C0BF82F880F8",
 -6786 => x"C0C0C0BF82F88082",
 -6785 => x"C0C0C0BF82F88092",
 -6784 => x"C0C0C0BF82F88099",
 -6783 => x"C0C0C0BF82F880B0",
 -6782 => x"C0C0C0BF82F880A4",
 -6781 => x"C0C0C0BF82F880F9",
 -6780 => x"C0C0C0BF82F880C0",
 -6779 => x"C0C0C0BF82F8F890",
 -6778 => x"C0C0C0BF82F8F880",
 -6777 => x"C0C0C0BF82F8F8F8",
 -6776 => x"C0C0C0BF82F8F882",
 -6775 => x"C0C0C0BF82F8F892",
 -6774 => x"C0C0C0BF82F8F899",
 -6773 => x"C0C0C0BF82F8F8B0",
 -6772 => x"C0C0C0BF82F8F8A4",
 -6771 => x"C0C0C0BF82F8F8F9",
 -6770 => x"C0C0C0BF82F8F8C0",
 -6769 => x"C0C0C0BF82F88290",
 -6768 => x"C0C0C0BF82F88280",
 -6767 => x"C0C0C0BF82F882F8",
 -6766 => x"C0C0C0BF82F88282",
 -6765 => x"C0C0C0BF82F88292",
 -6764 => x"C0C0C0BF82F88299",
 -6763 => x"C0C0C0BF82F882B0",
 -6762 => x"C0C0C0BF82F882A4",
 -6761 => x"C0C0C0BF82F882F9",
 -6760 => x"C0C0C0BF82F882C0",
 -6759 => x"C0C0C0BF82F89290",
 -6758 => x"C0C0C0BF82F89280",
 -6757 => x"C0C0C0BF82F892F8",
 -6756 => x"C0C0C0BF82F89282",
 -6755 => x"C0C0C0BF82F89292",
 -6754 => x"C0C0C0BF82F89299",
 -6753 => x"C0C0C0BF82F892B0",
 -6752 => x"C0C0C0BF82F892A4",
 -6751 => x"C0C0C0BF82F892F9",
 -6750 => x"C0C0C0BF82F892C0",
 -6749 => x"C0C0C0BF82F89990",
 -6748 => x"C0C0C0BF82F89980",
 -6747 => x"C0C0C0BF82F899F8",
 -6746 => x"C0C0C0BF82F89982",
 -6745 => x"C0C0C0BF82F89992",
 -6744 => x"C0C0C0BF82F89999",
 -6743 => x"C0C0C0BF82F899B0",
 -6742 => x"C0C0C0BF82F899A4",
 -6741 => x"C0C0C0BF82F899F9",
 -6740 => x"C0C0C0BF82F899C0",
 -6739 => x"C0C0C0BF82F8B090",
 -6738 => x"C0C0C0BF82F8B080",
 -6737 => x"C0C0C0BF82F8B0F8",
 -6736 => x"C0C0C0BF82F8B082",
 -6735 => x"C0C0C0BF82F8B092",
 -6734 => x"C0C0C0BF82F8B099",
 -6733 => x"C0C0C0BF82F8B0B0",
 -6732 => x"C0C0C0BF82F8B0A4",
 -6731 => x"C0C0C0BF82F8B0F9",
 -6730 => x"C0C0C0BF82F8B0C0",
 -6729 => x"C0C0C0BF82F8A490",
 -6728 => x"C0C0C0BF82F8A480",
 -6727 => x"C0C0C0BF82F8A4F8",
 -6726 => x"C0C0C0BF82F8A482",
 -6725 => x"C0C0C0BF82F8A492",
 -6724 => x"C0C0C0BF82F8A499",
 -6723 => x"C0C0C0BF82F8A4B0",
 -6722 => x"C0C0C0BF82F8A4A4",
 -6721 => x"C0C0C0BF82F8A4F9",
 -6720 => x"C0C0C0BF82F8A4C0",
 -6719 => x"C0C0C0BF82F8F990",
 -6718 => x"C0C0C0BF82F8F980",
 -6717 => x"C0C0C0BF82F8F9F8",
 -6716 => x"C0C0C0BF82F8F982",
 -6715 => x"C0C0C0BF82F8F992",
 -6714 => x"C0C0C0BF82F8F999",
 -6713 => x"C0C0C0BF82F8F9B0",
 -6712 => x"C0C0C0BF82F8F9A4",
 -6711 => x"C0C0C0BF82F8F9F9",
 -6710 => x"C0C0C0BF82F8F9C0",
 -6709 => x"C0C0C0BF82F8C090",
 -6708 => x"C0C0C0BF82F8C080",
 -6707 => x"C0C0C0BF82F8C0F8",
 -6706 => x"C0C0C0BF82F8C082",
 -6705 => x"C0C0C0BF82F8C092",
 -6704 => x"C0C0C0BF82F8C099",
 -6703 => x"C0C0C0BF82F8C0B0",
 -6702 => x"C0C0C0BF82F8C0A4",
 -6701 => x"C0C0C0BF82F8C0F9",
 -6700 => x"C0C0C0BF82F8C0C0",
 -6699 => x"C0C0C0BF82829090",
 -6698 => x"C0C0C0BF82829080",
 -6697 => x"C0C0C0BF828290F8",
 -6696 => x"C0C0C0BF82829082",
 -6695 => x"C0C0C0BF82829092",
 -6694 => x"C0C0C0BF82829099",
 -6693 => x"C0C0C0BF828290B0",
 -6692 => x"C0C0C0BF828290A4",
 -6691 => x"C0C0C0BF828290F9",
 -6690 => x"C0C0C0BF828290C0",
 -6689 => x"C0C0C0BF82828090",
 -6688 => x"C0C0C0BF82828080",
 -6687 => x"C0C0C0BF828280F8",
 -6686 => x"C0C0C0BF82828082",
 -6685 => x"C0C0C0BF82828092",
 -6684 => x"C0C0C0BF82828099",
 -6683 => x"C0C0C0BF828280B0",
 -6682 => x"C0C0C0BF828280A4",
 -6681 => x"C0C0C0BF828280F9",
 -6680 => x"C0C0C0BF828280C0",
 -6679 => x"C0C0C0BF8282F890",
 -6678 => x"C0C0C0BF8282F880",
 -6677 => x"C0C0C0BF8282F8F8",
 -6676 => x"C0C0C0BF8282F882",
 -6675 => x"C0C0C0BF8282F892",
 -6674 => x"C0C0C0BF8282F899",
 -6673 => x"C0C0C0BF8282F8B0",
 -6672 => x"C0C0C0BF8282F8A4",
 -6671 => x"C0C0C0BF8282F8F9",
 -6670 => x"C0C0C0BF8282F8C0",
 -6669 => x"C0C0C0BF82828290",
 -6668 => x"C0C0C0BF82828280",
 -6667 => x"C0C0C0BF828282F8",
 -6666 => x"C0C0C0BF82828282",
 -6665 => x"C0C0C0BF82828292",
 -6664 => x"C0C0C0BF82828299",
 -6663 => x"C0C0C0BF828282B0",
 -6662 => x"C0C0C0BF828282A4",
 -6661 => x"C0C0C0BF828282F9",
 -6660 => x"C0C0C0BF828282C0",
 -6659 => x"C0C0C0BF82829290",
 -6658 => x"C0C0C0BF82829280",
 -6657 => x"C0C0C0BF828292F8",
 -6656 => x"C0C0C0BF82829282",
 -6655 => x"C0C0C0BF82829292",
 -6654 => x"C0C0C0BF82829299",
 -6653 => x"C0C0C0BF828292B0",
 -6652 => x"C0C0C0BF828292A4",
 -6651 => x"C0C0C0BF828292F9",
 -6650 => x"C0C0C0BF828292C0",
 -6649 => x"C0C0C0BF82829990",
 -6648 => x"C0C0C0BF82829980",
 -6647 => x"C0C0C0BF828299F8",
 -6646 => x"C0C0C0BF82829982",
 -6645 => x"C0C0C0BF82829992",
 -6644 => x"C0C0C0BF82829999",
 -6643 => x"C0C0C0BF828299B0",
 -6642 => x"C0C0C0BF828299A4",
 -6641 => x"C0C0C0BF828299F9",
 -6640 => x"C0C0C0BF828299C0",
 -6639 => x"C0C0C0BF8282B090",
 -6638 => x"C0C0C0BF8282B080",
 -6637 => x"C0C0C0BF8282B0F8",
 -6636 => x"C0C0C0BF8282B082",
 -6635 => x"C0C0C0BF8282B092",
 -6634 => x"C0C0C0BF8282B099",
 -6633 => x"C0C0C0BF8282B0B0",
 -6632 => x"C0C0C0BF8282B0A4",
 -6631 => x"C0C0C0BF8282B0F9",
 -6630 => x"C0C0C0BF8282B0C0",
 -6629 => x"C0C0C0BF8282A490",
 -6628 => x"C0C0C0BF8282A480",
 -6627 => x"C0C0C0BF8282A4F8",
 -6626 => x"C0C0C0BF8282A482",
 -6625 => x"C0C0C0BF8282A492",
 -6624 => x"C0C0C0BF8282A499",
 -6623 => x"C0C0C0BF8282A4B0",
 -6622 => x"C0C0C0BF8282A4A4",
 -6621 => x"C0C0C0BF8282A4F9",
 -6620 => x"C0C0C0BF8282A4C0",
 -6619 => x"C0C0C0BF8282F990",
 -6618 => x"C0C0C0BF8282F980",
 -6617 => x"C0C0C0BF8282F9F8",
 -6616 => x"C0C0C0BF8282F982",
 -6615 => x"C0C0C0BF8282F992",
 -6614 => x"C0C0C0BF8282F999",
 -6613 => x"C0C0C0BF8282F9B0",
 -6612 => x"C0C0C0BF8282F9A4",
 -6611 => x"C0C0C0BF8282F9F9",
 -6610 => x"C0C0C0BF8282F9C0",
 -6609 => x"C0C0C0BF8282C090",
 -6608 => x"C0C0C0BF8282C080",
 -6607 => x"C0C0C0BF8282C0F8",
 -6606 => x"C0C0C0BF8282C082",
 -6605 => x"C0C0C0BF8282C092",
 -6604 => x"C0C0C0BF8282C099",
 -6603 => x"C0C0C0BF8282C0B0",
 -6602 => x"C0C0C0BF8282C0A4",
 -6601 => x"C0C0C0BF8282C0F9",
 -6600 => x"C0C0C0BF8282C0C0",
 -6599 => x"C0C0C0BF82929090",
 -6598 => x"C0C0C0BF82929080",
 -6597 => x"C0C0C0BF829290F8",
 -6596 => x"C0C0C0BF82929082",
 -6595 => x"C0C0C0BF82929092",
 -6594 => x"C0C0C0BF82929099",
 -6593 => x"C0C0C0BF829290B0",
 -6592 => x"C0C0C0BF829290A4",
 -6591 => x"C0C0C0BF829290F9",
 -6590 => x"C0C0C0BF829290C0",
 -6589 => x"C0C0C0BF82928090",
 -6588 => x"C0C0C0BF82928080",
 -6587 => x"C0C0C0BF829280F8",
 -6586 => x"C0C0C0BF82928082",
 -6585 => x"C0C0C0BF82928092",
 -6584 => x"C0C0C0BF82928099",
 -6583 => x"C0C0C0BF829280B0",
 -6582 => x"C0C0C0BF829280A4",
 -6581 => x"C0C0C0BF829280F9",
 -6580 => x"C0C0C0BF829280C0",
 -6579 => x"C0C0C0BF8292F890",
 -6578 => x"C0C0C0BF8292F880",
 -6577 => x"C0C0C0BF8292F8F8",
 -6576 => x"C0C0C0BF8292F882",
 -6575 => x"C0C0C0BF8292F892",
 -6574 => x"C0C0C0BF8292F899",
 -6573 => x"C0C0C0BF8292F8B0",
 -6572 => x"C0C0C0BF8292F8A4",
 -6571 => x"C0C0C0BF8292F8F9",
 -6570 => x"C0C0C0BF8292F8C0",
 -6569 => x"C0C0C0BF82928290",
 -6568 => x"C0C0C0BF82928280",
 -6567 => x"C0C0C0BF829282F8",
 -6566 => x"C0C0C0BF82928282",
 -6565 => x"C0C0C0BF82928292",
 -6564 => x"C0C0C0BF82928299",
 -6563 => x"C0C0C0BF829282B0",
 -6562 => x"C0C0C0BF829282A4",
 -6561 => x"C0C0C0BF829282F9",
 -6560 => x"C0C0C0BF829282C0",
 -6559 => x"C0C0C0BF82929290",
 -6558 => x"C0C0C0BF82929280",
 -6557 => x"C0C0C0BF829292F8",
 -6556 => x"C0C0C0BF82929282",
 -6555 => x"C0C0C0BF82929292",
 -6554 => x"C0C0C0BF82929299",
 -6553 => x"C0C0C0BF829292B0",
 -6552 => x"C0C0C0BF829292A4",
 -6551 => x"C0C0C0BF829292F9",
 -6550 => x"C0C0C0BF829292C0",
 -6549 => x"C0C0C0BF82929990",
 -6548 => x"C0C0C0BF82929980",
 -6547 => x"C0C0C0BF829299F8",
 -6546 => x"C0C0C0BF82929982",
 -6545 => x"C0C0C0BF82929992",
 -6544 => x"C0C0C0BF82929999",
 -6543 => x"C0C0C0BF829299B0",
 -6542 => x"C0C0C0BF829299A4",
 -6541 => x"C0C0C0BF829299F9",
 -6540 => x"C0C0C0BF829299C0",
 -6539 => x"C0C0C0BF8292B090",
 -6538 => x"C0C0C0BF8292B080",
 -6537 => x"C0C0C0BF8292B0F8",
 -6536 => x"C0C0C0BF8292B082",
 -6535 => x"C0C0C0BF8292B092",
 -6534 => x"C0C0C0BF8292B099",
 -6533 => x"C0C0C0BF8292B0B0",
 -6532 => x"C0C0C0BF8292B0A4",
 -6531 => x"C0C0C0BF8292B0F9",
 -6530 => x"C0C0C0BF8292B0C0",
 -6529 => x"C0C0C0BF8292A490",
 -6528 => x"C0C0C0BF8292A480",
 -6527 => x"C0C0C0BF8292A4F8",
 -6526 => x"C0C0C0BF8292A482",
 -6525 => x"C0C0C0BF8292A492",
 -6524 => x"C0C0C0BF8292A499",
 -6523 => x"C0C0C0BF8292A4B0",
 -6522 => x"C0C0C0BF8292A4A4",
 -6521 => x"C0C0C0BF8292A4F9",
 -6520 => x"C0C0C0BF8292A4C0",
 -6519 => x"C0C0C0BF8292F990",
 -6518 => x"C0C0C0BF8292F980",
 -6517 => x"C0C0C0BF8292F9F8",
 -6516 => x"C0C0C0BF8292F982",
 -6515 => x"C0C0C0BF8292F992",
 -6514 => x"C0C0C0BF8292F999",
 -6513 => x"C0C0C0BF8292F9B0",
 -6512 => x"C0C0C0BF8292F9A4",
 -6511 => x"C0C0C0BF8292F9F9",
 -6510 => x"C0C0C0BF8292F9C0",
 -6509 => x"C0C0C0BF8292C090",
 -6508 => x"C0C0C0BF8292C080",
 -6507 => x"C0C0C0BF8292C0F8",
 -6506 => x"C0C0C0BF8292C082",
 -6505 => x"C0C0C0BF8292C092",
 -6504 => x"C0C0C0BF8292C099",
 -6503 => x"C0C0C0BF8292C0B0",
 -6502 => x"C0C0C0BF8292C0A4",
 -6501 => x"C0C0C0BF8292C0F9",
 -6500 => x"C0C0C0BF8292C0C0",
 -6499 => x"C0C0C0BF82999090",
 -6498 => x"C0C0C0BF82999080",
 -6497 => x"C0C0C0BF829990F8",
 -6496 => x"C0C0C0BF82999082",
 -6495 => x"C0C0C0BF82999092",
 -6494 => x"C0C0C0BF82999099",
 -6493 => x"C0C0C0BF829990B0",
 -6492 => x"C0C0C0BF829990A4",
 -6491 => x"C0C0C0BF829990F9",
 -6490 => x"C0C0C0BF829990C0",
 -6489 => x"C0C0C0BF82998090",
 -6488 => x"C0C0C0BF82998080",
 -6487 => x"C0C0C0BF829980F8",
 -6486 => x"C0C0C0BF82998082",
 -6485 => x"C0C0C0BF82998092",
 -6484 => x"C0C0C0BF82998099",
 -6483 => x"C0C0C0BF829980B0",
 -6482 => x"C0C0C0BF829980A4",
 -6481 => x"C0C0C0BF829980F9",
 -6480 => x"C0C0C0BF829980C0",
 -6479 => x"C0C0C0BF8299F890",
 -6478 => x"C0C0C0BF8299F880",
 -6477 => x"C0C0C0BF8299F8F8",
 -6476 => x"C0C0C0BF8299F882",
 -6475 => x"C0C0C0BF8299F892",
 -6474 => x"C0C0C0BF8299F899",
 -6473 => x"C0C0C0BF8299F8B0",
 -6472 => x"C0C0C0BF8299F8A4",
 -6471 => x"C0C0C0BF8299F8F9",
 -6470 => x"C0C0C0BF8299F8C0",
 -6469 => x"C0C0C0BF82998290",
 -6468 => x"C0C0C0BF82998280",
 -6467 => x"C0C0C0BF829982F8",
 -6466 => x"C0C0C0BF82998282",
 -6465 => x"C0C0C0BF82998292",
 -6464 => x"C0C0C0BF82998299",
 -6463 => x"C0C0C0BF829982B0",
 -6462 => x"C0C0C0BF829982A4",
 -6461 => x"C0C0C0BF829982F9",
 -6460 => x"C0C0C0BF829982C0",
 -6459 => x"C0C0C0BF82999290",
 -6458 => x"C0C0C0BF82999280",
 -6457 => x"C0C0C0BF829992F8",
 -6456 => x"C0C0C0BF82999282",
 -6455 => x"C0C0C0BF82999292",
 -6454 => x"C0C0C0BF82999299",
 -6453 => x"C0C0C0BF829992B0",
 -6452 => x"C0C0C0BF829992A4",
 -6451 => x"C0C0C0BF829992F9",
 -6450 => x"C0C0C0BF829992C0",
 -6449 => x"C0C0C0BF82999990",
 -6448 => x"C0C0C0BF82999980",
 -6447 => x"C0C0C0BF829999F8",
 -6446 => x"C0C0C0BF82999982",
 -6445 => x"C0C0C0BF82999992",
 -6444 => x"C0C0C0BF82999999",
 -6443 => x"C0C0C0BF829999B0",
 -6442 => x"C0C0C0BF829999A4",
 -6441 => x"C0C0C0BF829999F9",
 -6440 => x"C0C0C0BF829999C0",
 -6439 => x"C0C0C0BF8299B090",
 -6438 => x"C0C0C0BF8299B080",
 -6437 => x"C0C0C0BF8299B0F8",
 -6436 => x"C0C0C0BF8299B082",
 -6435 => x"C0C0C0BF8299B092",
 -6434 => x"C0C0C0BF8299B099",
 -6433 => x"C0C0C0BF8299B0B0",
 -6432 => x"C0C0C0BF8299B0A4",
 -6431 => x"C0C0C0BF8299B0F9",
 -6430 => x"C0C0C0BF8299B0C0",
 -6429 => x"C0C0C0BF8299A490",
 -6428 => x"C0C0C0BF8299A480",
 -6427 => x"C0C0C0BF8299A4F8",
 -6426 => x"C0C0C0BF8299A482",
 -6425 => x"C0C0C0BF8299A492",
 -6424 => x"C0C0C0BF8299A499",
 -6423 => x"C0C0C0BF8299A4B0",
 -6422 => x"C0C0C0BF8299A4A4",
 -6421 => x"C0C0C0BF8299A4F9",
 -6420 => x"C0C0C0BF8299A4C0",
 -6419 => x"C0C0C0BF8299F990",
 -6418 => x"C0C0C0BF8299F980",
 -6417 => x"C0C0C0BF8299F9F8",
 -6416 => x"C0C0C0BF8299F982",
 -6415 => x"C0C0C0BF8299F992",
 -6414 => x"C0C0C0BF8299F999",
 -6413 => x"C0C0C0BF8299F9B0",
 -6412 => x"C0C0C0BF8299F9A4",
 -6411 => x"C0C0C0BF8299F9F9",
 -6410 => x"C0C0C0BF8299F9C0",
 -6409 => x"C0C0C0BF8299C090",
 -6408 => x"C0C0C0BF8299C080",
 -6407 => x"C0C0C0BF8299C0F8",
 -6406 => x"C0C0C0BF8299C082",
 -6405 => x"C0C0C0BF8299C092",
 -6404 => x"C0C0C0BF8299C099",
 -6403 => x"C0C0C0BF8299C0B0",
 -6402 => x"C0C0C0BF8299C0A4",
 -6401 => x"C0C0C0BF8299C0F9",
 -6400 => x"C0C0C0BF8299C0C0",
 -6399 => x"C0C0C0BF82B09090",
 -6398 => x"C0C0C0BF82B09080",
 -6397 => x"C0C0C0BF82B090F8",
 -6396 => x"C0C0C0BF82B09082",
 -6395 => x"C0C0C0BF82B09092",
 -6394 => x"C0C0C0BF82B09099",
 -6393 => x"C0C0C0BF82B090B0",
 -6392 => x"C0C0C0BF82B090A4",
 -6391 => x"C0C0C0BF82B090F9",
 -6390 => x"C0C0C0BF82B090C0",
 -6389 => x"C0C0C0BF82B08090",
 -6388 => x"C0C0C0BF82B08080",
 -6387 => x"C0C0C0BF82B080F8",
 -6386 => x"C0C0C0BF82B08082",
 -6385 => x"C0C0C0BF82B08092",
 -6384 => x"C0C0C0BF82B08099",
 -6383 => x"C0C0C0BF82B080B0",
 -6382 => x"C0C0C0BF82B080A4",
 -6381 => x"C0C0C0BF82B080F9",
 -6380 => x"C0C0C0BF82B080C0",
 -6379 => x"C0C0C0BF82B0F890",
 -6378 => x"C0C0C0BF82B0F880",
 -6377 => x"C0C0C0BF82B0F8F8",
 -6376 => x"C0C0C0BF82B0F882",
 -6375 => x"C0C0C0BF82B0F892",
 -6374 => x"C0C0C0BF82B0F899",
 -6373 => x"C0C0C0BF82B0F8B0",
 -6372 => x"C0C0C0BF82B0F8A4",
 -6371 => x"C0C0C0BF82B0F8F9",
 -6370 => x"C0C0C0BF82B0F8C0",
 -6369 => x"C0C0C0BF82B08290",
 -6368 => x"C0C0C0BF82B08280",
 -6367 => x"C0C0C0BF82B082F8",
 -6366 => x"C0C0C0BF82B08282",
 -6365 => x"C0C0C0BF82B08292",
 -6364 => x"C0C0C0BF82B08299",
 -6363 => x"C0C0C0BF82B082B0",
 -6362 => x"C0C0C0BF82B082A4",
 -6361 => x"C0C0C0BF82B082F9",
 -6360 => x"C0C0C0BF82B082C0",
 -6359 => x"C0C0C0BF82B09290",
 -6358 => x"C0C0C0BF82B09280",
 -6357 => x"C0C0C0BF82B092F8",
 -6356 => x"C0C0C0BF82B09282",
 -6355 => x"C0C0C0BF82B09292",
 -6354 => x"C0C0C0BF82B09299",
 -6353 => x"C0C0C0BF82B092B0",
 -6352 => x"C0C0C0BF82B092A4",
 -6351 => x"C0C0C0BF82B092F9",
 -6350 => x"C0C0C0BF82B092C0",
 -6349 => x"C0C0C0BF82B09990",
 -6348 => x"C0C0C0BF82B09980",
 -6347 => x"C0C0C0BF82B099F8",
 -6346 => x"C0C0C0BF82B09982",
 -6345 => x"C0C0C0BF82B09992",
 -6344 => x"C0C0C0BF82B09999",
 -6343 => x"C0C0C0BF82B099B0",
 -6342 => x"C0C0C0BF82B099A4",
 -6341 => x"C0C0C0BF82B099F9",
 -6340 => x"C0C0C0BF82B099C0",
 -6339 => x"C0C0C0BF82B0B090",
 -6338 => x"C0C0C0BF82B0B080",
 -6337 => x"C0C0C0BF82B0B0F8",
 -6336 => x"C0C0C0BF82B0B082",
 -6335 => x"C0C0C0BF82B0B092",
 -6334 => x"C0C0C0BF82B0B099",
 -6333 => x"C0C0C0BF82B0B0B0",
 -6332 => x"C0C0C0BF82B0B0A4",
 -6331 => x"C0C0C0BF82B0B0F9",
 -6330 => x"C0C0C0BF82B0B0C0",
 -6329 => x"C0C0C0BF82B0A490",
 -6328 => x"C0C0C0BF82B0A480",
 -6327 => x"C0C0C0BF82B0A4F8",
 -6326 => x"C0C0C0BF82B0A482",
 -6325 => x"C0C0C0BF82B0A492",
 -6324 => x"C0C0C0BF82B0A499",
 -6323 => x"C0C0C0BF82B0A4B0",
 -6322 => x"C0C0C0BF82B0A4A4",
 -6321 => x"C0C0C0BF82B0A4F9",
 -6320 => x"C0C0C0BF82B0A4C0",
 -6319 => x"C0C0C0BF82B0F990",
 -6318 => x"C0C0C0BF82B0F980",
 -6317 => x"C0C0C0BF82B0F9F8",
 -6316 => x"C0C0C0BF82B0F982",
 -6315 => x"C0C0C0BF82B0F992",
 -6314 => x"C0C0C0BF82B0F999",
 -6313 => x"C0C0C0BF82B0F9B0",
 -6312 => x"C0C0C0BF82B0F9A4",
 -6311 => x"C0C0C0BF82B0F9F9",
 -6310 => x"C0C0C0BF82B0F9C0",
 -6309 => x"C0C0C0BF82B0C090",
 -6308 => x"C0C0C0BF82B0C080",
 -6307 => x"C0C0C0BF82B0C0F8",
 -6306 => x"C0C0C0BF82B0C082",
 -6305 => x"C0C0C0BF82B0C092",
 -6304 => x"C0C0C0BF82B0C099",
 -6303 => x"C0C0C0BF82B0C0B0",
 -6302 => x"C0C0C0BF82B0C0A4",
 -6301 => x"C0C0C0BF82B0C0F9",
 -6300 => x"C0C0C0BF82B0C0C0",
 -6299 => x"C0C0C0BF82A49090",
 -6298 => x"C0C0C0BF82A49080",
 -6297 => x"C0C0C0BF82A490F8",
 -6296 => x"C0C0C0BF82A49082",
 -6295 => x"C0C0C0BF82A49092",
 -6294 => x"C0C0C0BF82A49099",
 -6293 => x"C0C0C0BF82A490B0",
 -6292 => x"C0C0C0BF82A490A4",
 -6291 => x"C0C0C0BF82A490F9",
 -6290 => x"C0C0C0BF82A490C0",
 -6289 => x"C0C0C0BF82A48090",
 -6288 => x"C0C0C0BF82A48080",
 -6287 => x"C0C0C0BF82A480F8",
 -6286 => x"C0C0C0BF82A48082",
 -6285 => x"C0C0C0BF82A48092",
 -6284 => x"C0C0C0BF82A48099",
 -6283 => x"C0C0C0BF82A480B0",
 -6282 => x"C0C0C0BF82A480A4",
 -6281 => x"C0C0C0BF82A480F9",
 -6280 => x"C0C0C0BF82A480C0",
 -6279 => x"C0C0C0BF82A4F890",
 -6278 => x"C0C0C0BF82A4F880",
 -6277 => x"C0C0C0BF82A4F8F8",
 -6276 => x"C0C0C0BF82A4F882",
 -6275 => x"C0C0C0BF82A4F892",
 -6274 => x"C0C0C0BF82A4F899",
 -6273 => x"C0C0C0BF82A4F8B0",
 -6272 => x"C0C0C0BF82A4F8A4",
 -6271 => x"C0C0C0BF82A4F8F9",
 -6270 => x"C0C0C0BF82A4F8C0",
 -6269 => x"C0C0C0BF82A48290",
 -6268 => x"C0C0C0BF82A48280",
 -6267 => x"C0C0C0BF82A482F8",
 -6266 => x"C0C0C0BF82A48282",
 -6265 => x"C0C0C0BF82A48292",
 -6264 => x"C0C0C0BF82A48299",
 -6263 => x"C0C0C0BF82A482B0",
 -6262 => x"C0C0C0BF82A482A4",
 -6261 => x"C0C0C0BF82A482F9",
 -6260 => x"C0C0C0BF82A482C0",
 -6259 => x"C0C0C0BF82A49290",
 -6258 => x"C0C0C0BF82A49280",
 -6257 => x"C0C0C0BF82A492F8",
 -6256 => x"C0C0C0BF82A49282",
 -6255 => x"C0C0C0BF82A49292",
 -6254 => x"C0C0C0BF82A49299",
 -6253 => x"C0C0C0BF82A492B0",
 -6252 => x"C0C0C0BF82A492A4",
 -6251 => x"C0C0C0BF82A492F9",
 -6250 => x"C0C0C0BF82A492C0",
 -6249 => x"C0C0C0BF82A49990",
 -6248 => x"C0C0C0BF82A49980",
 -6247 => x"C0C0C0BF82A499F8",
 -6246 => x"C0C0C0BF82A49982",
 -6245 => x"C0C0C0BF82A49992",
 -6244 => x"C0C0C0BF82A49999",
 -6243 => x"C0C0C0BF82A499B0",
 -6242 => x"C0C0C0BF82A499A4",
 -6241 => x"C0C0C0BF82A499F9",
 -6240 => x"C0C0C0BF82A499C0",
 -6239 => x"C0C0C0BF82A4B090",
 -6238 => x"C0C0C0BF82A4B080",
 -6237 => x"C0C0C0BF82A4B0F8",
 -6236 => x"C0C0C0BF82A4B082",
 -6235 => x"C0C0C0BF82A4B092",
 -6234 => x"C0C0C0BF82A4B099",
 -6233 => x"C0C0C0BF82A4B0B0",
 -6232 => x"C0C0C0BF82A4B0A4",
 -6231 => x"C0C0C0BF82A4B0F9",
 -6230 => x"C0C0C0BF82A4B0C0",
 -6229 => x"C0C0C0BF82A4A490",
 -6228 => x"C0C0C0BF82A4A480",
 -6227 => x"C0C0C0BF82A4A4F8",
 -6226 => x"C0C0C0BF82A4A482",
 -6225 => x"C0C0C0BF82A4A492",
 -6224 => x"C0C0C0BF82A4A499",
 -6223 => x"C0C0C0BF82A4A4B0",
 -6222 => x"C0C0C0BF82A4A4A4",
 -6221 => x"C0C0C0BF82A4A4F9",
 -6220 => x"C0C0C0BF82A4A4C0",
 -6219 => x"C0C0C0BF82A4F990",
 -6218 => x"C0C0C0BF82A4F980",
 -6217 => x"C0C0C0BF82A4F9F8",
 -6216 => x"C0C0C0BF82A4F982",
 -6215 => x"C0C0C0BF82A4F992",
 -6214 => x"C0C0C0BF82A4F999",
 -6213 => x"C0C0C0BF82A4F9B0",
 -6212 => x"C0C0C0BF82A4F9A4",
 -6211 => x"C0C0C0BF82A4F9F9",
 -6210 => x"C0C0C0BF82A4F9C0",
 -6209 => x"C0C0C0BF82A4C090",
 -6208 => x"C0C0C0BF82A4C080",
 -6207 => x"C0C0C0BF82A4C0F8",
 -6206 => x"C0C0C0BF82A4C082",
 -6205 => x"C0C0C0BF82A4C092",
 -6204 => x"C0C0C0BF82A4C099",
 -6203 => x"C0C0C0BF82A4C0B0",
 -6202 => x"C0C0C0BF82A4C0A4",
 -6201 => x"C0C0C0BF82A4C0F9",
 -6200 => x"C0C0C0BF82A4C0C0",
 -6199 => x"C0C0C0BF82F99090",
 -6198 => x"C0C0C0BF82F99080",
 -6197 => x"C0C0C0BF82F990F8",
 -6196 => x"C0C0C0BF82F99082",
 -6195 => x"C0C0C0BF82F99092",
 -6194 => x"C0C0C0BF82F99099",
 -6193 => x"C0C0C0BF82F990B0",
 -6192 => x"C0C0C0BF82F990A4",
 -6191 => x"C0C0C0BF82F990F9",
 -6190 => x"C0C0C0BF82F990C0",
 -6189 => x"C0C0C0BF82F98090",
 -6188 => x"C0C0C0BF82F98080",
 -6187 => x"C0C0C0BF82F980F8",
 -6186 => x"C0C0C0BF82F98082",
 -6185 => x"C0C0C0BF82F98092",
 -6184 => x"C0C0C0BF82F98099",
 -6183 => x"C0C0C0BF82F980B0",
 -6182 => x"C0C0C0BF82F980A4",
 -6181 => x"C0C0C0BF82F980F9",
 -6180 => x"C0C0C0BF82F980C0",
 -6179 => x"C0C0C0BF82F9F890",
 -6178 => x"C0C0C0BF82F9F880",
 -6177 => x"C0C0C0BF82F9F8F8",
 -6176 => x"C0C0C0BF82F9F882",
 -6175 => x"C0C0C0BF82F9F892",
 -6174 => x"C0C0C0BF82F9F899",
 -6173 => x"C0C0C0BF82F9F8B0",
 -6172 => x"C0C0C0BF82F9F8A4",
 -6171 => x"C0C0C0BF82F9F8F9",
 -6170 => x"C0C0C0BF82F9F8C0",
 -6169 => x"C0C0C0BF82F98290",
 -6168 => x"C0C0C0BF82F98280",
 -6167 => x"C0C0C0BF82F982F8",
 -6166 => x"C0C0C0BF82F98282",
 -6165 => x"C0C0C0BF82F98292",
 -6164 => x"C0C0C0BF82F98299",
 -6163 => x"C0C0C0BF82F982B0",
 -6162 => x"C0C0C0BF82F982A4",
 -6161 => x"C0C0C0BF82F982F9",
 -6160 => x"C0C0C0BF82F982C0",
 -6159 => x"C0C0C0BF82F99290",
 -6158 => x"C0C0C0BF82F99280",
 -6157 => x"C0C0C0BF82F992F8",
 -6156 => x"C0C0C0BF82F99282",
 -6155 => x"C0C0C0BF82F99292",
 -6154 => x"C0C0C0BF82F99299",
 -6153 => x"C0C0C0BF82F992B0",
 -6152 => x"C0C0C0BF82F992A4",
 -6151 => x"C0C0C0BF82F992F9",
 -6150 => x"C0C0C0BF82F992C0",
 -6149 => x"C0C0C0BF82F99990",
 -6148 => x"C0C0C0BF82F99980",
 -6147 => x"C0C0C0BF82F999F8",
 -6146 => x"C0C0C0BF82F99982",
 -6145 => x"C0C0C0BF82F99992",
 -6144 => x"C0C0C0BF82F99999",
 -6143 => x"C0C0C0BF82F999B0",
 -6142 => x"C0C0C0BF82F999A4",
 -6141 => x"C0C0C0BF82F999F9",
 -6140 => x"C0C0C0BF82F999C0",
 -6139 => x"C0C0C0BF82F9B090",
 -6138 => x"C0C0C0BF82F9B080",
 -6137 => x"C0C0C0BF82F9B0F8",
 -6136 => x"C0C0C0BF82F9B082",
 -6135 => x"C0C0C0BF82F9B092",
 -6134 => x"C0C0C0BF82F9B099",
 -6133 => x"C0C0C0BF82F9B0B0",
 -6132 => x"C0C0C0BF82F9B0A4",
 -6131 => x"C0C0C0BF82F9B0F9",
 -6130 => x"C0C0C0BF82F9B0C0",
 -6129 => x"C0C0C0BF82F9A490",
 -6128 => x"C0C0C0BF82F9A480",
 -6127 => x"C0C0C0BF82F9A4F8",
 -6126 => x"C0C0C0BF82F9A482",
 -6125 => x"C0C0C0BF82F9A492",
 -6124 => x"C0C0C0BF82F9A499",
 -6123 => x"C0C0C0BF82F9A4B0",
 -6122 => x"C0C0C0BF82F9A4A4",
 -6121 => x"C0C0C0BF82F9A4F9",
 -6120 => x"C0C0C0BF82F9A4C0",
 -6119 => x"C0C0C0BF82F9F990",
 -6118 => x"C0C0C0BF82F9F980",
 -6117 => x"C0C0C0BF82F9F9F8",
 -6116 => x"C0C0C0BF82F9F982",
 -6115 => x"C0C0C0BF82F9F992",
 -6114 => x"C0C0C0BF82F9F999",
 -6113 => x"C0C0C0BF82F9F9B0",
 -6112 => x"C0C0C0BF82F9F9A4",
 -6111 => x"C0C0C0BF82F9F9F9",
 -6110 => x"C0C0C0BF82F9F9C0",
 -6109 => x"C0C0C0BF82F9C090",
 -6108 => x"C0C0C0BF82F9C080",
 -6107 => x"C0C0C0BF82F9C0F8",
 -6106 => x"C0C0C0BF82F9C082",
 -6105 => x"C0C0C0BF82F9C092",
 -6104 => x"C0C0C0BF82F9C099",
 -6103 => x"C0C0C0BF82F9C0B0",
 -6102 => x"C0C0C0BF82F9C0A4",
 -6101 => x"C0C0C0BF82F9C0F9",
 -6100 => x"C0C0C0BF82F9C0C0",
 -6099 => x"C0C0C0BF82C09090",
 -6098 => x"C0C0C0BF82C09080",
 -6097 => x"C0C0C0BF82C090F8",
 -6096 => x"C0C0C0BF82C09082",
 -6095 => x"C0C0C0BF82C09092",
 -6094 => x"C0C0C0BF82C09099",
 -6093 => x"C0C0C0BF82C090B0",
 -6092 => x"C0C0C0BF82C090A4",
 -6091 => x"C0C0C0BF82C090F9",
 -6090 => x"C0C0C0BF82C090C0",
 -6089 => x"C0C0C0BF82C08090",
 -6088 => x"C0C0C0BF82C08080",
 -6087 => x"C0C0C0BF82C080F8",
 -6086 => x"C0C0C0BF82C08082",
 -6085 => x"C0C0C0BF82C08092",
 -6084 => x"C0C0C0BF82C08099",
 -6083 => x"C0C0C0BF82C080B0",
 -6082 => x"C0C0C0BF82C080A4",
 -6081 => x"C0C0C0BF82C080F9",
 -6080 => x"C0C0C0BF82C080C0",
 -6079 => x"C0C0C0BF82C0F890",
 -6078 => x"C0C0C0BF82C0F880",
 -6077 => x"C0C0C0BF82C0F8F8",
 -6076 => x"C0C0C0BF82C0F882",
 -6075 => x"C0C0C0BF82C0F892",
 -6074 => x"C0C0C0BF82C0F899",
 -6073 => x"C0C0C0BF82C0F8B0",
 -6072 => x"C0C0C0BF82C0F8A4",
 -6071 => x"C0C0C0BF82C0F8F9",
 -6070 => x"C0C0C0BF82C0F8C0",
 -6069 => x"C0C0C0BF82C08290",
 -6068 => x"C0C0C0BF82C08280",
 -6067 => x"C0C0C0BF82C082F8",
 -6066 => x"C0C0C0BF82C08282",
 -6065 => x"C0C0C0BF82C08292",
 -6064 => x"C0C0C0BF82C08299",
 -6063 => x"C0C0C0BF82C082B0",
 -6062 => x"C0C0C0BF82C082A4",
 -6061 => x"C0C0C0BF82C082F9",
 -6060 => x"C0C0C0BF82C082C0",
 -6059 => x"C0C0C0BF82C09290",
 -6058 => x"C0C0C0BF82C09280",
 -6057 => x"C0C0C0BF82C092F8",
 -6056 => x"C0C0C0BF82C09282",
 -6055 => x"C0C0C0BF82C09292",
 -6054 => x"C0C0C0BF82C09299",
 -6053 => x"C0C0C0BF82C092B0",
 -6052 => x"C0C0C0BF82C092A4",
 -6051 => x"C0C0C0BF82C092F9",
 -6050 => x"C0C0C0BF82C092C0",
 -6049 => x"C0C0C0BF82C09990",
 -6048 => x"C0C0C0BF82C09980",
 -6047 => x"C0C0C0BF82C099F8",
 -6046 => x"C0C0C0BF82C09982",
 -6045 => x"C0C0C0BF82C09992",
 -6044 => x"C0C0C0BF82C09999",
 -6043 => x"C0C0C0BF82C099B0",
 -6042 => x"C0C0C0BF82C099A4",
 -6041 => x"C0C0C0BF82C099F9",
 -6040 => x"C0C0C0BF82C099C0",
 -6039 => x"C0C0C0BF82C0B090",
 -6038 => x"C0C0C0BF82C0B080",
 -6037 => x"C0C0C0BF82C0B0F8",
 -6036 => x"C0C0C0BF82C0B082",
 -6035 => x"C0C0C0BF82C0B092",
 -6034 => x"C0C0C0BF82C0B099",
 -6033 => x"C0C0C0BF82C0B0B0",
 -6032 => x"C0C0C0BF82C0B0A4",
 -6031 => x"C0C0C0BF82C0B0F9",
 -6030 => x"C0C0C0BF82C0B0C0",
 -6029 => x"C0C0C0BF82C0A490",
 -6028 => x"C0C0C0BF82C0A480",
 -6027 => x"C0C0C0BF82C0A4F8",
 -6026 => x"C0C0C0BF82C0A482",
 -6025 => x"C0C0C0BF82C0A492",
 -6024 => x"C0C0C0BF82C0A499",
 -6023 => x"C0C0C0BF82C0A4B0",
 -6022 => x"C0C0C0BF82C0A4A4",
 -6021 => x"C0C0C0BF82C0A4F9",
 -6020 => x"C0C0C0BF82C0A4C0",
 -6019 => x"C0C0C0BF82C0F990",
 -6018 => x"C0C0C0BF82C0F980",
 -6017 => x"C0C0C0BF82C0F9F8",
 -6016 => x"C0C0C0BF82C0F982",
 -6015 => x"C0C0C0BF82C0F992",
 -6014 => x"C0C0C0BF82C0F999",
 -6013 => x"C0C0C0BF82C0F9B0",
 -6012 => x"C0C0C0BF82C0F9A4",
 -6011 => x"C0C0C0BF82C0F9F9",
 -6010 => x"C0C0C0BF82C0F9C0",
 -6009 => x"C0C0C0BF82C0C090",
 -6008 => x"C0C0C0BF82C0C080",
 -6007 => x"C0C0C0BF82C0C0F8",
 -6006 => x"C0C0C0BF82C0C082",
 -6005 => x"C0C0C0BF82C0C092",
 -6004 => x"C0C0C0BF82C0C099",
 -6003 => x"C0C0C0BF82C0C0B0",
 -6002 => x"C0C0C0BF82C0C0A4",
 -6001 => x"C0C0C0BF82C0C0F9",
 -6000 => x"C0C0C0BF82C0C0C0",
 -5999 => x"C0C0C0BF92909090",
 -5998 => x"C0C0C0BF92909080",
 -5997 => x"C0C0C0BF929090F8",
 -5996 => x"C0C0C0BF92909082",
 -5995 => x"C0C0C0BF92909092",
 -5994 => x"C0C0C0BF92909099",
 -5993 => x"C0C0C0BF929090B0",
 -5992 => x"C0C0C0BF929090A4",
 -5991 => x"C0C0C0BF929090F9",
 -5990 => x"C0C0C0BF929090C0",
 -5989 => x"C0C0C0BF92908090",
 -5988 => x"C0C0C0BF92908080",
 -5987 => x"C0C0C0BF929080F8",
 -5986 => x"C0C0C0BF92908082",
 -5985 => x"C0C0C0BF92908092",
 -5984 => x"C0C0C0BF92908099",
 -5983 => x"C0C0C0BF929080B0",
 -5982 => x"C0C0C0BF929080A4",
 -5981 => x"C0C0C0BF929080F9",
 -5980 => x"C0C0C0BF929080C0",
 -5979 => x"C0C0C0BF9290F890",
 -5978 => x"C0C0C0BF9290F880",
 -5977 => x"C0C0C0BF9290F8F8",
 -5976 => x"C0C0C0BF9290F882",
 -5975 => x"C0C0C0BF9290F892",
 -5974 => x"C0C0C0BF9290F899",
 -5973 => x"C0C0C0BF9290F8B0",
 -5972 => x"C0C0C0BF9290F8A4",
 -5971 => x"C0C0C0BF9290F8F9",
 -5970 => x"C0C0C0BF9290F8C0",
 -5969 => x"C0C0C0BF92908290",
 -5968 => x"C0C0C0BF92908280",
 -5967 => x"C0C0C0BF929082F8",
 -5966 => x"C0C0C0BF92908282",
 -5965 => x"C0C0C0BF92908292",
 -5964 => x"C0C0C0BF92908299",
 -5963 => x"C0C0C0BF929082B0",
 -5962 => x"C0C0C0BF929082A4",
 -5961 => x"C0C0C0BF929082F9",
 -5960 => x"C0C0C0BF929082C0",
 -5959 => x"C0C0C0BF92909290",
 -5958 => x"C0C0C0BF92909280",
 -5957 => x"C0C0C0BF929092F8",
 -5956 => x"C0C0C0BF92909282",
 -5955 => x"C0C0C0BF92909292",
 -5954 => x"C0C0C0BF92909299",
 -5953 => x"C0C0C0BF929092B0",
 -5952 => x"C0C0C0BF929092A4",
 -5951 => x"C0C0C0BF929092F9",
 -5950 => x"C0C0C0BF929092C0",
 -5949 => x"C0C0C0BF92909990",
 -5948 => x"C0C0C0BF92909980",
 -5947 => x"C0C0C0BF929099F8",
 -5946 => x"C0C0C0BF92909982",
 -5945 => x"C0C0C0BF92909992",
 -5944 => x"C0C0C0BF92909999",
 -5943 => x"C0C0C0BF929099B0",
 -5942 => x"C0C0C0BF929099A4",
 -5941 => x"C0C0C0BF929099F9",
 -5940 => x"C0C0C0BF929099C0",
 -5939 => x"C0C0C0BF9290B090",
 -5938 => x"C0C0C0BF9290B080",
 -5937 => x"C0C0C0BF9290B0F8",
 -5936 => x"C0C0C0BF9290B082",
 -5935 => x"C0C0C0BF9290B092",
 -5934 => x"C0C0C0BF9290B099",
 -5933 => x"C0C0C0BF9290B0B0",
 -5932 => x"C0C0C0BF9290B0A4",
 -5931 => x"C0C0C0BF9290B0F9",
 -5930 => x"C0C0C0BF9290B0C0",
 -5929 => x"C0C0C0BF9290A490",
 -5928 => x"C0C0C0BF9290A480",
 -5927 => x"C0C0C0BF9290A4F8",
 -5926 => x"C0C0C0BF9290A482",
 -5925 => x"C0C0C0BF9290A492",
 -5924 => x"C0C0C0BF9290A499",
 -5923 => x"C0C0C0BF9290A4B0",
 -5922 => x"C0C0C0BF9290A4A4",
 -5921 => x"C0C0C0BF9290A4F9",
 -5920 => x"C0C0C0BF9290A4C0",
 -5919 => x"C0C0C0BF9290F990",
 -5918 => x"C0C0C0BF9290F980",
 -5917 => x"C0C0C0BF9290F9F8",
 -5916 => x"C0C0C0BF9290F982",
 -5915 => x"C0C0C0BF9290F992",
 -5914 => x"C0C0C0BF9290F999",
 -5913 => x"C0C0C0BF9290F9B0",
 -5912 => x"C0C0C0BF9290F9A4",
 -5911 => x"C0C0C0BF9290F9F9",
 -5910 => x"C0C0C0BF9290F9C0",
 -5909 => x"C0C0C0BF9290C090",
 -5908 => x"C0C0C0BF9290C080",
 -5907 => x"C0C0C0BF9290C0F8",
 -5906 => x"C0C0C0BF9290C082",
 -5905 => x"C0C0C0BF9290C092",
 -5904 => x"C0C0C0BF9290C099",
 -5903 => x"C0C0C0BF9290C0B0",
 -5902 => x"C0C0C0BF9290C0A4",
 -5901 => x"C0C0C0BF9290C0F9",
 -5900 => x"C0C0C0BF9290C0C0",
 -5899 => x"C0C0C0BF92809090",
 -5898 => x"C0C0C0BF92809080",
 -5897 => x"C0C0C0BF928090F8",
 -5896 => x"C0C0C0BF92809082",
 -5895 => x"C0C0C0BF92809092",
 -5894 => x"C0C0C0BF92809099",
 -5893 => x"C0C0C0BF928090B0",
 -5892 => x"C0C0C0BF928090A4",
 -5891 => x"C0C0C0BF928090F9",
 -5890 => x"C0C0C0BF928090C0",
 -5889 => x"C0C0C0BF92808090",
 -5888 => x"C0C0C0BF92808080",
 -5887 => x"C0C0C0BF928080F8",
 -5886 => x"C0C0C0BF92808082",
 -5885 => x"C0C0C0BF92808092",
 -5884 => x"C0C0C0BF92808099",
 -5883 => x"C0C0C0BF928080B0",
 -5882 => x"C0C0C0BF928080A4",
 -5881 => x"C0C0C0BF928080F9",
 -5880 => x"C0C0C0BF928080C0",
 -5879 => x"C0C0C0BF9280F890",
 -5878 => x"C0C0C0BF9280F880",
 -5877 => x"C0C0C0BF9280F8F8",
 -5876 => x"C0C0C0BF9280F882",
 -5875 => x"C0C0C0BF9280F892",
 -5874 => x"C0C0C0BF9280F899",
 -5873 => x"C0C0C0BF9280F8B0",
 -5872 => x"C0C0C0BF9280F8A4",
 -5871 => x"C0C0C0BF9280F8F9",
 -5870 => x"C0C0C0BF9280F8C0",
 -5869 => x"C0C0C0BF92808290",
 -5868 => x"C0C0C0BF92808280",
 -5867 => x"C0C0C0BF928082F8",
 -5866 => x"C0C0C0BF92808282",
 -5865 => x"C0C0C0BF92808292",
 -5864 => x"C0C0C0BF92808299",
 -5863 => x"C0C0C0BF928082B0",
 -5862 => x"C0C0C0BF928082A4",
 -5861 => x"C0C0C0BF928082F9",
 -5860 => x"C0C0C0BF928082C0",
 -5859 => x"C0C0C0BF92809290",
 -5858 => x"C0C0C0BF92809280",
 -5857 => x"C0C0C0BF928092F8",
 -5856 => x"C0C0C0BF92809282",
 -5855 => x"C0C0C0BF92809292",
 -5854 => x"C0C0C0BF92809299",
 -5853 => x"C0C0C0BF928092B0",
 -5852 => x"C0C0C0BF928092A4",
 -5851 => x"C0C0C0BF928092F9",
 -5850 => x"C0C0C0BF928092C0",
 -5849 => x"C0C0C0BF92809990",
 -5848 => x"C0C0C0BF92809980",
 -5847 => x"C0C0C0BF928099F8",
 -5846 => x"C0C0C0BF92809982",
 -5845 => x"C0C0C0BF92809992",
 -5844 => x"C0C0C0BF92809999",
 -5843 => x"C0C0C0BF928099B0",
 -5842 => x"C0C0C0BF928099A4",
 -5841 => x"C0C0C0BF928099F9",
 -5840 => x"C0C0C0BF928099C0",
 -5839 => x"C0C0C0BF9280B090",
 -5838 => x"C0C0C0BF9280B080",
 -5837 => x"C0C0C0BF9280B0F8",
 -5836 => x"C0C0C0BF9280B082",
 -5835 => x"C0C0C0BF9280B092",
 -5834 => x"C0C0C0BF9280B099",
 -5833 => x"C0C0C0BF9280B0B0",
 -5832 => x"C0C0C0BF9280B0A4",
 -5831 => x"C0C0C0BF9280B0F9",
 -5830 => x"C0C0C0BF9280B0C0",
 -5829 => x"C0C0C0BF9280A490",
 -5828 => x"C0C0C0BF9280A480",
 -5827 => x"C0C0C0BF9280A4F8",
 -5826 => x"C0C0C0BF9280A482",
 -5825 => x"C0C0C0BF9280A492",
 -5824 => x"C0C0C0BF9280A499",
 -5823 => x"C0C0C0BF9280A4B0",
 -5822 => x"C0C0C0BF9280A4A4",
 -5821 => x"C0C0C0BF9280A4F9",
 -5820 => x"C0C0C0BF9280A4C0",
 -5819 => x"C0C0C0BF9280F990",
 -5818 => x"C0C0C0BF9280F980",
 -5817 => x"C0C0C0BF9280F9F8",
 -5816 => x"C0C0C0BF9280F982",
 -5815 => x"C0C0C0BF9280F992",
 -5814 => x"C0C0C0BF9280F999",
 -5813 => x"C0C0C0BF9280F9B0",
 -5812 => x"C0C0C0BF9280F9A4",
 -5811 => x"C0C0C0BF9280F9F9",
 -5810 => x"C0C0C0BF9280F9C0",
 -5809 => x"C0C0C0BF9280C090",
 -5808 => x"C0C0C0BF9280C080",
 -5807 => x"C0C0C0BF9280C0F8",
 -5806 => x"C0C0C0BF9280C082",
 -5805 => x"C0C0C0BF9280C092",
 -5804 => x"C0C0C0BF9280C099",
 -5803 => x"C0C0C0BF9280C0B0",
 -5802 => x"C0C0C0BF9280C0A4",
 -5801 => x"C0C0C0BF9280C0F9",
 -5800 => x"C0C0C0BF9280C0C0",
 -5799 => x"C0C0C0BF92F89090",
 -5798 => x"C0C0C0BF92F89080",
 -5797 => x"C0C0C0BF92F890F8",
 -5796 => x"C0C0C0BF92F89082",
 -5795 => x"C0C0C0BF92F89092",
 -5794 => x"C0C0C0BF92F89099",
 -5793 => x"C0C0C0BF92F890B0",
 -5792 => x"C0C0C0BF92F890A4",
 -5791 => x"C0C0C0BF92F890F9",
 -5790 => x"C0C0C0BF92F890C0",
 -5789 => x"C0C0C0BF92F88090",
 -5788 => x"C0C0C0BF92F88080",
 -5787 => x"C0C0C0BF92F880F8",
 -5786 => x"C0C0C0BF92F88082",
 -5785 => x"C0C0C0BF92F88092",
 -5784 => x"C0C0C0BF92F88099",
 -5783 => x"C0C0C0BF92F880B0",
 -5782 => x"C0C0C0BF92F880A4",
 -5781 => x"C0C0C0BF92F880F9",
 -5780 => x"C0C0C0BF92F880C0",
 -5779 => x"C0C0C0BF92F8F890",
 -5778 => x"C0C0C0BF92F8F880",
 -5777 => x"C0C0C0BF92F8F8F8",
 -5776 => x"C0C0C0BF92F8F882",
 -5775 => x"C0C0C0BF92F8F892",
 -5774 => x"C0C0C0BF92F8F899",
 -5773 => x"C0C0C0BF92F8F8B0",
 -5772 => x"C0C0C0BF92F8F8A4",
 -5771 => x"C0C0C0BF92F8F8F9",
 -5770 => x"C0C0C0BF92F8F8C0",
 -5769 => x"C0C0C0BF92F88290",
 -5768 => x"C0C0C0BF92F88280",
 -5767 => x"C0C0C0BF92F882F8",
 -5766 => x"C0C0C0BF92F88282",
 -5765 => x"C0C0C0BF92F88292",
 -5764 => x"C0C0C0BF92F88299",
 -5763 => x"C0C0C0BF92F882B0",
 -5762 => x"C0C0C0BF92F882A4",
 -5761 => x"C0C0C0BF92F882F9",
 -5760 => x"C0C0C0BF92F882C0",
 -5759 => x"C0C0C0BF92F89290",
 -5758 => x"C0C0C0BF92F89280",
 -5757 => x"C0C0C0BF92F892F8",
 -5756 => x"C0C0C0BF92F89282",
 -5755 => x"C0C0C0BF92F89292",
 -5754 => x"C0C0C0BF92F89299",
 -5753 => x"C0C0C0BF92F892B0",
 -5752 => x"C0C0C0BF92F892A4",
 -5751 => x"C0C0C0BF92F892F9",
 -5750 => x"C0C0C0BF92F892C0",
 -5749 => x"C0C0C0BF92F89990",
 -5748 => x"C0C0C0BF92F89980",
 -5747 => x"C0C0C0BF92F899F8",
 -5746 => x"C0C0C0BF92F89982",
 -5745 => x"C0C0C0BF92F89992",
 -5744 => x"C0C0C0BF92F89999",
 -5743 => x"C0C0C0BF92F899B0",
 -5742 => x"C0C0C0BF92F899A4",
 -5741 => x"C0C0C0BF92F899F9",
 -5740 => x"C0C0C0BF92F899C0",
 -5739 => x"C0C0C0BF92F8B090",
 -5738 => x"C0C0C0BF92F8B080",
 -5737 => x"C0C0C0BF92F8B0F8",
 -5736 => x"C0C0C0BF92F8B082",
 -5735 => x"C0C0C0BF92F8B092",
 -5734 => x"C0C0C0BF92F8B099",
 -5733 => x"C0C0C0BF92F8B0B0",
 -5732 => x"C0C0C0BF92F8B0A4",
 -5731 => x"C0C0C0BF92F8B0F9",
 -5730 => x"C0C0C0BF92F8B0C0",
 -5729 => x"C0C0C0BF92F8A490",
 -5728 => x"C0C0C0BF92F8A480",
 -5727 => x"C0C0C0BF92F8A4F8",
 -5726 => x"C0C0C0BF92F8A482",
 -5725 => x"C0C0C0BF92F8A492",
 -5724 => x"C0C0C0BF92F8A499",
 -5723 => x"C0C0C0BF92F8A4B0",
 -5722 => x"C0C0C0BF92F8A4A4",
 -5721 => x"C0C0C0BF92F8A4F9",
 -5720 => x"C0C0C0BF92F8A4C0",
 -5719 => x"C0C0C0BF92F8F990",
 -5718 => x"C0C0C0BF92F8F980",
 -5717 => x"C0C0C0BF92F8F9F8",
 -5716 => x"C0C0C0BF92F8F982",
 -5715 => x"C0C0C0BF92F8F992",
 -5714 => x"C0C0C0BF92F8F999",
 -5713 => x"C0C0C0BF92F8F9B0",
 -5712 => x"C0C0C0BF92F8F9A4",
 -5711 => x"C0C0C0BF92F8F9F9",
 -5710 => x"C0C0C0BF92F8F9C0",
 -5709 => x"C0C0C0BF92F8C090",
 -5708 => x"C0C0C0BF92F8C080",
 -5707 => x"C0C0C0BF92F8C0F8",
 -5706 => x"C0C0C0BF92F8C082",
 -5705 => x"C0C0C0BF92F8C092",
 -5704 => x"C0C0C0BF92F8C099",
 -5703 => x"C0C0C0BF92F8C0B0",
 -5702 => x"C0C0C0BF92F8C0A4",
 -5701 => x"C0C0C0BF92F8C0F9",
 -5700 => x"C0C0C0BF92F8C0C0",
 -5699 => x"C0C0C0BF92829090",
 -5698 => x"C0C0C0BF92829080",
 -5697 => x"C0C0C0BF928290F8",
 -5696 => x"C0C0C0BF92829082",
 -5695 => x"C0C0C0BF92829092",
 -5694 => x"C0C0C0BF92829099",
 -5693 => x"C0C0C0BF928290B0",
 -5692 => x"C0C0C0BF928290A4",
 -5691 => x"C0C0C0BF928290F9",
 -5690 => x"C0C0C0BF928290C0",
 -5689 => x"C0C0C0BF92828090",
 -5688 => x"C0C0C0BF92828080",
 -5687 => x"C0C0C0BF928280F8",
 -5686 => x"C0C0C0BF92828082",
 -5685 => x"C0C0C0BF92828092",
 -5684 => x"C0C0C0BF92828099",
 -5683 => x"C0C0C0BF928280B0",
 -5682 => x"C0C0C0BF928280A4",
 -5681 => x"C0C0C0BF928280F9",
 -5680 => x"C0C0C0BF928280C0",
 -5679 => x"C0C0C0BF9282F890",
 -5678 => x"C0C0C0BF9282F880",
 -5677 => x"C0C0C0BF9282F8F8",
 -5676 => x"C0C0C0BF9282F882",
 -5675 => x"C0C0C0BF9282F892",
 -5674 => x"C0C0C0BF9282F899",
 -5673 => x"C0C0C0BF9282F8B0",
 -5672 => x"C0C0C0BF9282F8A4",
 -5671 => x"C0C0C0BF9282F8F9",
 -5670 => x"C0C0C0BF9282F8C0",
 -5669 => x"C0C0C0BF92828290",
 -5668 => x"C0C0C0BF92828280",
 -5667 => x"C0C0C0BF928282F8",
 -5666 => x"C0C0C0BF92828282",
 -5665 => x"C0C0C0BF92828292",
 -5664 => x"C0C0C0BF92828299",
 -5663 => x"C0C0C0BF928282B0",
 -5662 => x"C0C0C0BF928282A4",
 -5661 => x"C0C0C0BF928282F9",
 -5660 => x"C0C0C0BF928282C0",
 -5659 => x"C0C0C0BF92829290",
 -5658 => x"C0C0C0BF92829280",
 -5657 => x"C0C0C0BF928292F8",
 -5656 => x"C0C0C0BF92829282",
 -5655 => x"C0C0C0BF92829292",
 -5654 => x"C0C0C0BF92829299",
 -5653 => x"C0C0C0BF928292B0",
 -5652 => x"C0C0C0BF928292A4",
 -5651 => x"C0C0C0BF928292F9",
 -5650 => x"C0C0C0BF928292C0",
 -5649 => x"C0C0C0BF92829990",
 -5648 => x"C0C0C0BF92829980",
 -5647 => x"C0C0C0BF928299F8",
 -5646 => x"C0C0C0BF92829982",
 -5645 => x"C0C0C0BF92829992",
 -5644 => x"C0C0C0BF92829999",
 -5643 => x"C0C0C0BF928299B0",
 -5642 => x"C0C0C0BF928299A4",
 -5641 => x"C0C0C0BF928299F9",
 -5640 => x"C0C0C0BF928299C0",
 -5639 => x"C0C0C0BF9282B090",
 -5638 => x"C0C0C0BF9282B080",
 -5637 => x"C0C0C0BF9282B0F8",
 -5636 => x"C0C0C0BF9282B082",
 -5635 => x"C0C0C0BF9282B092",
 -5634 => x"C0C0C0BF9282B099",
 -5633 => x"C0C0C0BF9282B0B0",
 -5632 => x"C0C0C0BF9282B0A4",
 -5631 => x"C0C0C0BF9282B0F9",
 -5630 => x"C0C0C0BF9282B0C0",
 -5629 => x"C0C0C0BF9282A490",
 -5628 => x"C0C0C0BF9282A480",
 -5627 => x"C0C0C0BF9282A4F8",
 -5626 => x"C0C0C0BF9282A482",
 -5625 => x"C0C0C0BF9282A492",
 -5624 => x"C0C0C0BF9282A499",
 -5623 => x"C0C0C0BF9282A4B0",
 -5622 => x"C0C0C0BF9282A4A4",
 -5621 => x"C0C0C0BF9282A4F9",
 -5620 => x"C0C0C0BF9282A4C0",
 -5619 => x"C0C0C0BF9282F990",
 -5618 => x"C0C0C0BF9282F980",
 -5617 => x"C0C0C0BF9282F9F8",
 -5616 => x"C0C0C0BF9282F982",
 -5615 => x"C0C0C0BF9282F992",
 -5614 => x"C0C0C0BF9282F999",
 -5613 => x"C0C0C0BF9282F9B0",
 -5612 => x"C0C0C0BF9282F9A4",
 -5611 => x"C0C0C0BF9282F9F9",
 -5610 => x"C0C0C0BF9282F9C0",
 -5609 => x"C0C0C0BF9282C090",
 -5608 => x"C0C0C0BF9282C080",
 -5607 => x"C0C0C0BF9282C0F8",
 -5606 => x"C0C0C0BF9282C082",
 -5605 => x"C0C0C0BF9282C092",
 -5604 => x"C0C0C0BF9282C099",
 -5603 => x"C0C0C0BF9282C0B0",
 -5602 => x"C0C0C0BF9282C0A4",
 -5601 => x"C0C0C0BF9282C0F9",
 -5600 => x"C0C0C0BF9282C0C0",
 -5599 => x"C0C0C0BF92929090",
 -5598 => x"C0C0C0BF92929080",
 -5597 => x"C0C0C0BF929290F8",
 -5596 => x"C0C0C0BF92929082",
 -5595 => x"C0C0C0BF92929092",
 -5594 => x"C0C0C0BF92929099",
 -5593 => x"C0C0C0BF929290B0",
 -5592 => x"C0C0C0BF929290A4",
 -5591 => x"C0C0C0BF929290F9",
 -5590 => x"C0C0C0BF929290C0",
 -5589 => x"C0C0C0BF92928090",
 -5588 => x"C0C0C0BF92928080",
 -5587 => x"C0C0C0BF929280F8",
 -5586 => x"C0C0C0BF92928082",
 -5585 => x"C0C0C0BF92928092",
 -5584 => x"C0C0C0BF92928099",
 -5583 => x"C0C0C0BF929280B0",
 -5582 => x"C0C0C0BF929280A4",
 -5581 => x"C0C0C0BF929280F9",
 -5580 => x"C0C0C0BF929280C0",
 -5579 => x"C0C0C0BF9292F890",
 -5578 => x"C0C0C0BF9292F880",
 -5577 => x"C0C0C0BF9292F8F8",
 -5576 => x"C0C0C0BF9292F882",
 -5575 => x"C0C0C0BF9292F892",
 -5574 => x"C0C0C0BF9292F899",
 -5573 => x"C0C0C0BF9292F8B0",
 -5572 => x"C0C0C0BF9292F8A4",
 -5571 => x"C0C0C0BF9292F8F9",
 -5570 => x"C0C0C0BF9292F8C0",
 -5569 => x"C0C0C0BF92928290",
 -5568 => x"C0C0C0BF92928280",
 -5567 => x"C0C0C0BF929282F8",
 -5566 => x"C0C0C0BF92928282",
 -5565 => x"C0C0C0BF92928292",
 -5564 => x"C0C0C0BF92928299",
 -5563 => x"C0C0C0BF929282B0",
 -5562 => x"C0C0C0BF929282A4",
 -5561 => x"C0C0C0BF929282F9",
 -5560 => x"C0C0C0BF929282C0",
 -5559 => x"C0C0C0BF92929290",
 -5558 => x"C0C0C0BF92929280",
 -5557 => x"C0C0C0BF929292F8",
 -5556 => x"C0C0C0BF92929282",
 -5555 => x"C0C0C0BF92929292",
 -5554 => x"C0C0C0BF92929299",
 -5553 => x"C0C0C0BF929292B0",
 -5552 => x"C0C0C0BF929292A4",
 -5551 => x"C0C0C0BF929292F9",
 -5550 => x"C0C0C0BF929292C0",
 -5549 => x"C0C0C0BF92929990",
 -5548 => x"C0C0C0BF92929980",
 -5547 => x"C0C0C0BF929299F8",
 -5546 => x"C0C0C0BF92929982",
 -5545 => x"C0C0C0BF92929992",
 -5544 => x"C0C0C0BF92929999",
 -5543 => x"C0C0C0BF929299B0",
 -5542 => x"C0C0C0BF929299A4",
 -5541 => x"C0C0C0BF929299F9",
 -5540 => x"C0C0C0BF929299C0",
 -5539 => x"C0C0C0BF9292B090",
 -5538 => x"C0C0C0BF9292B080",
 -5537 => x"C0C0C0BF9292B0F8",
 -5536 => x"C0C0C0BF9292B082",
 -5535 => x"C0C0C0BF9292B092",
 -5534 => x"C0C0C0BF9292B099",
 -5533 => x"C0C0C0BF9292B0B0",
 -5532 => x"C0C0C0BF9292B0A4",
 -5531 => x"C0C0C0BF9292B0F9",
 -5530 => x"C0C0C0BF9292B0C0",
 -5529 => x"C0C0C0BF9292A490",
 -5528 => x"C0C0C0BF9292A480",
 -5527 => x"C0C0C0BF9292A4F8",
 -5526 => x"C0C0C0BF9292A482",
 -5525 => x"C0C0C0BF9292A492",
 -5524 => x"C0C0C0BF9292A499",
 -5523 => x"C0C0C0BF9292A4B0",
 -5522 => x"C0C0C0BF9292A4A4",
 -5521 => x"C0C0C0BF9292A4F9",
 -5520 => x"C0C0C0BF9292A4C0",
 -5519 => x"C0C0C0BF9292F990",
 -5518 => x"C0C0C0BF9292F980",
 -5517 => x"C0C0C0BF9292F9F8",
 -5516 => x"C0C0C0BF9292F982",
 -5515 => x"C0C0C0BF9292F992",
 -5514 => x"C0C0C0BF9292F999",
 -5513 => x"C0C0C0BF9292F9B0",
 -5512 => x"C0C0C0BF9292F9A4",
 -5511 => x"C0C0C0BF9292F9F9",
 -5510 => x"C0C0C0BF9292F9C0",
 -5509 => x"C0C0C0BF9292C090",
 -5508 => x"C0C0C0BF9292C080",
 -5507 => x"C0C0C0BF9292C0F8",
 -5506 => x"C0C0C0BF9292C082",
 -5505 => x"C0C0C0BF9292C092",
 -5504 => x"C0C0C0BF9292C099",
 -5503 => x"C0C0C0BF9292C0B0",
 -5502 => x"C0C0C0BF9292C0A4",
 -5501 => x"C0C0C0BF9292C0F9",
 -5500 => x"C0C0C0BF9292C0C0",
 -5499 => x"C0C0C0BF92999090",
 -5498 => x"C0C0C0BF92999080",
 -5497 => x"C0C0C0BF929990F8",
 -5496 => x"C0C0C0BF92999082",
 -5495 => x"C0C0C0BF92999092",
 -5494 => x"C0C0C0BF92999099",
 -5493 => x"C0C0C0BF929990B0",
 -5492 => x"C0C0C0BF929990A4",
 -5491 => x"C0C0C0BF929990F9",
 -5490 => x"C0C0C0BF929990C0",
 -5489 => x"C0C0C0BF92998090",
 -5488 => x"C0C0C0BF92998080",
 -5487 => x"C0C0C0BF929980F8",
 -5486 => x"C0C0C0BF92998082",
 -5485 => x"C0C0C0BF92998092",
 -5484 => x"C0C0C0BF92998099",
 -5483 => x"C0C0C0BF929980B0",
 -5482 => x"C0C0C0BF929980A4",
 -5481 => x"C0C0C0BF929980F9",
 -5480 => x"C0C0C0BF929980C0",
 -5479 => x"C0C0C0BF9299F890",
 -5478 => x"C0C0C0BF9299F880",
 -5477 => x"C0C0C0BF9299F8F8",
 -5476 => x"C0C0C0BF9299F882",
 -5475 => x"C0C0C0BF9299F892",
 -5474 => x"C0C0C0BF9299F899",
 -5473 => x"C0C0C0BF9299F8B0",
 -5472 => x"C0C0C0BF9299F8A4",
 -5471 => x"C0C0C0BF9299F8F9",
 -5470 => x"C0C0C0BF9299F8C0",
 -5469 => x"C0C0C0BF92998290",
 -5468 => x"C0C0C0BF92998280",
 -5467 => x"C0C0C0BF929982F8",
 -5466 => x"C0C0C0BF92998282",
 -5465 => x"C0C0C0BF92998292",
 -5464 => x"C0C0C0BF92998299",
 -5463 => x"C0C0C0BF929982B0",
 -5462 => x"C0C0C0BF929982A4",
 -5461 => x"C0C0C0BF929982F9",
 -5460 => x"C0C0C0BF929982C0",
 -5459 => x"C0C0C0BF92999290",
 -5458 => x"C0C0C0BF92999280",
 -5457 => x"C0C0C0BF929992F8",
 -5456 => x"C0C0C0BF92999282",
 -5455 => x"C0C0C0BF92999292",
 -5454 => x"C0C0C0BF92999299",
 -5453 => x"C0C0C0BF929992B0",
 -5452 => x"C0C0C0BF929992A4",
 -5451 => x"C0C0C0BF929992F9",
 -5450 => x"C0C0C0BF929992C0",
 -5449 => x"C0C0C0BF92999990",
 -5448 => x"C0C0C0BF92999980",
 -5447 => x"C0C0C0BF929999F8",
 -5446 => x"C0C0C0BF92999982",
 -5445 => x"C0C0C0BF92999992",
 -5444 => x"C0C0C0BF92999999",
 -5443 => x"C0C0C0BF929999B0",
 -5442 => x"C0C0C0BF929999A4",
 -5441 => x"C0C0C0BF929999F9",
 -5440 => x"C0C0C0BF929999C0",
 -5439 => x"C0C0C0BF9299B090",
 -5438 => x"C0C0C0BF9299B080",
 -5437 => x"C0C0C0BF9299B0F8",
 -5436 => x"C0C0C0BF9299B082",
 -5435 => x"C0C0C0BF9299B092",
 -5434 => x"C0C0C0BF9299B099",
 -5433 => x"C0C0C0BF9299B0B0",
 -5432 => x"C0C0C0BF9299B0A4",
 -5431 => x"C0C0C0BF9299B0F9",
 -5430 => x"C0C0C0BF9299B0C0",
 -5429 => x"C0C0C0BF9299A490",
 -5428 => x"C0C0C0BF9299A480",
 -5427 => x"C0C0C0BF9299A4F8",
 -5426 => x"C0C0C0BF9299A482",
 -5425 => x"C0C0C0BF9299A492",
 -5424 => x"C0C0C0BF9299A499",
 -5423 => x"C0C0C0BF9299A4B0",
 -5422 => x"C0C0C0BF9299A4A4",
 -5421 => x"C0C0C0BF9299A4F9",
 -5420 => x"C0C0C0BF9299A4C0",
 -5419 => x"C0C0C0BF9299F990",
 -5418 => x"C0C0C0BF9299F980",
 -5417 => x"C0C0C0BF9299F9F8",
 -5416 => x"C0C0C0BF9299F982",
 -5415 => x"C0C0C0BF9299F992",
 -5414 => x"C0C0C0BF9299F999",
 -5413 => x"C0C0C0BF9299F9B0",
 -5412 => x"C0C0C0BF9299F9A4",
 -5411 => x"C0C0C0BF9299F9F9",
 -5410 => x"C0C0C0BF9299F9C0",
 -5409 => x"C0C0C0BF9299C090",
 -5408 => x"C0C0C0BF9299C080",
 -5407 => x"C0C0C0BF9299C0F8",
 -5406 => x"C0C0C0BF9299C082",
 -5405 => x"C0C0C0BF9299C092",
 -5404 => x"C0C0C0BF9299C099",
 -5403 => x"C0C0C0BF9299C0B0",
 -5402 => x"C0C0C0BF9299C0A4",
 -5401 => x"C0C0C0BF9299C0F9",
 -5400 => x"C0C0C0BF9299C0C0",
 -5399 => x"C0C0C0BF92B09090",
 -5398 => x"C0C0C0BF92B09080",
 -5397 => x"C0C0C0BF92B090F8",
 -5396 => x"C0C0C0BF92B09082",
 -5395 => x"C0C0C0BF92B09092",
 -5394 => x"C0C0C0BF92B09099",
 -5393 => x"C0C0C0BF92B090B0",
 -5392 => x"C0C0C0BF92B090A4",
 -5391 => x"C0C0C0BF92B090F9",
 -5390 => x"C0C0C0BF92B090C0",
 -5389 => x"C0C0C0BF92B08090",
 -5388 => x"C0C0C0BF92B08080",
 -5387 => x"C0C0C0BF92B080F8",
 -5386 => x"C0C0C0BF92B08082",
 -5385 => x"C0C0C0BF92B08092",
 -5384 => x"C0C0C0BF92B08099",
 -5383 => x"C0C0C0BF92B080B0",
 -5382 => x"C0C0C0BF92B080A4",
 -5381 => x"C0C0C0BF92B080F9",
 -5380 => x"C0C0C0BF92B080C0",
 -5379 => x"C0C0C0BF92B0F890",
 -5378 => x"C0C0C0BF92B0F880",
 -5377 => x"C0C0C0BF92B0F8F8",
 -5376 => x"C0C0C0BF92B0F882",
 -5375 => x"C0C0C0BF92B0F892",
 -5374 => x"C0C0C0BF92B0F899",
 -5373 => x"C0C0C0BF92B0F8B0",
 -5372 => x"C0C0C0BF92B0F8A4",
 -5371 => x"C0C0C0BF92B0F8F9",
 -5370 => x"C0C0C0BF92B0F8C0",
 -5369 => x"C0C0C0BF92B08290",
 -5368 => x"C0C0C0BF92B08280",
 -5367 => x"C0C0C0BF92B082F8",
 -5366 => x"C0C0C0BF92B08282",
 -5365 => x"C0C0C0BF92B08292",
 -5364 => x"C0C0C0BF92B08299",
 -5363 => x"C0C0C0BF92B082B0",
 -5362 => x"C0C0C0BF92B082A4",
 -5361 => x"C0C0C0BF92B082F9",
 -5360 => x"C0C0C0BF92B082C0",
 -5359 => x"C0C0C0BF92B09290",
 -5358 => x"C0C0C0BF92B09280",
 -5357 => x"C0C0C0BF92B092F8",
 -5356 => x"C0C0C0BF92B09282",
 -5355 => x"C0C0C0BF92B09292",
 -5354 => x"C0C0C0BF92B09299",
 -5353 => x"C0C0C0BF92B092B0",
 -5352 => x"C0C0C0BF92B092A4",
 -5351 => x"C0C0C0BF92B092F9",
 -5350 => x"C0C0C0BF92B092C0",
 -5349 => x"C0C0C0BF92B09990",
 -5348 => x"C0C0C0BF92B09980",
 -5347 => x"C0C0C0BF92B099F8",
 -5346 => x"C0C0C0BF92B09982",
 -5345 => x"C0C0C0BF92B09992",
 -5344 => x"C0C0C0BF92B09999",
 -5343 => x"C0C0C0BF92B099B0",
 -5342 => x"C0C0C0BF92B099A4",
 -5341 => x"C0C0C0BF92B099F9",
 -5340 => x"C0C0C0BF92B099C0",
 -5339 => x"C0C0C0BF92B0B090",
 -5338 => x"C0C0C0BF92B0B080",
 -5337 => x"C0C0C0BF92B0B0F8",
 -5336 => x"C0C0C0BF92B0B082",
 -5335 => x"C0C0C0BF92B0B092",
 -5334 => x"C0C0C0BF92B0B099",
 -5333 => x"C0C0C0BF92B0B0B0",
 -5332 => x"C0C0C0BF92B0B0A4",
 -5331 => x"C0C0C0BF92B0B0F9",
 -5330 => x"C0C0C0BF92B0B0C0",
 -5329 => x"C0C0C0BF92B0A490",
 -5328 => x"C0C0C0BF92B0A480",
 -5327 => x"C0C0C0BF92B0A4F8",
 -5326 => x"C0C0C0BF92B0A482",
 -5325 => x"C0C0C0BF92B0A492",
 -5324 => x"C0C0C0BF92B0A499",
 -5323 => x"C0C0C0BF92B0A4B0",
 -5322 => x"C0C0C0BF92B0A4A4",
 -5321 => x"C0C0C0BF92B0A4F9",
 -5320 => x"C0C0C0BF92B0A4C0",
 -5319 => x"C0C0C0BF92B0F990",
 -5318 => x"C0C0C0BF92B0F980",
 -5317 => x"C0C0C0BF92B0F9F8",
 -5316 => x"C0C0C0BF92B0F982",
 -5315 => x"C0C0C0BF92B0F992",
 -5314 => x"C0C0C0BF92B0F999",
 -5313 => x"C0C0C0BF92B0F9B0",
 -5312 => x"C0C0C0BF92B0F9A4",
 -5311 => x"C0C0C0BF92B0F9F9",
 -5310 => x"C0C0C0BF92B0F9C0",
 -5309 => x"C0C0C0BF92B0C090",
 -5308 => x"C0C0C0BF92B0C080",
 -5307 => x"C0C0C0BF92B0C0F8",
 -5306 => x"C0C0C0BF92B0C082",
 -5305 => x"C0C0C0BF92B0C092",
 -5304 => x"C0C0C0BF92B0C099",
 -5303 => x"C0C0C0BF92B0C0B0",
 -5302 => x"C0C0C0BF92B0C0A4",
 -5301 => x"C0C0C0BF92B0C0F9",
 -5300 => x"C0C0C0BF92B0C0C0",
 -5299 => x"C0C0C0BF92A49090",
 -5298 => x"C0C0C0BF92A49080",
 -5297 => x"C0C0C0BF92A490F8",
 -5296 => x"C0C0C0BF92A49082",
 -5295 => x"C0C0C0BF92A49092",
 -5294 => x"C0C0C0BF92A49099",
 -5293 => x"C0C0C0BF92A490B0",
 -5292 => x"C0C0C0BF92A490A4",
 -5291 => x"C0C0C0BF92A490F9",
 -5290 => x"C0C0C0BF92A490C0",
 -5289 => x"C0C0C0BF92A48090",
 -5288 => x"C0C0C0BF92A48080",
 -5287 => x"C0C0C0BF92A480F8",
 -5286 => x"C0C0C0BF92A48082",
 -5285 => x"C0C0C0BF92A48092",
 -5284 => x"C0C0C0BF92A48099",
 -5283 => x"C0C0C0BF92A480B0",
 -5282 => x"C0C0C0BF92A480A4",
 -5281 => x"C0C0C0BF92A480F9",
 -5280 => x"C0C0C0BF92A480C0",
 -5279 => x"C0C0C0BF92A4F890",
 -5278 => x"C0C0C0BF92A4F880",
 -5277 => x"C0C0C0BF92A4F8F8",
 -5276 => x"C0C0C0BF92A4F882",
 -5275 => x"C0C0C0BF92A4F892",
 -5274 => x"C0C0C0BF92A4F899",
 -5273 => x"C0C0C0BF92A4F8B0",
 -5272 => x"C0C0C0BF92A4F8A4",
 -5271 => x"C0C0C0BF92A4F8F9",
 -5270 => x"C0C0C0BF92A4F8C0",
 -5269 => x"C0C0C0BF92A48290",
 -5268 => x"C0C0C0BF92A48280",
 -5267 => x"C0C0C0BF92A482F8",
 -5266 => x"C0C0C0BF92A48282",
 -5265 => x"C0C0C0BF92A48292",
 -5264 => x"C0C0C0BF92A48299",
 -5263 => x"C0C0C0BF92A482B0",
 -5262 => x"C0C0C0BF92A482A4",
 -5261 => x"C0C0C0BF92A482F9",
 -5260 => x"C0C0C0BF92A482C0",
 -5259 => x"C0C0C0BF92A49290",
 -5258 => x"C0C0C0BF92A49280",
 -5257 => x"C0C0C0BF92A492F8",
 -5256 => x"C0C0C0BF92A49282",
 -5255 => x"C0C0C0BF92A49292",
 -5254 => x"C0C0C0BF92A49299",
 -5253 => x"C0C0C0BF92A492B0",
 -5252 => x"C0C0C0BF92A492A4",
 -5251 => x"C0C0C0BF92A492F9",
 -5250 => x"C0C0C0BF92A492C0",
 -5249 => x"C0C0C0BF92A49990",
 -5248 => x"C0C0C0BF92A49980",
 -5247 => x"C0C0C0BF92A499F8",
 -5246 => x"C0C0C0BF92A49982",
 -5245 => x"C0C0C0BF92A49992",
 -5244 => x"C0C0C0BF92A49999",
 -5243 => x"C0C0C0BF92A499B0",
 -5242 => x"C0C0C0BF92A499A4",
 -5241 => x"C0C0C0BF92A499F9",
 -5240 => x"C0C0C0BF92A499C0",
 -5239 => x"C0C0C0BF92A4B090",
 -5238 => x"C0C0C0BF92A4B080",
 -5237 => x"C0C0C0BF92A4B0F8",
 -5236 => x"C0C0C0BF92A4B082",
 -5235 => x"C0C0C0BF92A4B092",
 -5234 => x"C0C0C0BF92A4B099",
 -5233 => x"C0C0C0BF92A4B0B0",
 -5232 => x"C0C0C0BF92A4B0A4",
 -5231 => x"C0C0C0BF92A4B0F9",
 -5230 => x"C0C0C0BF92A4B0C0",
 -5229 => x"C0C0C0BF92A4A490",
 -5228 => x"C0C0C0BF92A4A480",
 -5227 => x"C0C0C0BF92A4A4F8",
 -5226 => x"C0C0C0BF92A4A482",
 -5225 => x"C0C0C0BF92A4A492",
 -5224 => x"C0C0C0BF92A4A499",
 -5223 => x"C0C0C0BF92A4A4B0",
 -5222 => x"C0C0C0BF92A4A4A4",
 -5221 => x"C0C0C0BF92A4A4F9",
 -5220 => x"C0C0C0BF92A4A4C0",
 -5219 => x"C0C0C0BF92A4F990",
 -5218 => x"C0C0C0BF92A4F980",
 -5217 => x"C0C0C0BF92A4F9F8",
 -5216 => x"C0C0C0BF92A4F982",
 -5215 => x"C0C0C0BF92A4F992",
 -5214 => x"C0C0C0BF92A4F999",
 -5213 => x"C0C0C0BF92A4F9B0",
 -5212 => x"C0C0C0BF92A4F9A4",
 -5211 => x"C0C0C0BF92A4F9F9",
 -5210 => x"C0C0C0BF92A4F9C0",
 -5209 => x"C0C0C0BF92A4C090",
 -5208 => x"C0C0C0BF92A4C080",
 -5207 => x"C0C0C0BF92A4C0F8",
 -5206 => x"C0C0C0BF92A4C082",
 -5205 => x"C0C0C0BF92A4C092",
 -5204 => x"C0C0C0BF92A4C099",
 -5203 => x"C0C0C0BF92A4C0B0",
 -5202 => x"C0C0C0BF92A4C0A4",
 -5201 => x"C0C0C0BF92A4C0F9",
 -5200 => x"C0C0C0BF92A4C0C0",
 -5199 => x"C0C0C0BF92F99090",
 -5198 => x"C0C0C0BF92F99080",
 -5197 => x"C0C0C0BF92F990F8",
 -5196 => x"C0C0C0BF92F99082",
 -5195 => x"C0C0C0BF92F99092",
 -5194 => x"C0C0C0BF92F99099",
 -5193 => x"C0C0C0BF92F990B0",
 -5192 => x"C0C0C0BF92F990A4",
 -5191 => x"C0C0C0BF92F990F9",
 -5190 => x"C0C0C0BF92F990C0",
 -5189 => x"C0C0C0BF92F98090",
 -5188 => x"C0C0C0BF92F98080",
 -5187 => x"C0C0C0BF92F980F8",
 -5186 => x"C0C0C0BF92F98082",
 -5185 => x"C0C0C0BF92F98092",
 -5184 => x"C0C0C0BF92F98099",
 -5183 => x"C0C0C0BF92F980B0",
 -5182 => x"C0C0C0BF92F980A4",
 -5181 => x"C0C0C0BF92F980F9",
 -5180 => x"C0C0C0BF92F980C0",
 -5179 => x"C0C0C0BF92F9F890",
 -5178 => x"C0C0C0BF92F9F880",
 -5177 => x"C0C0C0BF92F9F8F8",
 -5176 => x"C0C0C0BF92F9F882",
 -5175 => x"C0C0C0BF92F9F892",
 -5174 => x"C0C0C0BF92F9F899",
 -5173 => x"C0C0C0BF92F9F8B0",
 -5172 => x"C0C0C0BF92F9F8A4",
 -5171 => x"C0C0C0BF92F9F8F9",
 -5170 => x"C0C0C0BF92F9F8C0",
 -5169 => x"C0C0C0BF92F98290",
 -5168 => x"C0C0C0BF92F98280",
 -5167 => x"C0C0C0BF92F982F8",
 -5166 => x"C0C0C0BF92F98282",
 -5165 => x"C0C0C0BF92F98292",
 -5164 => x"C0C0C0BF92F98299",
 -5163 => x"C0C0C0BF92F982B0",
 -5162 => x"C0C0C0BF92F982A4",
 -5161 => x"C0C0C0BF92F982F9",
 -5160 => x"C0C0C0BF92F982C0",
 -5159 => x"C0C0C0BF92F99290",
 -5158 => x"C0C0C0BF92F99280",
 -5157 => x"C0C0C0BF92F992F8",
 -5156 => x"C0C0C0BF92F99282",
 -5155 => x"C0C0C0BF92F99292",
 -5154 => x"C0C0C0BF92F99299",
 -5153 => x"C0C0C0BF92F992B0",
 -5152 => x"C0C0C0BF92F992A4",
 -5151 => x"C0C0C0BF92F992F9",
 -5150 => x"C0C0C0BF92F992C0",
 -5149 => x"C0C0C0BF92F99990",
 -5148 => x"C0C0C0BF92F99980",
 -5147 => x"C0C0C0BF92F999F8",
 -5146 => x"C0C0C0BF92F99982",
 -5145 => x"C0C0C0BF92F99992",
 -5144 => x"C0C0C0BF92F99999",
 -5143 => x"C0C0C0BF92F999B0",
 -5142 => x"C0C0C0BF92F999A4",
 -5141 => x"C0C0C0BF92F999F9",
 -5140 => x"C0C0C0BF92F999C0",
 -5139 => x"C0C0C0BF92F9B090",
 -5138 => x"C0C0C0BF92F9B080",
 -5137 => x"C0C0C0BF92F9B0F8",
 -5136 => x"C0C0C0BF92F9B082",
 -5135 => x"C0C0C0BF92F9B092",
 -5134 => x"C0C0C0BF92F9B099",
 -5133 => x"C0C0C0BF92F9B0B0",
 -5132 => x"C0C0C0BF92F9B0A4",
 -5131 => x"C0C0C0BF92F9B0F9",
 -5130 => x"C0C0C0BF92F9B0C0",
 -5129 => x"C0C0C0BF92F9A490",
 -5128 => x"C0C0C0BF92F9A480",
 -5127 => x"C0C0C0BF92F9A4F8",
 -5126 => x"C0C0C0BF92F9A482",
 -5125 => x"C0C0C0BF92F9A492",
 -5124 => x"C0C0C0BF92F9A499",
 -5123 => x"C0C0C0BF92F9A4B0",
 -5122 => x"C0C0C0BF92F9A4A4",
 -5121 => x"C0C0C0BF92F9A4F9",
 -5120 => x"C0C0C0BF92F9A4C0",
 -5119 => x"C0C0C0BF92F9F990",
 -5118 => x"C0C0C0BF92F9F980",
 -5117 => x"C0C0C0BF92F9F9F8",
 -5116 => x"C0C0C0BF92F9F982",
 -5115 => x"C0C0C0BF92F9F992",
 -5114 => x"C0C0C0BF92F9F999",
 -5113 => x"C0C0C0BF92F9F9B0",
 -5112 => x"C0C0C0BF92F9F9A4",
 -5111 => x"C0C0C0BF92F9F9F9",
 -5110 => x"C0C0C0BF92F9F9C0",
 -5109 => x"C0C0C0BF92F9C090",
 -5108 => x"C0C0C0BF92F9C080",
 -5107 => x"C0C0C0BF92F9C0F8",
 -5106 => x"C0C0C0BF92F9C082",
 -5105 => x"C0C0C0BF92F9C092",
 -5104 => x"C0C0C0BF92F9C099",
 -5103 => x"C0C0C0BF92F9C0B0",
 -5102 => x"C0C0C0BF92F9C0A4",
 -5101 => x"C0C0C0BF92F9C0F9",
 -5100 => x"C0C0C0BF92F9C0C0",
 -5099 => x"C0C0C0BF92C09090",
 -5098 => x"C0C0C0BF92C09080",
 -5097 => x"C0C0C0BF92C090F8",
 -5096 => x"C0C0C0BF92C09082",
 -5095 => x"C0C0C0BF92C09092",
 -5094 => x"C0C0C0BF92C09099",
 -5093 => x"C0C0C0BF92C090B0",
 -5092 => x"C0C0C0BF92C090A4",
 -5091 => x"C0C0C0BF92C090F9",
 -5090 => x"C0C0C0BF92C090C0",
 -5089 => x"C0C0C0BF92C08090",
 -5088 => x"C0C0C0BF92C08080",
 -5087 => x"C0C0C0BF92C080F8",
 -5086 => x"C0C0C0BF92C08082",
 -5085 => x"C0C0C0BF92C08092",
 -5084 => x"C0C0C0BF92C08099",
 -5083 => x"C0C0C0BF92C080B0",
 -5082 => x"C0C0C0BF92C080A4",
 -5081 => x"C0C0C0BF92C080F9",
 -5080 => x"C0C0C0BF92C080C0",
 -5079 => x"C0C0C0BF92C0F890",
 -5078 => x"C0C0C0BF92C0F880",
 -5077 => x"C0C0C0BF92C0F8F8",
 -5076 => x"C0C0C0BF92C0F882",
 -5075 => x"C0C0C0BF92C0F892",
 -5074 => x"C0C0C0BF92C0F899",
 -5073 => x"C0C0C0BF92C0F8B0",
 -5072 => x"C0C0C0BF92C0F8A4",
 -5071 => x"C0C0C0BF92C0F8F9",
 -5070 => x"C0C0C0BF92C0F8C0",
 -5069 => x"C0C0C0BF92C08290",
 -5068 => x"C0C0C0BF92C08280",
 -5067 => x"C0C0C0BF92C082F8",
 -5066 => x"C0C0C0BF92C08282",
 -5065 => x"C0C0C0BF92C08292",
 -5064 => x"C0C0C0BF92C08299",
 -5063 => x"C0C0C0BF92C082B0",
 -5062 => x"C0C0C0BF92C082A4",
 -5061 => x"C0C0C0BF92C082F9",
 -5060 => x"C0C0C0BF92C082C0",
 -5059 => x"C0C0C0BF92C09290",
 -5058 => x"C0C0C0BF92C09280",
 -5057 => x"C0C0C0BF92C092F8",
 -5056 => x"C0C0C0BF92C09282",
 -5055 => x"C0C0C0BF92C09292",
 -5054 => x"C0C0C0BF92C09299",
 -5053 => x"C0C0C0BF92C092B0",
 -5052 => x"C0C0C0BF92C092A4",
 -5051 => x"C0C0C0BF92C092F9",
 -5050 => x"C0C0C0BF92C092C0",
 -5049 => x"C0C0C0BF92C09990",
 -5048 => x"C0C0C0BF92C09980",
 -5047 => x"C0C0C0BF92C099F8",
 -5046 => x"C0C0C0BF92C09982",
 -5045 => x"C0C0C0BF92C09992",
 -5044 => x"C0C0C0BF92C09999",
 -5043 => x"C0C0C0BF92C099B0",
 -5042 => x"C0C0C0BF92C099A4",
 -5041 => x"C0C0C0BF92C099F9",
 -5040 => x"C0C0C0BF92C099C0",
 -5039 => x"C0C0C0BF92C0B090",
 -5038 => x"C0C0C0BF92C0B080",
 -5037 => x"C0C0C0BF92C0B0F8",
 -5036 => x"C0C0C0BF92C0B082",
 -5035 => x"C0C0C0BF92C0B092",
 -5034 => x"C0C0C0BF92C0B099",
 -5033 => x"C0C0C0BF92C0B0B0",
 -5032 => x"C0C0C0BF92C0B0A4",
 -5031 => x"C0C0C0BF92C0B0F9",
 -5030 => x"C0C0C0BF92C0B0C0",
 -5029 => x"C0C0C0BF92C0A490",
 -5028 => x"C0C0C0BF92C0A480",
 -5027 => x"C0C0C0BF92C0A4F8",
 -5026 => x"C0C0C0BF92C0A482",
 -5025 => x"C0C0C0BF92C0A492",
 -5024 => x"C0C0C0BF92C0A499",
 -5023 => x"C0C0C0BF92C0A4B0",
 -5022 => x"C0C0C0BF92C0A4A4",
 -5021 => x"C0C0C0BF92C0A4F9",
 -5020 => x"C0C0C0BF92C0A4C0",
 -5019 => x"C0C0C0BF92C0F990",
 -5018 => x"C0C0C0BF92C0F980",
 -5017 => x"C0C0C0BF92C0F9F8",
 -5016 => x"C0C0C0BF92C0F982",
 -5015 => x"C0C0C0BF92C0F992",
 -5014 => x"C0C0C0BF92C0F999",
 -5013 => x"C0C0C0BF92C0F9B0",
 -5012 => x"C0C0C0BF92C0F9A4",
 -5011 => x"C0C0C0BF92C0F9F9",
 -5010 => x"C0C0C0BF92C0F9C0",
 -5009 => x"C0C0C0BF92C0C090",
 -5008 => x"C0C0C0BF92C0C080",
 -5007 => x"C0C0C0BF92C0C0F8",
 -5006 => x"C0C0C0BF92C0C082",
 -5005 => x"C0C0C0BF92C0C092",
 -5004 => x"C0C0C0BF92C0C099",
 -5003 => x"C0C0C0BF92C0C0B0",
 -5002 => x"C0C0C0BF92C0C0A4",
 -5001 => x"C0C0C0BF92C0C0F9",
 -5000 => x"C0C0C0BF92C0C0C0",
 -4999 => x"C0C0C0BF99909090",
 -4998 => x"C0C0C0BF99909080",
 -4997 => x"C0C0C0BF999090F8",
 -4996 => x"C0C0C0BF99909082",
 -4995 => x"C0C0C0BF99909092",
 -4994 => x"C0C0C0BF99909099",
 -4993 => x"C0C0C0BF999090B0",
 -4992 => x"C0C0C0BF999090A4",
 -4991 => x"C0C0C0BF999090F9",
 -4990 => x"C0C0C0BF999090C0",
 -4989 => x"C0C0C0BF99908090",
 -4988 => x"C0C0C0BF99908080",
 -4987 => x"C0C0C0BF999080F8",
 -4986 => x"C0C0C0BF99908082",
 -4985 => x"C0C0C0BF99908092",
 -4984 => x"C0C0C0BF99908099",
 -4983 => x"C0C0C0BF999080B0",
 -4982 => x"C0C0C0BF999080A4",
 -4981 => x"C0C0C0BF999080F9",
 -4980 => x"C0C0C0BF999080C0",
 -4979 => x"C0C0C0BF9990F890",
 -4978 => x"C0C0C0BF9990F880",
 -4977 => x"C0C0C0BF9990F8F8",
 -4976 => x"C0C0C0BF9990F882",
 -4975 => x"C0C0C0BF9990F892",
 -4974 => x"C0C0C0BF9990F899",
 -4973 => x"C0C0C0BF9990F8B0",
 -4972 => x"C0C0C0BF9990F8A4",
 -4971 => x"C0C0C0BF9990F8F9",
 -4970 => x"C0C0C0BF9990F8C0",
 -4969 => x"C0C0C0BF99908290",
 -4968 => x"C0C0C0BF99908280",
 -4967 => x"C0C0C0BF999082F8",
 -4966 => x"C0C0C0BF99908282",
 -4965 => x"C0C0C0BF99908292",
 -4964 => x"C0C0C0BF99908299",
 -4963 => x"C0C0C0BF999082B0",
 -4962 => x"C0C0C0BF999082A4",
 -4961 => x"C0C0C0BF999082F9",
 -4960 => x"C0C0C0BF999082C0",
 -4959 => x"C0C0C0BF99909290",
 -4958 => x"C0C0C0BF99909280",
 -4957 => x"C0C0C0BF999092F8",
 -4956 => x"C0C0C0BF99909282",
 -4955 => x"C0C0C0BF99909292",
 -4954 => x"C0C0C0BF99909299",
 -4953 => x"C0C0C0BF999092B0",
 -4952 => x"C0C0C0BF999092A4",
 -4951 => x"C0C0C0BF999092F9",
 -4950 => x"C0C0C0BF999092C0",
 -4949 => x"C0C0C0BF99909990",
 -4948 => x"C0C0C0BF99909980",
 -4947 => x"C0C0C0BF999099F8",
 -4946 => x"C0C0C0BF99909982",
 -4945 => x"C0C0C0BF99909992",
 -4944 => x"C0C0C0BF99909999",
 -4943 => x"C0C0C0BF999099B0",
 -4942 => x"C0C0C0BF999099A4",
 -4941 => x"C0C0C0BF999099F9",
 -4940 => x"C0C0C0BF999099C0",
 -4939 => x"C0C0C0BF9990B090",
 -4938 => x"C0C0C0BF9990B080",
 -4937 => x"C0C0C0BF9990B0F8",
 -4936 => x"C0C0C0BF9990B082",
 -4935 => x"C0C0C0BF9990B092",
 -4934 => x"C0C0C0BF9990B099",
 -4933 => x"C0C0C0BF9990B0B0",
 -4932 => x"C0C0C0BF9990B0A4",
 -4931 => x"C0C0C0BF9990B0F9",
 -4930 => x"C0C0C0BF9990B0C0",
 -4929 => x"C0C0C0BF9990A490",
 -4928 => x"C0C0C0BF9990A480",
 -4927 => x"C0C0C0BF9990A4F8",
 -4926 => x"C0C0C0BF9990A482",
 -4925 => x"C0C0C0BF9990A492",
 -4924 => x"C0C0C0BF9990A499",
 -4923 => x"C0C0C0BF9990A4B0",
 -4922 => x"C0C0C0BF9990A4A4",
 -4921 => x"C0C0C0BF9990A4F9",
 -4920 => x"C0C0C0BF9990A4C0",
 -4919 => x"C0C0C0BF9990F990",
 -4918 => x"C0C0C0BF9990F980",
 -4917 => x"C0C0C0BF9990F9F8",
 -4916 => x"C0C0C0BF9990F982",
 -4915 => x"C0C0C0BF9990F992",
 -4914 => x"C0C0C0BF9990F999",
 -4913 => x"C0C0C0BF9990F9B0",
 -4912 => x"C0C0C0BF9990F9A4",
 -4911 => x"C0C0C0BF9990F9F9",
 -4910 => x"C0C0C0BF9990F9C0",
 -4909 => x"C0C0C0BF9990C090",
 -4908 => x"C0C0C0BF9990C080",
 -4907 => x"C0C0C0BF9990C0F8",
 -4906 => x"C0C0C0BF9990C082",
 -4905 => x"C0C0C0BF9990C092",
 -4904 => x"C0C0C0BF9990C099",
 -4903 => x"C0C0C0BF9990C0B0",
 -4902 => x"C0C0C0BF9990C0A4",
 -4901 => x"C0C0C0BF9990C0F9",
 -4900 => x"C0C0C0BF9990C0C0",
 -4899 => x"C0C0C0BF99809090",
 -4898 => x"C0C0C0BF99809080",
 -4897 => x"C0C0C0BF998090F8",
 -4896 => x"C0C0C0BF99809082",
 -4895 => x"C0C0C0BF99809092",
 -4894 => x"C0C0C0BF99809099",
 -4893 => x"C0C0C0BF998090B0",
 -4892 => x"C0C0C0BF998090A4",
 -4891 => x"C0C0C0BF998090F9",
 -4890 => x"C0C0C0BF998090C0",
 -4889 => x"C0C0C0BF99808090",
 -4888 => x"C0C0C0BF99808080",
 -4887 => x"C0C0C0BF998080F8",
 -4886 => x"C0C0C0BF99808082",
 -4885 => x"C0C0C0BF99808092",
 -4884 => x"C0C0C0BF99808099",
 -4883 => x"C0C0C0BF998080B0",
 -4882 => x"C0C0C0BF998080A4",
 -4881 => x"C0C0C0BF998080F9",
 -4880 => x"C0C0C0BF998080C0",
 -4879 => x"C0C0C0BF9980F890",
 -4878 => x"C0C0C0BF9980F880",
 -4877 => x"C0C0C0BF9980F8F8",
 -4876 => x"C0C0C0BF9980F882",
 -4875 => x"C0C0C0BF9980F892",
 -4874 => x"C0C0C0BF9980F899",
 -4873 => x"C0C0C0BF9980F8B0",
 -4872 => x"C0C0C0BF9980F8A4",
 -4871 => x"C0C0C0BF9980F8F9",
 -4870 => x"C0C0C0BF9980F8C0",
 -4869 => x"C0C0C0BF99808290",
 -4868 => x"C0C0C0BF99808280",
 -4867 => x"C0C0C0BF998082F8",
 -4866 => x"C0C0C0BF99808282",
 -4865 => x"C0C0C0BF99808292",
 -4864 => x"C0C0C0BF99808299",
 -4863 => x"C0C0C0BF998082B0",
 -4862 => x"C0C0C0BF998082A4",
 -4861 => x"C0C0C0BF998082F9",
 -4860 => x"C0C0C0BF998082C0",
 -4859 => x"C0C0C0BF99809290",
 -4858 => x"C0C0C0BF99809280",
 -4857 => x"C0C0C0BF998092F8",
 -4856 => x"C0C0C0BF99809282",
 -4855 => x"C0C0C0BF99809292",
 -4854 => x"C0C0C0BF99809299",
 -4853 => x"C0C0C0BF998092B0",
 -4852 => x"C0C0C0BF998092A4",
 -4851 => x"C0C0C0BF998092F9",
 -4850 => x"C0C0C0BF998092C0",
 -4849 => x"C0C0C0BF99809990",
 -4848 => x"C0C0C0BF99809980",
 -4847 => x"C0C0C0BF998099F8",
 -4846 => x"C0C0C0BF99809982",
 -4845 => x"C0C0C0BF99809992",
 -4844 => x"C0C0C0BF99809999",
 -4843 => x"C0C0C0BF998099B0",
 -4842 => x"C0C0C0BF998099A4",
 -4841 => x"C0C0C0BF998099F9",
 -4840 => x"C0C0C0BF998099C0",
 -4839 => x"C0C0C0BF9980B090",
 -4838 => x"C0C0C0BF9980B080",
 -4837 => x"C0C0C0BF9980B0F8",
 -4836 => x"C0C0C0BF9980B082",
 -4835 => x"C0C0C0BF9980B092",
 -4834 => x"C0C0C0BF9980B099",
 -4833 => x"C0C0C0BF9980B0B0",
 -4832 => x"C0C0C0BF9980B0A4",
 -4831 => x"C0C0C0BF9980B0F9",
 -4830 => x"C0C0C0BF9980B0C0",
 -4829 => x"C0C0C0BF9980A490",
 -4828 => x"C0C0C0BF9980A480",
 -4827 => x"C0C0C0BF9980A4F8",
 -4826 => x"C0C0C0BF9980A482",
 -4825 => x"C0C0C0BF9980A492",
 -4824 => x"C0C0C0BF9980A499",
 -4823 => x"C0C0C0BF9980A4B0",
 -4822 => x"C0C0C0BF9980A4A4",
 -4821 => x"C0C0C0BF9980A4F9",
 -4820 => x"C0C0C0BF9980A4C0",
 -4819 => x"C0C0C0BF9980F990",
 -4818 => x"C0C0C0BF9980F980",
 -4817 => x"C0C0C0BF9980F9F8",
 -4816 => x"C0C0C0BF9980F982",
 -4815 => x"C0C0C0BF9980F992",
 -4814 => x"C0C0C0BF9980F999",
 -4813 => x"C0C0C0BF9980F9B0",
 -4812 => x"C0C0C0BF9980F9A4",
 -4811 => x"C0C0C0BF9980F9F9",
 -4810 => x"C0C0C0BF9980F9C0",
 -4809 => x"C0C0C0BF9980C090",
 -4808 => x"C0C0C0BF9980C080",
 -4807 => x"C0C0C0BF9980C0F8",
 -4806 => x"C0C0C0BF9980C082",
 -4805 => x"C0C0C0BF9980C092",
 -4804 => x"C0C0C0BF9980C099",
 -4803 => x"C0C0C0BF9980C0B0",
 -4802 => x"C0C0C0BF9980C0A4",
 -4801 => x"C0C0C0BF9980C0F9",
 -4800 => x"C0C0C0BF9980C0C0",
 -4799 => x"C0C0C0BF99F89090",
 -4798 => x"C0C0C0BF99F89080",
 -4797 => x"C0C0C0BF99F890F8",
 -4796 => x"C0C0C0BF99F89082",
 -4795 => x"C0C0C0BF99F89092",
 -4794 => x"C0C0C0BF99F89099",
 -4793 => x"C0C0C0BF99F890B0",
 -4792 => x"C0C0C0BF99F890A4",
 -4791 => x"C0C0C0BF99F890F9",
 -4790 => x"C0C0C0BF99F890C0",
 -4789 => x"C0C0C0BF99F88090",
 -4788 => x"C0C0C0BF99F88080",
 -4787 => x"C0C0C0BF99F880F8",
 -4786 => x"C0C0C0BF99F88082",
 -4785 => x"C0C0C0BF99F88092",
 -4784 => x"C0C0C0BF99F88099",
 -4783 => x"C0C0C0BF99F880B0",
 -4782 => x"C0C0C0BF99F880A4",
 -4781 => x"C0C0C0BF99F880F9",
 -4780 => x"C0C0C0BF99F880C0",
 -4779 => x"C0C0C0BF99F8F890",
 -4778 => x"C0C0C0BF99F8F880",
 -4777 => x"C0C0C0BF99F8F8F8",
 -4776 => x"C0C0C0BF99F8F882",
 -4775 => x"C0C0C0BF99F8F892",
 -4774 => x"C0C0C0BF99F8F899",
 -4773 => x"C0C0C0BF99F8F8B0",
 -4772 => x"C0C0C0BF99F8F8A4",
 -4771 => x"C0C0C0BF99F8F8F9",
 -4770 => x"C0C0C0BF99F8F8C0",
 -4769 => x"C0C0C0BF99F88290",
 -4768 => x"C0C0C0BF99F88280",
 -4767 => x"C0C0C0BF99F882F8",
 -4766 => x"C0C0C0BF99F88282",
 -4765 => x"C0C0C0BF99F88292",
 -4764 => x"C0C0C0BF99F88299",
 -4763 => x"C0C0C0BF99F882B0",
 -4762 => x"C0C0C0BF99F882A4",
 -4761 => x"C0C0C0BF99F882F9",
 -4760 => x"C0C0C0BF99F882C0",
 -4759 => x"C0C0C0BF99F89290",
 -4758 => x"C0C0C0BF99F89280",
 -4757 => x"C0C0C0BF99F892F8",
 -4756 => x"C0C0C0BF99F89282",
 -4755 => x"C0C0C0BF99F89292",
 -4754 => x"C0C0C0BF99F89299",
 -4753 => x"C0C0C0BF99F892B0",
 -4752 => x"C0C0C0BF99F892A4",
 -4751 => x"C0C0C0BF99F892F9",
 -4750 => x"C0C0C0BF99F892C0",
 -4749 => x"C0C0C0BF99F89990",
 -4748 => x"C0C0C0BF99F89980",
 -4747 => x"C0C0C0BF99F899F8",
 -4746 => x"C0C0C0BF99F89982",
 -4745 => x"C0C0C0BF99F89992",
 -4744 => x"C0C0C0BF99F89999",
 -4743 => x"C0C0C0BF99F899B0",
 -4742 => x"C0C0C0BF99F899A4",
 -4741 => x"C0C0C0BF99F899F9",
 -4740 => x"C0C0C0BF99F899C0",
 -4739 => x"C0C0C0BF99F8B090",
 -4738 => x"C0C0C0BF99F8B080",
 -4737 => x"C0C0C0BF99F8B0F8",
 -4736 => x"C0C0C0BF99F8B082",
 -4735 => x"C0C0C0BF99F8B092",
 -4734 => x"C0C0C0BF99F8B099",
 -4733 => x"C0C0C0BF99F8B0B0",
 -4732 => x"C0C0C0BF99F8B0A4",
 -4731 => x"C0C0C0BF99F8B0F9",
 -4730 => x"C0C0C0BF99F8B0C0",
 -4729 => x"C0C0C0BF99F8A490",
 -4728 => x"C0C0C0BF99F8A480",
 -4727 => x"C0C0C0BF99F8A4F8",
 -4726 => x"C0C0C0BF99F8A482",
 -4725 => x"C0C0C0BF99F8A492",
 -4724 => x"C0C0C0BF99F8A499",
 -4723 => x"C0C0C0BF99F8A4B0",
 -4722 => x"C0C0C0BF99F8A4A4",
 -4721 => x"C0C0C0BF99F8A4F9",
 -4720 => x"C0C0C0BF99F8A4C0",
 -4719 => x"C0C0C0BF99F8F990",
 -4718 => x"C0C0C0BF99F8F980",
 -4717 => x"C0C0C0BF99F8F9F8",
 -4716 => x"C0C0C0BF99F8F982",
 -4715 => x"C0C0C0BF99F8F992",
 -4714 => x"C0C0C0BF99F8F999",
 -4713 => x"C0C0C0BF99F8F9B0",
 -4712 => x"C0C0C0BF99F8F9A4",
 -4711 => x"C0C0C0BF99F8F9F9",
 -4710 => x"C0C0C0BF99F8F9C0",
 -4709 => x"C0C0C0BF99F8C090",
 -4708 => x"C0C0C0BF99F8C080",
 -4707 => x"C0C0C0BF99F8C0F8",
 -4706 => x"C0C0C0BF99F8C082",
 -4705 => x"C0C0C0BF99F8C092",
 -4704 => x"C0C0C0BF99F8C099",
 -4703 => x"C0C0C0BF99F8C0B0",
 -4702 => x"C0C0C0BF99F8C0A4",
 -4701 => x"C0C0C0BF99F8C0F9",
 -4700 => x"C0C0C0BF99F8C0C0",
 -4699 => x"C0C0C0BF99829090",
 -4698 => x"C0C0C0BF99829080",
 -4697 => x"C0C0C0BF998290F8",
 -4696 => x"C0C0C0BF99829082",
 -4695 => x"C0C0C0BF99829092",
 -4694 => x"C0C0C0BF99829099",
 -4693 => x"C0C0C0BF998290B0",
 -4692 => x"C0C0C0BF998290A4",
 -4691 => x"C0C0C0BF998290F9",
 -4690 => x"C0C0C0BF998290C0",
 -4689 => x"C0C0C0BF99828090",
 -4688 => x"C0C0C0BF99828080",
 -4687 => x"C0C0C0BF998280F8",
 -4686 => x"C0C0C0BF99828082",
 -4685 => x"C0C0C0BF99828092",
 -4684 => x"C0C0C0BF99828099",
 -4683 => x"C0C0C0BF998280B0",
 -4682 => x"C0C0C0BF998280A4",
 -4681 => x"C0C0C0BF998280F9",
 -4680 => x"C0C0C0BF998280C0",
 -4679 => x"C0C0C0BF9982F890",
 -4678 => x"C0C0C0BF9982F880",
 -4677 => x"C0C0C0BF9982F8F8",
 -4676 => x"C0C0C0BF9982F882",
 -4675 => x"C0C0C0BF9982F892",
 -4674 => x"C0C0C0BF9982F899",
 -4673 => x"C0C0C0BF9982F8B0",
 -4672 => x"C0C0C0BF9982F8A4",
 -4671 => x"C0C0C0BF9982F8F9",
 -4670 => x"C0C0C0BF9982F8C0",
 -4669 => x"C0C0C0BF99828290",
 -4668 => x"C0C0C0BF99828280",
 -4667 => x"C0C0C0BF998282F8",
 -4666 => x"C0C0C0BF99828282",
 -4665 => x"C0C0C0BF99828292",
 -4664 => x"C0C0C0BF99828299",
 -4663 => x"C0C0C0BF998282B0",
 -4662 => x"C0C0C0BF998282A4",
 -4661 => x"C0C0C0BF998282F9",
 -4660 => x"C0C0C0BF998282C0",
 -4659 => x"C0C0C0BF99829290",
 -4658 => x"C0C0C0BF99829280",
 -4657 => x"C0C0C0BF998292F8",
 -4656 => x"C0C0C0BF99829282",
 -4655 => x"C0C0C0BF99829292",
 -4654 => x"C0C0C0BF99829299",
 -4653 => x"C0C0C0BF998292B0",
 -4652 => x"C0C0C0BF998292A4",
 -4651 => x"C0C0C0BF998292F9",
 -4650 => x"C0C0C0BF998292C0",
 -4649 => x"C0C0C0BF99829990",
 -4648 => x"C0C0C0BF99829980",
 -4647 => x"C0C0C0BF998299F8",
 -4646 => x"C0C0C0BF99829982",
 -4645 => x"C0C0C0BF99829992",
 -4644 => x"C0C0C0BF99829999",
 -4643 => x"C0C0C0BF998299B0",
 -4642 => x"C0C0C0BF998299A4",
 -4641 => x"C0C0C0BF998299F9",
 -4640 => x"C0C0C0BF998299C0",
 -4639 => x"C0C0C0BF9982B090",
 -4638 => x"C0C0C0BF9982B080",
 -4637 => x"C0C0C0BF9982B0F8",
 -4636 => x"C0C0C0BF9982B082",
 -4635 => x"C0C0C0BF9982B092",
 -4634 => x"C0C0C0BF9982B099",
 -4633 => x"C0C0C0BF9982B0B0",
 -4632 => x"C0C0C0BF9982B0A4",
 -4631 => x"C0C0C0BF9982B0F9",
 -4630 => x"C0C0C0BF9982B0C0",
 -4629 => x"C0C0C0BF9982A490",
 -4628 => x"C0C0C0BF9982A480",
 -4627 => x"C0C0C0BF9982A4F8",
 -4626 => x"C0C0C0BF9982A482",
 -4625 => x"C0C0C0BF9982A492",
 -4624 => x"C0C0C0BF9982A499",
 -4623 => x"C0C0C0BF9982A4B0",
 -4622 => x"C0C0C0BF9982A4A4",
 -4621 => x"C0C0C0BF9982A4F9",
 -4620 => x"C0C0C0BF9982A4C0",
 -4619 => x"C0C0C0BF9982F990",
 -4618 => x"C0C0C0BF9982F980",
 -4617 => x"C0C0C0BF9982F9F8",
 -4616 => x"C0C0C0BF9982F982",
 -4615 => x"C0C0C0BF9982F992",
 -4614 => x"C0C0C0BF9982F999",
 -4613 => x"C0C0C0BF9982F9B0",
 -4612 => x"C0C0C0BF9982F9A4",
 -4611 => x"C0C0C0BF9982F9F9",
 -4610 => x"C0C0C0BF9982F9C0",
 -4609 => x"C0C0C0BF9982C090",
 -4608 => x"C0C0C0BF9982C080",
 -4607 => x"C0C0C0BF9982C0F8",
 -4606 => x"C0C0C0BF9982C082",
 -4605 => x"C0C0C0BF9982C092",
 -4604 => x"C0C0C0BF9982C099",
 -4603 => x"C0C0C0BF9982C0B0",
 -4602 => x"C0C0C0BF9982C0A4",
 -4601 => x"C0C0C0BF9982C0F9",
 -4600 => x"C0C0C0BF9982C0C0",
 -4599 => x"C0C0C0BF99929090",
 -4598 => x"C0C0C0BF99929080",
 -4597 => x"C0C0C0BF999290F8",
 -4596 => x"C0C0C0BF99929082",
 -4595 => x"C0C0C0BF99929092",
 -4594 => x"C0C0C0BF99929099",
 -4593 => x"C0C0C0BF999290B0",
 -4592 => x"C0C0C0BF999290A4",
 -4591 => x"C0C0C0BF999290F9",
 -4590 => x"C0C0C0BF999290C0",
 -4589 => x"C0C0C0BF99928090",
 -4588 => x"C0C0C0BF99928080",
 -4587 => x"C0C0C0BF999280F8",
 -4586 => x"C0C0C0BF99928082",
 -4585 => x"C0C0C0BF99928092",
 -4584 => x"C0C0C0BF99928099",
 -4583 => x"C0C0C0BF999280B0",
 -4582 => x"C0C0C0BF999280A4",
 -4581 => x"C0C0C0BF999280F9",
 -4580 => x"C0C0C0BF999280C0",
 -4579 => x"C0C0C0BF9992F890",
 -4578 => x"C0C0C0BF9992F880",
 -4577 => x"C0C0C0BF9992F8F8",
 -4576 => x"C0C0C0BF9992F882",
 -4575 => x"C0C0C0BF9992F892",
 -4574 => x"C0C0C0BF9992F899",
 -4573 => x"C0C0C0BF9992F8B0",
 -4572 => x"C0C0C0BF9992F8A4",
 -4571 => x"C0C0C0BF9992F8F9",
 -4570 => x"C0C0C0BF9992F8C0",
 -4569 => x"C0C0C0BF99928290",
 -4568 => x"C0C0C0BF99928280",
 -4567 => x"C0C0C0BF999282F8",
 -4566 => x"C0C0C0BF99928282",
 -4565 => x"C0C0C0BF99928292",
 -4564 => x"C0C0C0BF99928299",
 -4563 => x"C0C0C0BF999282B0",
 -4562 => x"C0C0C0BF999282A4",
 -4561 => x"C0C0C0BF999282F9",
 -4560 => x"C0C0C0BF999282C0",
 -4559 => x"C0C0C0BF99929290",
 -4558 => x"C0C0C0BF99929280",
 -4557 => x"C0C0C0BF999292F8",
 -4556 => x"C0C0C0BF99929282",
 -4555 => x"C0C0C0BF99929292",
 -4554 => x"C0C0C0BF99929299",
 -4553 => x"C0C0C0BF999292B0",
 -4552 => x"C0C0C0BF999292A4",
 -4551 => x"C0C0C0BF999292F9",
 -4550 => x"C0C0C0BF999292C0",
 -4549 => x"C0C0C0BF99929990",
 -4548 => x"C0C0C0BF99929980",
 -4547 => x"C0C0C0BF999299F8",
 -4546 => x"C0C0C0BF99929982",
 -4545 => x"C0C0C0BF99929992",
 -4544 => x"C0C0C0BF99929999",
 -4543 => x"C0C0C0BF999299B0",
 -4542 => x"C0C0C0BF999299A4",
 -4541 => x"C0C0C0BF999299F9",
 -4540 => x"C0C0C0BF999299C0",
 -4539 => x"C0C0C0BF9992B090",
 -4538 => x"C0C0C0BF9992B080",
 -4537 => x"C0C0C0BF9992B0F8",
 -4536 => x"C0C0C0BF9992B082",
 -4535 => x"C0C0C0BF9992B092",
 -4534 => x"C0C0C0BF9992B099",
 -4533 => x"C0C0C0BF9992B0B0",
 -4532 => x"C0C0C0BF9992B0A4",
 -4531 => x"C0C0C0BF9992B0F9",
 -4530 => x"C0C0C0BF9992B0C0",
 -4529 => x"C0C0C0BF9992A490",
 -4528 => x"C0C0C0BF9992A480",
 -4527 => x"C0C0C0BF9992A4F8",
 -4526 => x"C0C0C0BF9992A482",
 -4525 => x"C0C0C0BF9992A492",
 -4524 => x"C0C0C0BF9992A499",
 -4523 => x"C0C0C0BF9992A4B0",
 -4522 => x"C0C0C0BF9992A4A4",
 -4521 => x"C0C0C0BF9992A4F9",
 -4520 => x"C0C0C0BF9992A4C0",
 -4519 => x"C0C0C0BF9992F990",
 -4518 => x"C0C0C0BF9992F980",
 -4517 => x"C0C0C0BF9992F9F8",
 -4516 => x"C0C0C0BF9992F982",
 -4515 => x"C0C0C0BF9992F992",
 -4514 => x"C0C0C0BF9992F999",
 -4513 => x"C0C0C0BF9992F9B0",
 -4512 => x"C0C0C0BF9992F9A4",
 -4511 => x"C0C0C0BF9992F9F9",
 -4510 => x"C0C0C0BF9992F9C0",
 -4509 => x"C0C0C0BF9992C090",
 -4508 => x"C0C0C0BF9992C080",
 -4507 => x"C0C0C0BF9992C0F8",
 -4506 => x"C0C0C0BF9992C082",
 -4505 => x"C0C0C0BF9992C092",
 -4504 => x"C0C0C0BF9992C099",
 -4503 => x"C0C0C0BF9992C0B0",
 -4502 => x"C0C0C0BF9992C0A4",
 -4501 => x"C0C0C0BF9992C0F9",
 -4500 => x"C0C0C0BF9992C0C0",
 -4499 => x"C0C0C0BF99999090",
 -4498 => x"C0C0C0BF99999080",
 -4497 => x"C0C0C0BF999990F8",
 -4496 => x"C0C0C0BF99999082",
 -4495 => x"C0C0C0BF99999092",
 -4494 => x"C0C0C0BF99999099",
 -4493 => x"C0C0C0BF999990B0",
 -4492 => x"C0C0C0BF999990A4",
 -4491 => x"C0C0C0BF999990F9",
 -4490 => x"C0C0C0BF999990C0",
 -4489 => x"C0C0C0BF99998090",
 -4488 => x"C0C0C0BF99998080",
 -4487 => x"C0C0C0BF999980F8",
 -4486 => x"C0C0C0BF99998082",
 -4485 => x"C0C0C0BF99998092",
 -4484 => x"C0C0C0BF99998099",
 -4483 => x"C0C0C0BF999980B0",
 -4482 => x"C0C0C0BF999980A4",
 -4481 => x"C0C0C0BF999980F9",
 -4480 => x"C0C0C0BF999980C0",
 -4479 => x"C0C0C0BF9999F890",
 -4478 => x"C0C0C0BF9999F880",
 -4477 => x"C0C0C0BF9999F8F8",
 -4476 => x"C0C0C0BF9999F882",
 -4475 => x"C0C0C0BF9999F892",
 -4474 => x"C0C0C0BF9999F899",
 -4473 => x"C0C0C0BF9999F8B0",
 -4472 => x"C0C0C0BF9999F8A4",
 -4471 => x"C0C0C0BF9999F8F9",
 -4470 => x"C0C0C0BF9999F8C0",
 -4469 => x"C0C0C0BF99998290",
 -4468 => x"C0C0C0BF99998280",
 -4467 => x"C0C0C0BF999982F8",
 -4466 => x"C0C0C0BF99998282",
 -4465 => x"C0C0C0BF99998292",
 -4464 => x"C0C0C0BF99998299",
 -4463 => x"C0C0C0BF999982B0",
 -4462 => x"C0C0C0BF999982A4",
 -4461 => x"C0C0C0BF999982F9",
 -4460 => x"C0C0C0BF999982C0",
 -4459 => x"C0C0C0BF99999290",
 -4458 => x"C0C0C0BF99999280",
 -4457 => x"C0C0C0BF999992F8",
 -4456 => x"C0C0C0BF99999282",
 -4455 => x"C0C0C0BF99999292",
 -4454 => x"C0C0C0BF99999299",
 -4453 => x"C0C0C0BF999992B0",
 -4452 => x"C0C0C0BF999992A4",
 -4451 => x"C0C0C0BF999992F9",
 -4450 => x"C0C0C0BF999992C0",
 -4449 => x"C0C0C0BF99999990",
 -4448 => x"C0C0C0BF99999980",
 -4447 => x"C0C0C0BF999999F8",
 -4446 => x"C0C0C0BF99999982",
 -4445 => x"C0C0C0BF99999992",
 -4444 => x"C0C0C0BF99999999",
 -4443 => x"C0C0C0BF999999B0",
 -4442 => x"C0C0C0BF999999A4",
 -4441 => x"C0C0C0BF999999F9",
 -4440 => x"C0C0C0BF999999C0",
 -4439 => x"C0C0C0BF9999B090",
 -4438 => x"C0C0C0BF9999B080",
 -4437 => x"C0C0C0BF9999B0F8",
 -4436 => x"C0C0C0BF9999B082",
 -4435 => x"C0C0C0BF9999B092",
 -4434 => x"C0C0C0BF9999B099",
 -4433 => x"C0C0C0BF9999B0B0",
 -4432 => x"C0C0C0BF9999B0A4",
 -4431 => x"C0C0C0BF9999B0F9",
 -4430 => x"C0C0C0BF9999B0C0",
 -4429 => x"C0C0C0BF9999A490",
 -4428 => x"C0C0C0BF9999A480",
 -4427 => x"C0C0C0BF9999A4F8",
 -4426 => x"C0C0C0BF9999A482",
 -4425 => x"C0C0C0BF9999A492",
 -4424 => x"C0C0C0BF9999A499",
 -4423 => x"C0C0C0BF9999A4B0",
 -4422 => x"C0C0C0BF9999A4A4",
 -4421 => x"C0C0C0BF9999A4F9",
 -4420 => x"C0C0C0BF9999A4C0",
 -4419 => x"C0C0C0BF9999F990",
 -4418 => x"C0C0C0BF9999F980",
 -4417 => x"C0C0C0BF9999F9F8",
 -4416 => x"C0C0C0BF9999F982",
 -4415 => x"C0C0C0BF9999F992",
 -4414 => x"C0C0C0BF9999F999",
 -4413 => x"C0C0C0BF9999F9B0",
 -4412 => x"C0C0C0BF9999F9A4",
 -4411 => x"C0C0C0BF9999F9F9",
 -4410 => x"C0C0C0BF9999F9C0",
 -4409 => x"C0C0C0BF9999C090",
 -4408 => x"C0C0C0BF9999C080",
 -4407 => x"C0C0C0BF9999C0F8",
 -4406 => x"C0C0C0BF9999C082",
 -4405 => x"C0C0C0BF9999C092",
 -4404 => x"C0C0C0BF9999C099",
 -4403 => x"C0C0C0BF9999C0B0",
 -4402 => x"C0C0C0BF9999C0A4",
 -4401 => x"C0C0C0BF9999C0F9",
 -4400 => x"C0C0C0BF9999C0C0",
 -4399 => x"C0C0C0BF99B09090",
 -4398 => x"C0C0C0BF99B09080",
 -4397 => x"C0C0C0BF99B090F8",
 -4396 => x"C0C0C0BF99B09082",
 -4395 => x"C0C0C0BF99B09092",
 -4394 => x"C0C0C0BF99B09099",
 -4393 => x"C0C0C0BF99B090B0",
 -4392 => x"C0C0C0BF99B090A4",
 -4391 => x"C0C0C0BF99B090F9",
 -4390 => x"C0C0C0BF99B090C0",
 -4389 => x"C0C0C0BF99B08090",
 -4388 => x"C0C0C0BF99B08080",
 -4387 => x"C0C0C0BF99B080F8",
 -4386 => x"C0C0C0BF99B08082",
 -4385 => x"C0C0C0BF99B08092",
 -4384 => x"C0C0C0BF99B08099",
 -4383 => x"C0C0C0BF99B080B0",
 -4382 => x"C0C0C0BF99B080A4",
 -4381 => x"C0C0C0BF99B080F9",
 -4380 => x"C0C0C0BF99B080C0",
 -4379 => x"C0C0C0BF99B0F890",
 -4378 => x"C0C0C0BF99B0F880",
 -4377 => x"C0C0C0BF99B0F8F8",
 -4376 => x"C0C0C0BF99B0F882",
 -4375 => x"C0C0C0BF99B0F892",
 -4374 => x"C0C0C0BF99B0F899",
 -4373 => x"C0C0C0BF99B0F8B0",
 -4372 => x"C0C0C0BF99B0F8A4",
 -4371 => x"C0C0C0BF99B0F8F9",
 -4370 => x"C0C0C0BF99B0F8C0",
 -4369 => x"C0C0C0BF99B08290",
 -4368 => x"C0C0C0BF99B08280",
 -4367 => x"C0C0C0BF99B082F8",
 -4366 => x"C0C0C0BF99B08282",
 -4365 => x"C0C0C0BF99B08292",
 -4364 => x"C0C0C0BF99B08299",
 -4363 => x"C0C0C0BF99B082B0",
 -4362 => x"C0C0C0BF99B082A4",
 -4361 => x"C0C0C0BF99B082F9",
 -4360 => x"C0C0C0BF99B082C0",
 -4359 => x"C0C0C0BF99B09290",
 -4358 => x"C0C0C0BF99B09280",
 -4357 => x"C0C0C0BF99B092F8",
 -4356 => x"C0C0C0BF99B09282",
 -4355 => x"C0C0C0BF99B09292",
 -4354 => x"C0C0C0BF99B09299",
 -4353 => x"C0C0C0BF99B092B0",
 -4352 => x"C0C0C0BF99B092A4",
 -4351 => x"C0C0C0BF99B092F9",
 -4350 => x"C0C0C0BF99B092C0",
 -4349 => x"C0C0C0BF99B09990",
 -4348 => x"C0C0C0BF99B09980",
 -4347 => x"C0C0C0BF99B099F8",
 -4346 => x"C0C0C0BF99B09982",
 -4345 => x"C0C0C0BF99B09992",
 -4344 => x"C0C0C0BF99B09999",
 -4343 => x"C0C0C0BF99B099B0",
 -4342 => x"C0C0C0BF99B099A4",
 -4341 => x"C0C0C0BF99B099F9",
 -4340 => x"C0C0C0BF99B099C0",
 -4339 => x"C0C0C0BF99B0B090",
 -4338 => x"C0C0C0BF99B0B080",
 -4337 => x"C0C0C0BF99B0B0F8",
 -4336 => x"C0C0C0BF99B0B082",
 -4335 => x"C0C0C0BF99B0B092",
 -4334 => x"C0C0C0BF99B0B099",
 -4333 => x"C0C0C0BF99B0B0B0",
 -4332 => x"C0C0C0BF99B0B0A4",
 -4331 => x"C0C0C0BF99B0B0F9",
 -4330 => x"C0C0C0BF99B0B0C0",
 -4329 => x"C0C0C0BF99B0A490",
 -4328 => x"C0C0C0BF99B0A480",
 -4327 => x"C0C0C0BF99B0A4F8",
 -4326 => x"C0C0C0BF99B0A482",
 -4325 => x"C0C0C0BF99B0A492",
 -4324 => x"C0C0C0BF99B0A499",
 -4323 => x"C0C0C0BF99B0A4B0",
 -4322 => x"C0C0C0BF99B0A4A4",
 -4321 => x"C0C0C0BF99B0A4F9",
 -4320 => x"C0C0C0BF99B0A4C0",
 -4319 => x"C0C0C0BF99B0F990",
 -4318 => x"C0C0C0BF99B0F980",
 -4317 => x"C0C0C0BF99B0F9F8",
 -4316 => x"C0C0C0BF99B0F982",
 -4315 => x"C0C0C0BF99B0F992",
 -4314 => x"C0C0C0BF99B0F999",
 -4313 => x"C0C0C0BF99B0F9B0",
 -4312 => x"C0C0C0BF99B0F9A4",
 -4311 => x"C0C0C0BF99B0F9F9",
 -4310 => x"C0C0C0BF99B0F9C0",
 -4309 => x"C0C0C0BF99B0C090",
 -4308 => x"C0C0C0BF99B0C080",
 -4307 => x"C0C0C0BF99B0C0F8",
 -4306 => x"C0C0C0BF99B0C082",
 -4305 => x"C0C0C0BF99B0C092",
 -4304 => x"C0C0C0BF99B0C099",
 -4303 => x"C0C0C0BF99B0C0B0",
 -4302 => x"C0C0C0BF99B0C0A4",
 -4301 => x"C0C0C0BF99B0C0F9",
 -4300 => x"C0C0C0BF99B0C0C0",
 -4299 => x"C0C0C0BF99A49090",
 -4298 => x"C0C0C0BF99A49080",
 -4297 => x"C0C0C0BF99A490F8",
 -4296 => x"C0C0C0BF99A49082",
 -4295 => x"C0C0C0BF99A49092",
 -4294 => x"C0C0C0BF99A49099",
 -4293 => x"C0C0C0BF99A490B0",
 -4292 => x"C0C0C0BF99A490A4",
 -4291 => x"C0C0C0BF99A490F9",
 -4290 => x"C0C0C0BF99A490C0",
 -4289 => x"C0C0C0BF99A48090",
 -4288 => x"C0C0C0BF99A48080",
 -4287 => x"C0C0C0BF99A480F8",
 -4286 => x"C0C0C0BF99A48082",
 -4285 => x"C0C0C0BF99A48092",
 -4284 => x"C0C0C0BF99A48099",
 -4283 => x"C0C0C0BF99A480B0",
 -4282 => x"C0C0C0BF99A480A4",
 -4281 => x"C0C0C0BF99A480F9",
 -4280 => x"C0C0C0BF99A480C0",
 -4279 => x"C0C0C0BF99A4F890",
 -4278 => x"C0C0C0BF99A4F880",
 -4277 => x"C0C0C0BF99A4F8F8",
 -4276 => x"C0C0C0BF99A4F882",
 -4275 => x"C0C0C0BF99A4F892",
 -4274 => x"C0C0C0BF99A4F899",
 -4273 => x"C0C0C0BF99A4F8B0",
 -4272 => x"C0C0C0BF99A4F8A4",
 -4271 => x"C0C0C0BF99A4F8F9",
 -4270 => x"C0C0C0BF99A4F8C0",
 -4269 => x"C0C0C0BF99A48290",
 -4268 => x"C0C0C0BF99A48280",
 -4267 => x"C0C0C0BF99A482F8",
 -4266 => x"C0C0C0BF99A48282",
 -4265 => x"C0C0C0BF99A48292",
 -4264 => x"C0C0C0BF99A48299",
 -4263 => x"C0C0C0BF99A482B0",
 -4262 => x"C0C0C0BF99A482A4",
 -4261 => x"C0C0C0BF99A482F9",
 -4260 => x"C0C0C0BF99A482C0",
 -4259 => x"C0C0C0BF99A49290",
 -4258 => x"C0C0C0BF99A49280",
 -4257 => x"C0C0C0BF99A492F8",
 -4256 => x"C0C0C0BF99A49282",
 -4255 => x"C0C0C0BF99A49292",
 -4254 => x"C0C0C0BF99A49299",
 -4253 => x"C0C0C0BF99A492B0",
 -4252 => x"C0C0C0BF99A492A4",
 -4251 => x"C0C0C0BF99A492F9",
 -4250 => x"C0C0C0BF99A492C0",
 -4249 => x"C0C0C0BF99A49990",
 -4248 => x"C0C0C0BF99A49980",
 -4247 => x"C0C0C0BF99A499F8",
 -4246 => x"C0C0C0BF99A49982",
 -4245 => x"C0C0C0BF99A49992",
 -4244 => x"C0C0C0BF99A49999",
 -4243 => x"C0C0C0BF99A499B0",
 -4242 => x"C0C0C0BF99A499A4",
 -4241 => x"C0C0C0BF99A499F9",
 -4240 => x"C0C0C0BF99A499C0",
 -4239 => x"C0C0C0BF99A4B090",
 -4238 => x"C0C0C0BF99A4B080",
 -4237 => x"C0C0C0BF99A4B0F8",
 -4236 => x"C0C0C0BF99A4B082",
 -4235 => x"C0C0C0BF99A4B092",
 -4234 => x"C0C0C0BF99A4B099",
 -4233 => x"C0C0C0BF99A4B0B0",
 -4232 => x"C0C0C0BF99A4B0A4",
 -4231 => x"C0C0C0BF99A4B0F9",
 -4230 => x"C0C0C0BF99A4B0C0",
 -4229 => x"C0C0C0BF99A4A490",
 -4228 => x"C0C0C0BF99A4A480",
 -4227 => x"C0C0C0BF99A4A4F8",
 -4226 => x"C0C0C0BF99A4A482",
 -4225 => x"C0C0C0BF99A4A492",
 -4224 => x"C0C0C0BF99A4A499",
 -4223 => x"C0C0C0BF99A4A4B0",
 -4222 => x"C0C0C0BF99A4A4A4",
 -4221 => x"C0C0C0BF99A4A4F9",
 -4220 => x"C0C0C0BF99A4A4C0",
 -4219 => x"C0C0C0BF99A4F990",
 -4218 => x"C0C0C0BF99A4F980",
 -4217 => x"C0C0C0BF99A4F9F8",
 -4216 => x"C0C0C0BF99A4F982",
 -4215 => x"C0C0C0BF99A4F992",
 -4214 => x"C0C0C0BF99A4F999",
 -4213 => x"C0C0C0BF99A4F9B0",
 -4212 => x"C0C0C0BF99A4F9A4",
 -4211 => x"C0C0C0BF99A4F9F9",
 -4210 => x"C0C0C0BF99A4F9C0",
 -4209 => x"C0C0C0BF99A4C090",
 -4208 => x"C0C0C0BF99A4C080",
 -4207 => x"C0C0C0BF99A4C0F8",
 -4206 => x"C0C0C0BF99A4C082",
 -4205 => x"C0C0C0BF99A4C092",
 -4204 => x"C0C0C0BF99A4C099",
 -4203 => x"C0C0C0BF99A4C0B0",
 -4202 => x"C0C0C0BF99A4C0A4",
 -4201 => x"C0C0C0BF99A4C0F9",
 -4200 => x"C0C0C0BF99A4C0C0",
 -4199 => x"C0C0C0BF99F99090",
 -4198 => x"C0C0C0BF99F99080",
 -4197 => x"C0C0C0BF99F990F8",
 -4196 => x"C0C0C0BF99F99082",
 -4195 => x"C0C0C0BF99F99092",
 -4194 => x"C0C0C0BF99F99099",
 -4193 => x"C0C0C0BF99F990B0",
 -4192 => x"C0C0C0BF99F990A4",
 -4191 => x"C0C0C0BF99F990F9",
 -4190 => x"C0C0C0BF99F990C0",
 -4189 => x"C0C0C0BF99F98090",
 -4188 => x"C0C0C0BF99F98080",
 -4187 => x"C0C0C0BF99F980F8",
 -4186 => x"C0C0C0BF99F98082",
 -4185 => x"C0C0C0BF99F98092",
 -4184 => x"C0C0C0BF99F98099",
 -4183 => x"C0C0C0BF99F980B0",
 -4182 => x"C0C0C0BF99F980A4",
 -4181 => x"C0C0C0BF99F980F9",
 -4180 => x"C0C0C0BF99F980C0",
 -4179 => x"C0C0C0BF99F9F890",
 -4178 => x"C0C0C0BF99F9F880",
 -4177 => x"C0C0C0BF99F9F8F8",
 -4176 => x"C0C0C0BF99F9F882",
 -4175 => x"C0C0C0BF99F9F892",
 -4174 => x"C0C0C0BF99F9F899",
 -4173 => x"C0C0C0BF99F9F8B0",
 -4172 => x"C0C0C0BF99F9F8A4",
 -4171 => x"C0C0C0BF99F9F8F9",
 -4170 => x"C0C0C0BF99F9F8C0",
 -4169 => x"C0C0C0BF99F98290",
 -4168 => x"C0C0C0BF99F98280",
 -4167 => x"C0C0C0BF99F982F8",
 -4166 => x"C0C0C0BF99F98282",
 -4165 => x"C0C0C0BF99F98292",
 -4164 => x"C0C0C0BF99F98299",
 -4163 => x"C0C0C0BF99F982B0",
 -4162 => x"C0C0C0BF99F982A4",
 -4161 => x"C0C0C0BF99F982F9",
 -4160 => x"C0C0C0BF99F982C0",
 -4159 => x"C0C0C0BF99F99290",
 -4158 => x"C0C0C0BF99F99280",
 -4157 => x"C0C0C0BF99F992F8",
 -4156 => x"C0C0C0BF99F99282",
 -4155 => x"C0C0C0BF99F99292",
 -4154 => x"C0C0C0BF99F99299",
 -4153 => x"C0C0C0BF99F992B0",
 -4152 => x"C0C0C0BF99F992A4",
 -4151 => x"C0C0C0BF99F992F9",
 -4150 => x"C0C0C0BF99F992C0",
 -4149 => x"C0C0C0BF99F99990",
 -4148 => x"C0C0C0BF99F99980",
 -4147 => x"C0C0C0BF99F999F8",
 -4146 => x"C0C0C0BF99F99982",
 -4145 => x"C0C0C0BF99F99992",
 -4144 => x"C0C0C0BF99F99999",
 -4143 => x"C0C0C0BF99F999B0",
 -4142 => x"C0C0C0BF99F999A4",
 -4141 => x"C0C0C0BF99F999F9",
 -4140 => x"C0C0C0BF99F999C0",
 -4139 => x"C0C0C0BF99F9B090",
 -4138 => x"C0C0C0BF99F9B080",
 -4137 => x"C0C0C0BF99F9B0F8",
 -4136 => x"C0C0C0BF99F9B082",
 -4135 => x"C0C0C0BF99F9B092",
 -4134 => x"C0C0C0BF99F9B099",
 -4133 => x"C0C0C0BF99F9B0B0",
 -4132 => x"C0C0C0BF99F9B0A4",
 -4131 => x"C0C0C0BF99F9B0F9",
 -4130 => x"C0C0C0BF99F9B0C0",
 -4129 => x"C0C0C0BF99F9A490",
 -4128 => x"C0C0C0BF99F9A480",
 -4127 => x"C0C0C0BF99F9A4F8",
 -4126 => x"C0C0C0BF99F9A482",
 -4125 => x"C0C0C0BF99F9A492",
 -4124 => x"C0C0C0BF99F9A499",
 -4123 => x"C0C0C0BF99F9A4B0",
 -4122 => x"C0C0C0BF99F9A4A4",
 -4121 => x"C0C0C0BF99F9A4F9",
 -4120 => x"C0C0C0BF99F9A4C0",
 -4119 => x"C0C0C0BF99F9F990",
 -4118 => x"C0C0C0BF99F9F980",
 -4117 => x"C0C0C0BF99F9F9F8",
 -4116 => x"C0C0C0BF99F9F982",
 -4115 => x"C0C0C0BF99F9F992",
 -4114 => x"C0C0C0BF99F9F999",
 -4113 => x"C0C0C0BF99F9F9B0",
 -4112 => x"C0C0C0BF99F9F9A4",
 -4111 => x"C0C0C0BF99F9F9F9",
 -4110 => x"C0C0C0BF99F9F9C0",
 -4109 => x"C0C0C0BF99F9C090",
 -4108 => x"C0C0C0BF99F9C080",
 -4107 => x"C0C0C0BF99F9C0F8",
 -4106 => x"C0C0C0BF99F9C082",
 -4105 => x"C0C0C0BF99F9C092",
 -4104 => x"C0C0C0BF99F9C099",
 -4103 => x"C0C0C0BF99F9C0B0",
 -4102 => x"C0C0C0BF99F9C0A4",
 -4101 => x"C0C0C0BF99F9C0F9",
 -4100 => x"C0C0C0BF99F9C0C0",
 -4099 => x"C0C0C0BF99C09090",
 -4098 => x"C0C0C0BF99C09080",
 -4097 => x"C0C0C0BF99C090F8",
 -4096 => x"C0C0C0BF99C09082",
 -4095 => x"C0C0C0BF99C09092",
 -4094 => x"C0C0C0BF99C09099",
 -4093 => x"C0C0C0BF99C090B0",
 -4092 => x"C0C0C0BF99C090A4",
 -4091 => x"C0C0C0BF99C090F9",
 -4090 => x"C0C0C0BF99C090C0",
 -4089 => x"C0C0C0BF99C08090",
 -4088 => x"C0C0C0BF99C08080",
 -4087 => x"C0C0C0BF99C080F8",
 -4086 => x"C0C0C0BF99C08082",
 -4085 => x"C0C0C0BF99C08092",
 -4084 => x"C0C0C0BF99C08099",
 -4083 => x"C0C0C0BF99C080B0",
 -4082 => x"C0C0C0BF99C080A4",
 -4081 => x"C0C0C0BF99C080F9",
 -4080 => x"C0C0C0BF99C080C0",
 -4079 => x"C0C0C0BF99C0F890",
 -4078 => x"C0C0C0BF99C0F880",
 -4077 => x"C0C0C0BF99C0F8F8",
 -4076 => x"C0C0C0BF99C0F882",
 -4075 => x"C0C0C0BF99C0F892",
 -4074 => x"C0C0C0BF99C0F899",
 -4073 => x"C0C0C0BF99C0F8B0",
 -4072 => x"C0C0C0BF99C0F8A4",
 -4071 => x"C0C0C0BF99C0F8F9",
 -4070 => x"C0C0C0BF99C0F8C0",
 -4069 => x"C0C0C0BF99C08290",
 -4068 => x"C0C0C0BF99C08280",
 -4067 => x"C0C0C0BF99C082F8",
 -4066 => x"C0C0C0BF99C08282",
 -4065 => x"C0C0C0BF99C08292",
 -4064 => x"C0C0C0BF99C08299",
 -4063 => x"C0C0C0BF99C082B0",
 -4062 => x"C0C0C0BF99C082A4",
 -4061 => x"C0C0C0BF99C082F9",
 -4060 => x"C0C0C0BF99C082C0",
 -4059 => x"C0C0C0BF99C09290",
 -4058 => x"C0C0C0BF99C09280",
 -4057 => x"C0C0C0BF99C092F8",
 -4056 => x"C0C0C0BF99C09282",
 -4055 => x"C0C0C0BF99C09292",
 -4054 => x"C0C0C0BF99C09299",
 -4053 => x"C0C0C0BF99C092B0",
 -4052 => x"C0C0C0BF99C092A4",
 -4051 => x"C0C0C0BF99C092F9",
 -4050 => x"C0C0C0BF99C092C0",
 -4049 => x"C0C0C0BF99C09990",
 -4048 => x"C0C0C0BF99C09980",
 -4047 => x"C0C0C0BF99C099F8",
 -4046 => x"C0C0C0BF99C09982",
 -4045 => x"C0C0C0BF99C09992",
 -4044 => x"C0C0C0BF99C09999",
 -4043 => x"C0C0C0BF99C099B0",
 -4042 => x"C0C0C0BF99C099A4",
 -4041 => x"C0C0C0BF99C099F9",
 -4040 => x"C0C0C0BF99C099C0",
 -4039 => x"C0C0C0BF99C0B090",
 -4038 => x"C0C0C0BF99C0B080",
 -4037 => x"C0C0C0BF99C0B0F8",
 -4036 => x"C0C0C0BF99C0B082",
 -4035 => x"C0C0C0BF99C0B092",
 -4034 => x"C0C0C0BF99C0B099",
 -4033 => x"C0C0C0BF99C0B0B0",
 -4032 => x"C0C0C0BF99C0B0A4",
 -4031 => x"C0C0C0BF99C0B0F9",
 -4030 => x"C0C0C0BF99C0B0C0",
 -4029 => x"C0C0C0BF99C0A490",
 -4028 => x"C0C0C0BF99C0A480",
 -4027 => x"C0C0C0BF99C0A4F8",
 -4026 => x"C0C0C0BF99C0A482",
 -4025 => x"C0C0C0BF99C0A492",
 -4024 => x"C0C0C0BF99C0A499",
 -4023 => x"C0C0C0BF99C0A4B0",
 -4022 => x"C0C0C0BF99C0A4A4",
 -4021 => x"C0C0C0BF99C0A4F9",
 -4020 => x"C0C0C0BF99C0A4C0",
 -4019 => x"C0C0C0BF99C0F990",
 -4018 => x"C0C0C0BF99C0F980",
 -4017 => x"C0C0C0BF99C0F9F8",
 -4016 => x"C0C0C0BF99C0F982",
 -4015 => x"C0C0C0BF99C0F992",
 -4014 => x"C0C0C0BF99C0F999",
 -4013 => x"C0C0C0BF99C0F9B0",
 -4012 => x"C0C0C0BF99C0F9A4",
 -4011 => x"C0C0C0BF99C0F9F9",
 -4010 => x"C0C0C0BF99C0F9C0",
 -4009 => x"C0C0C0BF99C0C090",
 -4008 => x"C0C0C0BF99C0C080",
 -4007 => x"C0C0C0BF99C0C0F8",
 -4006 => x"C0C0C0BF99C0C082",
 -4005 => x"C0C0C0BF99C0C092",
 -4004 => x"C0C0C0BF99C0C099",
 -4003 => x"C0C0C0BF99C0C0B0",
 -4002 => x"C0C0C0BF99C0C0A4",
 -4001 => x"C0C0C0BF99C0C0F9",
 -4000 => x"C0C0C0BF99C0C0C0",
 -3999 => x"C0C0C0BFB0909090",
 -3998 => x"C0C0C0BFB0909080",
 -3997 => x"C0C0C0BFB09090F8",
 -3996 => x"C0C0C0BFB0909082",
 -3995 => x"C0C0C0BFB0909092",
 -3994 => x"C0C0C0BFB0909099",
 -3993 => x"C0C0C0BFB09090B0",
 -3992 => x"C0C0C0BFB09090A4",
 -3991 => x"C0C0C0BFB09090F9",
 -3990 => x"C0C0C0BFB09090C0",
 -3989 => x"C0C0C0BFB0908090",
 -3988 => x"C0C0C0BFB0908080",
 -3987 => x"C0C0C0BFB09080F8",
 -3986 => x"C0C0C0BFB0908082",
 -3985 => x"C0C0C0BFB0908092",
 -3984 => x"C0C0C0BFB0908099",
 -3983 => x"C0C0C0BFB09080B0",
 -3982 => x"C0C0C0BFB09080A4",
 -3981 => x"C0C0C0BFB09080F9",
 -3980 => x"C0C0C0BFB09080C0",
 -3979 => x"C0C0C0BFB090F890",
 -3978 => x"C0C0C0BFB090F880",
 -3977 => x"C0C0C0BFB090F8F8",
 -3976 => x"C0C0C0BFB090F882",
 -3975 => x"C0C0C0BFB090F892",
 -3974 => x"C0C0C0BFB090F899",
 -3973 => x"C0C0C0BFB090F8B0",
 -3972 => x"C0C0C0BFB090F8A4",
 -3971 => x"C0C0C0BFB090F8F9",
 -3970 => x"C0C0C0BFB090F8C0",
 -3969 => x"C0C0C0BFB0908290",
 -3968 => x"C0C0C0BFB0908280",
 -3967 => x"C0C0C0BFB09082F8",
 -3966 => x"C0C0C0BFB0908282",
 -3965 => x"C0C0C0BFB0908292",
 -3964 => x"C0C0C0BFB0908299",
 -3963 => x"C0C0C0BFB09082B0",
 -3962 => x"C0C0C0BFB09082A4",
 -3961 => x"C0C0C0BFB09082F9",
 -3960 => x"C0C0C0BFB09082C0",
 -3959 => x"C0C0C0BFB0909290",
 -3958 => x"C0C0C0BFB0909280",
 -3957 => x"C0C0C0BFB09092F8",
 -3956 => x"C0C0C0BFB0909282",
 -3955 => x"C0C0C0BFB0909292",
 -3954 => x"C0C0C0BFB0909299",
 -3953 => x"C0C0C0BFB09092B0",
 -3952 => x"C0C0C0BFB09092A4",
 -3951 => x"C0C0C0BFB09092F9",
 -3950 => x"C0C0C0BFB09092C0",
 -3949 => x"C0C0C0BFB0909990",
 -3948 => x"C0C0C0BFB0909980",
 -3947 => x"C0C0C0BFB09099F8",
 -3946 => x"C0C0C0BFB0909982",
 -3945 => x"C0C0C0BFB0909992",
 -3944 => x"C0C0C0BFB0909999",
 -3943 => x"C0C0C0BFB09099B0",
 -3942 => x"C0C0C0BFB09099A4",
 -3941 => x"C0C0C0BFB09099F9",
 -3940 => x"C0C0C0BFB09099C0",
 -3939 => x"C0C0C0BFB090B090",
 -3938 => x"C0C0C0BFB090B080",
 -3937 => x"C0C0C0BFB090B0F8",
 -3936 => x"C0C0C0BFB090B082",
 -3935 => x"C0C0C0BFB090B092",
 -3934 => x"C0C0C0BFB090B099",
 -3933 => x"C0C0C0BFB090B0B0",
 -3932 => x"C0C0C0BFB090B0A4",
 -3931 => x"C0C0C0BFB090B0F9",
 -3930 => x"C0C0C0BFB090B0C0",
 -3929 => x"C0C0C0BFB090A490",
 -3928 => x"C0C0C0BFB090A480",
 -3927 => x"C0C0C0BFB090A4F8",
 -3926 => x"C0C0C0BFB090A482",
 -3925 => x"C0C0C0BFB090A492",
 -3924 => x"C0C0C0BFB090A499",
 -3923 => x"C0C0C0BFB090A4B0",
 -3922 => x"C0C0C0BFB090A4A4",
 -3921 => x"C0C0C0BFB090A4F9",
 -3920 => x"C0C0C0BFB090A4C0",
 -3919 => x"C0C0C0BFB090F990",
 -3918 => x"C0C0C0BFB090F980",
 -3917 => x"C0C0C0BFB090F9F8",
 -3916 => x"C0C0C0BFB090F982",
 -3915 => x"C0C0C0BFB090F992",
 -3914 => x"C0C0C0BFB090F999",
 -3913 => x"C0C0C0BFB090F9B0",
 -3912 => x"C0C0C0BFB090F9A4",
 -3911 => x"C0C0C0BFB090F9F9",
 -3910 => x"C0C0C0BFB090F9C0",
 -3909 => x"C0C0C0BFB090C090",
 -3908 => x"C0C0C0BFB090C080",
 -3907 => x"C0C0C0BFB090C0F8",
 -3906 => x"C0C0C0BFB090C082",
 -3905 => x"C0C0C0BFB090C092",
 -3904 => x"C0C0C0BFB090C099",
 -3903 => x"C0C0C0BFB090C0B0",
 -3902 => x"C0C0C0BFB090C0A4",
 -3901 => x"C0C0C0BFB090C0F9",
 -3900 => x"C0C0C0BFB090C0C0",
 -3899 => x"C0C0C0BFB0809090",
 -3898 => x"C0C0C0BFB0809080",
 -3897 => x"C0C0C0BFB08090F8",
 -3896 => x"C0C0C0BFB0809082",
 -3895 => x"C0C0C0BFB0809092",
 -3894 => x"C0C0C0BFB0809099",
 -3893 => x"C0C0C0BFB08090B0",
 -3892 => x"C0C0C0BFB08090A4",
 -3891 => x"C0C0C0BFB08090F9",
 -3890 => x"C0C0C0BFB08090C0",
 -3889 => x"C0C0C0BFB0808090",
 -3888 => x"C0C0C0BFB0808080",
 -3887 => x"C0C0C0BFB08080F8",
 -3886 => x"C0C0C0BFB0808082",
 -3885 => x"C0C0C0BFB0808092",
 -3884 => x"C0C0C0BFB0808099",
 -3883 => x"C0C0C0BFB08080B0",
 -3882 => x"C0C0C0BFB08080A4",
 -3881 => x"C0C0C0BFB08080F9",
 -3880 => x"C0C0C0BFB08080C0",
 -3879 => x"C0C0C0BFB080F890",
 -3878 => x"C0C0C0BFB080F880",
 -3877 => x"C0C0C0BFB080F8F8",
 -3876 => x"C0C0C0BFB080F882",
 -3875 => x"C0C0C0BFB080F892",
 -3874 => x"C0C0C0BFB080F899",
 -3873 => x"C0C0C0BFB080F8B0",
 -3872 => x"C0C0C0BFB080F8A4",
 -3871 => x"C0C0C0BFB080F8F9",
 -3870 => x"C0C0C0BFB080F8C0",
 -3869 => x"C0C0C0BFB0808290",
 -3868 => x"C0C0C0BFB0808280",
 -3867 => x"C0C0C0BFB08082F8",
 -3866 => x"C0C0C0BFB0808282",
 -3865 => x"C0C0C0BFB0808292",
 -3864 => x"C0C0C0BFB0808299",
 -3863 => x"C0C0C0BFB08082B0",
 -3862 => x"C0C0C0BFB08082A4",
 -3861 => x"C0C0C0BFB08082F9",
 -3860 => x"C0C0C0BFB08082C0",
 -3859 => x"C0C0C0BFB0809290",
 -3858 => x"C0C0C0BFB0809280",
 -3857 => x"C0C0C0BFB08092F8",
 -3856 => x"C0C0C0BFB0809282",
 -3855 => x"C0C0C0BFB0809292",
 -3854 => x"C0C0C0BFB0809299",
 -3853 => x"C0C0C0BFB08092B0",
 -3852 => x"C0C0C0BFB08092A4",
 -3851 => x"C0C0C0BFB08092F9",
 -3850 => x"C0C0C0BFB08092C0",
 -3849 => x"C0C0C0BFB0809990",
 -3848 => x"C0C0C0BFB0809980",
 -3847 => x"C0C0C0BFB08099F8",
 -3846 => x"C0C0C0BFB0809982",
 -3845 => x"C0C0C0BFB0809992",
 -3844 => x"C0C0C0BFB0809999",
 -3843 => x"C0C0C0BFB08099B0",
 -3842 => x"C0C0C0BFB08099A4",
 -3841 => x"C0C0C0BFB08099F9",
 -3840 => x"C0C0C0BFB08099C0",
 -3839 => x"C0C0C0BFB080B090",
 -3838 => x"C0C0C0BFB080B080",
 -3837 => x"C0C0C0BFB080B0F8",
 -3836 => x"C0C0C0BFB080B082",
 -3835 => x"C0C0C0BFB080B092",
 -3834 => x"C0C0C0BFB080B099",
 -3833 => x"C0C0C0BFB080B0B0",
 -3832 => x"C0C0C0BFB080B0A4",
 -3831 => x"C0C0C0BFB080B0F9",
 -3830 => x"C0C0C0BFB080B0C0",
 -3829 => x"C0C0C0BFB080A490",
 -3828 => x"C0C0C0BFB080A480",
 -3827 => x"C0C0C0BFB080A4F8",
 -3826 => x"C0C0C0BFB080A482",
 -3825 => x"C0C0C0BFB080A492",
 -3824 => x"C0C0C0BFB080A499",
 -3823 => x"C0C0C0BFB080A4B0",
 -3822 => x"C0C0C0BFB080A4A4",
 -3821 => x"C0C0C0BFB080A4F9",
 -3820 => x"C0C0C0BFB080A4C0",
 -3819 => x"C0C0C0BFB080F990",
 -3818 => x"C0C0C0BFB080F980",
 -3817 => x"C0C0C0BFB080F9F8",
 -3816 => x"C0C0C0BFB080F982",
 -3815 => x"C0C0C0BFB080F992",
 -3814 => x"C0C0C0BFB080F999",
 -3813 => x"C0C0C0BFB080F9B0",
 -3812 => x"C0C0C0BFB080F9A4",
 -3811 => x"C0C0C0BFB080F9F9",
 -3810 => x"C0C0C0BFB080F9C0",
 -3809 => x"C0C0C0BFB080C090",
 -3808 => x"C0C0C0BFB080C080",
 -3807 => x"C0C0C0BFB080C0F8",
 -3806 => x"C0C0C0BFB080C082",
 -3805 => x"C0C0C0BFB080C092",
 -3804 => x"C0C0C0BFB080C099",
 -3803 => x"C0C0C0BFB080C0B0",
 -3802 => x"C0C0C0BFB080C0A4",
 -3801 => x"C0C0C0BFB080C0F9",
 -3800 => x"C0C0C0BFB080C0C0",
 -3799 => x"C0C0C0BFB0F89090",
 -3798 => x"C0C0C0BFB0F89080",
 -3797 => x"C0C0C0BFB0F890F8",
 -3796 => x"C0C0C0BFB0F89082",
 -3795 => x"C0C0C0BFB0F89092",
 -3794 => x"C0C0C0BFB0F89099",
 -3793 => x"C0C0C0BFB0F890B0",
 -3792 => x"C0C0C0BFB0F890A4",
 -3791 => x"C0C0C0BFB0F890F9",
 -3790 => x"C0C0C0BFB0F890C0",
 -3789 => x"C0C0C0BFB0F88090",
 -3788 => x"C0C0C0BFB0F88080",
 -3787 => x"C0C0C0BFB0F880F8",
 -3786 => x"C0C0C0BFB0F88082",
 -3785 => x"C0C0C0BFB0F88092",
 -3784 => x"C0C0C0BFB0F88099",
 -3783 => x"C0C0C0BFB0F880B0",
 -3782 => x"C0C0C0BFB0F880A4",
 -3781 => x"C0C0C0BFB0F880F9",
 -3780 => x"C0C0C0BFB0F880C0",
 -3779 => x"C0C0C0BFB0F8F890",
 -3778 => x"C0C0C0BFB0F8F880",
 -3777 => x"C0C0C0BFB0F8F8F8",
 -3776 => x"C0C0C0BFB0F8F882",
 -3775 => x"C0C0C0BFB0F8F892",
 -3774 => x"C0C0C0BFB0F8F899",
 -3773 => x"C0C0C0BFB0F8F8B0",
 -3772 => x"C0C0C0BFB0F8F8A4",
 -3771 => x"C0C0C0BFB0F8F8F9",
 -3770 => x"C0C0C0BFB0F8F8C0",
 -3769 => x"C0C0C0BFB0F88290",
 -3768 => x"C0C0C0BFB0F88280",
 -3767 => x"C0C0C0BFB0F882F8",
 -3766 => x"C0C0C0BFB0F88282",
 -3765 => x"C0C0C0BFB0F88292",
 -3764 => x"C0C0C0BFB0F88299",
 -3763 => x"C0C0C0BFB0F882B0",
 -3762 => x"C0C0C0BFB0F882A4",
 -3761 => x"C0C0C0BFB0F882F9",
 -3760 => x"C0C0C0BFB0F882C0",
 -3759 => x"C0C0C0BFB0F89290",
 -3758 => x"C0C0C0BFB0F89280",
 -3757 => x"C0C0C0BFB0F892F8",
 -3756 => x"C0C0C0BFB0F89282",
 -3755 => x"C0C0C0BFB0F89292",
 -3754 => x"C0C0C0BFB0F89299",
 -3753 => x"C0C0C0BFB0F892B0",
 -3752 => x"C0C0C0BFB0F892A4",
 -3751 => x"C0C0C0BFB0F892F9",
 -3750 => x"C0C0C0BFB0F892C0",
 -3749 => x"C0C0C0BFB0F89990",
 -3748 => x"C0C0C0BFB0F89980",
 -3747 => x"C0C0C0BFB0F899F8",
 -3746 => x"C0C0C0BFB0F89982",
 -3745 => x"C0C0C0BFB0F89992",
 -3744 => x"C0C0C0BFB0F89999",
 -3743 => x"C0C0C0BFB0F899B0",
 -3742 => x"C0C0C0BFB0F899A4",
 -3741 => x"C0C0C0BFB0F899F9",
 -3740 => x"C0C0C0BFB0F899C0",
 -3739 => x"C0C0C0BFB0F8B090",
 -3738 => x"C0C0C0BFB0F8B080",
 -3737 => x"C0C0C0BFB0F8B0F8",
 -3736 => x"C0C0C0BFB0F8B082",
 -3735 => x"C0C0C0BFB0F8B092",
 -3734 => x"C0C0C0BFB0F8B099",
 -3733 => x"C0C0C0BFB0F8B0B0",
 -3732 => x"C0C0C0BFB0F8B0A4",
 -3731 => x"C0C0C0BFB0F8B0F9",
 -3730 => x"C0C0C0BFB0F8B0C0",
 -3729 => x"C0C0C0BFB0F8A490",
 -3728 => x"C0C0C0BFB0F8A480",
 -3727 => x"C0C0C0BFB0F8A4F8",
 -3726 => x"C0C0C0BFB0F8A482",
 -3725 => x"C0C0C0BFB0F8A492",
 -3724 => x"C0C0C0BFB0F8A499",
 -3723 => x"C0C0C0BFB0F8A4B0",
 -3722 => x"C0C0C0BFB0F8A4A4",
 -3721 => x"C0C0C0BFB0F8A4F9",
 -3720 => x"C0C0C0BFB0F8A4C0",
 -3719 => x"C0C0C0BFB0F8F990",
 -3718 => x"C0C0C0BFB0F8F980",
 -3717 => x"C0C0C0BFB0F8F9F8",
 -3716 => x"C0C0C0BFB0F8F982",
 -3715 => x"C0C0C0BFB0F8F992",
 -3714 => x"C0C0C0BFB0F8F999",
 -3713 => x"C0C0C0BFB0F8F9B0",
 -3712 => x"C0C0C0BFB0F8F9A4",
 -3711 => x"C0C0C0BFB0F8F9F9",
 -3710 => x"C0C0C0BFB0F8F9C0",
 -3709 => x"C0C0C0BFB0F8C090",
 -3708 => x"C0C0C0BFB0F8C080",
 -3707 => x"C0C0C0BFB0F8C0F8",
 -3706 => x"C0C0C0BFB0F8C082",
 -3705 => x"C0C0C0BFB0F8C092",
 -3704 => x"C0C0C0BFB0F8C099",
 -3703 => x"C0C0C0BFB0F8C0B0",
 -3702 => x"C0C0C0BFB0F8C0A4",
 -3701 => x"C0C0C0BFB0F8C0F9",
 -3700 => x"C0C0C0BFB0F8C0C0",
 -3699 => x"C0C0C0BFB0829090",
 -3698 => x"C0C0C0BFB0829080",
 -3697 => x"C0C0C0BFB08290F8",
 -3696 => x"C0C0C0BFB0829082",
 -3695 => x"C0C0C0BFB0829092",
 -3694 => x"C0C0C0BFB0829099",
 -3693 => x"C0C0C0BFB08290B0",
 -3692 => x"C0C0C0BFB08290A4",
 -3691 => x"C0C0C0BFB08290F9",
 -3690 => x"C0C0C0BFB08290C0",
 -3689 => x"C0C0C0BFB0828090",
 -3688 => x"C0C0C0BFB0828080",
 -3687 => x"C0C0C0BFB08280F8",
 -3686 => x"C0C0C0BFB0828082",
 -3685 => x"C0C0C0BFB0828092",
 -3684 => x"C0C0C0BFB0828099",
 -3683 => x"C0C0C0BFB08280B0",
 -3682 => x"C0C0C0BFB08280A4",
 -3681 => x"C0C0C0BFB08280F9",
 -3680 => x"C0C0C0BFB08280C0",
 -3679 => x"C0C0C0BFB082F890",
 -3678 => x"C0C0C0BFB082F880",
 -3677 => x"C0C0C0BFB082F8F8",
 -3676 => x"C0C0C0BFB082F882",
 -3675 => x"C0C0C0BFB082F892",
 -3674 => x"C0C0C0BFB082F899",
 -3673 => x"C0C0C0BFB082F8B0",
 -3672 => x"C0C0C0BFB082F8A4",
 -3671 => x"C0C0C0BFB082F8F9",
 -3670 => x"C0C0C0BFB082F8C0",
 -3669 => x"C0C0C0BFB0828290",
 -3668 => x"C0C0C0BFB0828280",
 -3667 => x"C0C0C0BFB08282F8",
 -3666 => x"C0C0C0BFB0828282",
 -3665 => x"C0C0C0BFB0828292",
 -3664 => x"C0C0C0BFB0828299",
 -3663 => x"C0C0C0BFB08282B0",
 -3662 => x"C0C0C0BFB08282A4",
 -3661 => x"C0C0C0BFB08282F9",
 -3660 => x"C0C0C0BFB08282C0",
 -3659 => x"C0C0C0BFB0829290",
 -3658 => x"C0C0C0BFB0829280",
 -3657 => x"C0C0C0BFB08292F8",
 -3656 => x"C0C0C0BFB0829282",
 -3655 => x"C0C0C0BFB0829292",
 -3654 => x"C0C0C0BFB0829299",
 -3653 => x"C0C0C0BFB08292B0",
 -3652 => x"C0C0C0BFB08292A4",
 -3651 => x"C0C0C0BFB08292F9",
 -3650 => x"C0C0C0BFB08292C0",
 -3649 => x"C0C0C0BFB0829990",
 -3648 => x"C0C0C0BFB0829980",
 -3647 => x"C0C0C0BFB08299F8",
 -3646 => x"C0C0C0BFB0829982",
 -3645 => x"C0C0C0BFB0829992",
 -3644 => x"C0C0C0BFB0829999",
 -3643 => x"C0C0C0BFB08299B0",
 -3642 => x"C0C0C0BFB08299A4",
 -3641 => x"C0C0C0BFB08299F9",
 -3640 => x"C0C0C0BFB08299C0",
 -3639 => x"C0C0C0BFB082B090",
 -3638 => x"C0C0C0BFB082B080",
 -3637 => x"C0C0C0BFB082B0F8",
 -3636 => x"C0C0C0BFB082B082",
 -3635 => x"C0C0C0BFB082B092",
 -3634 => x"C0C0C0BFB082B099",
 -3633 => x"C0C0C0BFB082B0B0",
 -3632 => x"C0C0C0BFB082B0A4",
 -3631 => x"C0C0C0BFB082B0F9",
 -3630 => x"C0C0C0BFB082B0C0",
 -3629 => x"C0C0C0BFB082A490",
 -3628 => x"C0C0C0BFB082A480",
 -3627 => x"C0C0C0BFB082A4F8",
 -3626 => x"C0C0C0BFB082A482",
 -3625 => x"C0C0C0BFB082A492",
 -3624 => x"C0C0C0BFB082A499",
 -3623 => x"C0C0C0BFB082A4B0",
 -3622 => x"C0C0C0BFB082A4A4",
 -3621 => x"C0C0C0BFB082A4F9",
 -3620 => x"C0C0C0BFB082A4C0",
 -3619 => x"C0C0C0BFB082F990",
 -3618 => x"C0C0C0BFB082F980",
 -3617 => x"C0C0C0BFB082F9F8",
 -3616 => x"C0C0C0BFB082F982",
 -3615 => x"C0C0C0BFB082F992",
 -3614 => x"C0C0C0BFB082F999",
 -3613 => x"C0C0C0BFB082F9B0",
 -3612 => x"C0C0C0BFB082F9A4",
 -3611 => x"C0C0C0BFB082F9F9",
 -3610 => x"C0C0C0BFB082F9C0",
 -3609 => x"C0C0C0BFB082C090",
 -3608 => x"C0C0C0BFB082C080",
 -3607 => x"C0C0C0BFB082C0F8",
 -3606 => x"C0C0C0BFB082C082",
 -3605 => x"C0C0C0BFB082C092",
 -3604 => x"C0C0C0BFB082C099",
 -3603 => x"C0C0C0BFB082C0B0",
 -3602 => x"C0C0C0BFB082C0A4",
 -3601 => x"C0C0C0BFB082C0F9",
 -3600 => x"C0C0C0BFB082C0C0",
 -3599 => x"C0C0C0BFB0929090",
 -3598 => x"C0C0C0BFB0929080",
 -3597 => x"C0C0C0BFB09290F8",
 -3596 => x"C0C0C0BFB0929082",
 -3595 => x"C0C0C0BFB0929092",
 -3594 => x"C0C0C0BFB0929099",
 -3593 => x"C0C0C0BFB09290B0",
 -3592 => x"C0C0C0BFB09290A4",
 -3591 => x"C0C0C0BFB09290F9",
 -3590 => x"C0C0C0BFB09290C0",
 -3589 => x"C0C0C0BFB0928090",
 -3588 => x"C0C0C0BFB0928080",
 -3587 => x"C0C0C0BFB09280F8",
 -3586 => x"C0C0C0BFB0928082",
 -3585 => x"C0C0C0BFB0928092",
 -3584 => x"C0C0C0BFB0928099",
 -3583 => x"C0C0C0BFB09280B0",
 -3582 => x"C0C0C0BFB09280A4",
 -3581 => x"C0C0C0BFB09280F9",
 -3580 => x"C0C0C0BFB09280C0",
 -3579 => x"C0C0C0BFB092F890",
 -3578 => x"C0C0C0BFB092F880",
 -3577 => x"C0C0C0BFB092F8F8",
 -3576 => x"C0C0C0BFB092F882",
 -3575 => x"C0C0C0BFB092F892",
 -3574 => x"C0C0C0BFB092F899",
 -3573 => x"C0C0C0BFB092F8B0",
 -3572 => x"C0C0C0BFB092F8A4",
 -3571 => x"C0C0C0BFB092F8F9",
 -3570 => x"C0C0C0BFB092F8C0",
 -3569 => x"C0C0C0BFB0928290",
 -3568 => x"C0C0C0BFB0928280",
 -3567 => x"C0C0C0BFB09282F8",
 -3566 => x"C0C0C0BFB0928282",
 -3565 => x"C0C0C0BFB0928292",
 -3564 => x"C0C0C0BFB0928299",
 -3563 => x"C0C0C0BFB09282B0",
 -3562 => x"C0C0C0BFB09282A4",
 -3561 => x"C0C0C0BFB09282F9",
 -3560 => x"C0C0C0BFB09282C0",
 -3559 => x"C0C0C0BFB0929290",
 -3558 => x"C0C0C0BFB0929280",
 -3557 => x"C0C0C0BFB09292F8",
 -3556 => x"C0C0C0BFB0929282",
 -3555 => x"C0C0C0BFB0929292",
 -3554 => x"C0C0C0BFB0929299",
 -3553 => x"C0C0C0BFB09292B0",
 -3552 => x"C0C0C0BFB09292A4",
 -3551 => x"C0C0C0BFB09292F9",
 -3550 => x"C0C0C0BFB09292C0",
 -3549 => x"C0C0C0BFB0929990",
 -3548 => x"C0C0C0BFB0929980",
 -3547 => x"C0C0C0BFB09299F8",
 -3546 => x"C0C0C0BFB0929982",
 -3545 => x"C0C0C0BFB0929992",
 -3544 => x"C0C0C0BFB0929999",
 -3543 => x"C0C0C0BFB09299B0",
 -3542 => x"C0C0C0BFB09299A4",
 -3541 => x"C0C0C0BFB09299F9",
 -3540 => x"C0C0C0BFB09299C0",
 -3539 => x"C0C0C0BFB092B090",
 -3538 => x"C0C0C0BFB092B080",
 -3537 => x"C0C0C0BFB092B0F8",
 -3536 => x"C0C0C0BFB092B082",
 -3535 => x"C0C0C0BFB092B092",
 -3534 => x"C0C0C0BFB092B099",
 -3533 => x"C0C0C0BFB092B0B0",
 -3532 => x"C0C0C0BFB092B0A4",
 -3531 => x"C0C0C0BFB092B0F9",
 -3530 => x"C0C0C0BFB092B0C0",
 -3529 => x"C0C0C0BFB092A490",
 -3528 => x"C0C0C0BFB092A480",
 -3527 => x"C0C0C0BFB092A4F8",
 -3526 => x"C0C0C0BFB092A482",
 -3525 => x"C0C0C0BFB092A492",
 -3524 => x"C0C0C0BFB092A499",
 -3523 => x"C0C0C0BFB092A4B0",
 -3522 => x"C0C0C0BFB092A4A4",
 -3521 => x"C0C0C0BFB092A4F9",
 -3520 => x"C0C0C0BFB092A4C0",
 -3519 => x"C0C0C0BFB092F990",
 -3518 => x"C0C0C0BFB092F980",
 -3517 => x"C0C0C0BFB092F9F8",
 -3516 => x"C0C0C0BFB092F982",
 -3515 => x"C0C0C0BFB092F992",
 -3514 => x"C0C0C0BFB092F999",
 -3513 => x"C0C0C0BFB092F9B0",
 -3512 => x"C0C0C0BFB092F9A4",
 -3511 => x"C0C0C0BFB092F9F9",
 -3510 => x"C0C0C0BFB092F9C0",
 -3509 => x"C0C0C0BFB092C090",
 -3508 => x"C0C0C0BFB092C080",
 -3507 => x"C0C0C0BFB092C0F8",
 -3506 => x"C0C0C0BFB092C082",
 -3505 => x"C0C0C0BFB092C092",
 -3504 => x"C0C0C0BFB092C099",
 -3503 => x"C0C0C0BFB092C0B0",
 -3502 => x"C0C0C0BFB092C0A4",
 -3501 => x"C0C0C0BFB092C0F9",
 -3500 => x"C0C0C0BFB092C0C0",
 -3499 => x"C0C0C0BFB0999090",
 -3498 => x"C0C0C0BFB0999080",
 -3497 => x"C0C0C0BFB09990F8",
 -3496 => x"C0C0C0BFB0999082",
 -3495 => x"C0C0C0BFB0999092",
 -3494 => x"C0C0C0BFB0999099",
 -3493 => x"C0C0C0BFB09990B0",
 -3492 => x"C0C0C0BFB09990A4",
 -3491 => x"C0C0C0BFB09990F9",
 -3490 => x"C0C0C0BFB09990C0",
 -3489 => x"C0C0C0BFB0998090",
 -3488 => x"C0C0C0BFB0998080",
 -3487 => x"C0C0C0BFB09980F8",
 -3486 => x"C0C0C0BFB0998082",
 -3485 => x"C0C0C0BFB0998092",
 -3484 => x"C0C0C0BFB0998099",
 -3483 => x"C0C0C0BFB09980B0",
 -3482 => x"C0C0C0BFB09980A4",
 -3481 => x"C0C0C0BFB09980F9",
 -3480 => x"C0C0C0BFB09980C0",
 -3479 => x"C0C0C0BFB099F890",
 -3478 => x"C0C0C0BFB099F880",
 -3477 => x"C0C0C0BFB099F8F8",
 -3476 => x"C0C0C0BFB099F882",
 -3475 => x"C0C0C0BFB099F892",
 -3474 => x"C0C0C0BFB099F899",
 -3473 => x"C0C0C0BFB099F8B0",
 -3472 => x"C0C0C0BFB099F8A4",
 -3471 => x"C0C0C0BFB099F8F9",
 -3470 => x"C0C0C0BFB099F8C0",
 -3469 => x"C0C0C0BFB0998290",
 -3468 => x"C0C0C0BFB0998280",
 -3467 => x"C0C0C0BFB09982F8",
 -3466 => x"C0C0C0BFB0998282",
 -3465 => x"C0C0C0BFB0998292",
 -3464 => x"C0C0C0BFB0998299",
 -3463 => x"C0C0C0BFB09982B0",
 -3462 => x"C0C0C0BFB09982A4",
 -3461 => x"C0C0C0BFB09982F9",
 -3460 => x"C0C0C0BFB09982C0",
 -3459 => x"C0C0C0BFB0999290",
 -3458 => x"C0C0C0BFB0999280",
 -3457 => x"C0C0C0BFB09992F8",
 -3456 => x"C0C0C0BFB0999282",
 -3455 => x"C0C0C0BFB0999292",
 -3454 => x"C0C0C0BFB0999299",
 -3453 => x"C0C0C0BFB09992B0",
 -3452 => x"C0C0C0BFB09992A4",
 -3451 => x"C0C0C0BFB09992F9",
 -3450 => x"C0C0C0BFB09992C0",
 -3449 => x"C0C0C0BFB0999990",
 -3448 => x"C0C0C0BFB0999980",
 -3447 => x"C0C0C0BFB09999F8",
 -3446 => x"C0C0C0BFB0999982",
 -3445 => x"C0C0C0BFB0999992",
 -3444 => x"C0C0C0BFB0999999",
 -3443 => x"C0C0C0BFB09999B0",
 -3442 => x"C0C0C0BFB09999A4",
 -3441 => x"C0C0C0BFB09999F9",
 -3440 => x"C0C0C0BFB09999C0",
 -3439 => x"C0C0C0BFB099B090",
 -3438 => x"C0C0C0BFB099B080",
 -3437 => x"C0C0C0BFB099B0F8",
 -3436 => x"C0C0C0BFB099B082",
 -3435 => x"C0C0C0BFB099B092",
 -3434 => x"C0C0C0BFB099B099",
 -3433 => x"C0C0C0BFB099B0B0",
 -3432 => x"C0C0C0BFB099B0A4",
 -3431 => x"C0C0C0BFB099B0F9",
 -3430 => x"C0C0C0BFB099B0C0",
 -3429 => x"C0C0C0BFB099A490",
 -3428 => x"C0C0C0BFB099A480",
 -3427 => x"C0C0C0BFB099A4F8",
 -3426 => x"C0C0C0BFB099A482",
 -3425 => x"C0C0C0BFB099A492",
 -3424 => x"C0C0C0BFB099A499",
 -3423 => x"C0C0C0BFB099A4B0",
 -3422 => x"C0C0C0BFB099A4A4",
 -3421 => x"C0C0C0BFB099A4F9",
 -3420 => x"C0C0C0BFB099A4C0",
 -3419 => x"C0C0C0BFB099F990",
 -3418 => x"C0C0C0BFB099F980",
 -3417 => x"C0C0C0BFB099F9F8",
 -3416 => x"C0C0C0BFB099F982",
 -3415 => x"C0C0C0BFB099F992",
 -3414 => x"C0C0C0BFB099F999",
 -3413 => x"C0C0C0BFB099F9B0",
 -3412 => x"C0C0C0BFB099F9A4",
 -3411 => x"C0C0C0BFB099F9F9",
 -3410 => x"C0C0C0BFB099F9C0",
 -3409 => x"C0C0C0BFB099C090",
 -3408 => x"C0C0C0BFB099C080",
 -3407 => x"C0C0C0BFB099C0F8",
 -3406 => x"C0C0C0BFB099C082",
 -3405 => x"C0C0C0BFB099C092",
 -3404 => x"C0C0C0BFB099C099",
 -3403 => x"C0C0C0BFB099C0B0",
 -3402 => x"C0C0C0BFB099C0A4",
 -3401 => x"C0C0C0BFB099C0F9",
 -3400 => x"C0C0C0BFB099C0C0",
 -3399 => x"C0C0C0BFB0B09090",
 -3398 => x"C0C0C0BFB0B09080",
 -3397 => x"C0C0C0BFB0B090F8",
 -3396 => x"C0C0C0BFB0B09082",
 -3395 => x"C0C0C0BFB0B09092",
 -3394 => x"C0C0C0BFB0B09099",
 -3393 => x"C0C0C0BFB0B090B0",
 -3392 => x"C0C0C0BFB0B090A4",
 -3391 => x"C0C0C0BFB0B090F9",
 -3390 => x"C0C0C0BFB0B090C0",
 -3389 => x"C0C0C0BFB0B08090",
 -3388 => x"C0C0C0BFB0B08080",
 -3387 => x"C0C0C0BFB0B080F8",
 -3386 => x"C0C0C0BFB0B08082",
 -3385 => x"C0C0C0BFB0B08092",
 -3384 => x"C0C0C0BFB0B08099",
 -3383 => x"C0C0C0BFB0B080B0",
 -3382 => x"C0C0C0BFB0B080A4",
 -3381 => x"C0C0C0BFB0B080F9",
 -3380 => x"C0C0C0BFB0B080C0",
 -3379 => x"C0C0C0BFB0B0F890",
 -3378 => x"C0C0C0BFB0B0F880",
 -3377 => x"C0C0C0BFB0B0F8F8",
 -3376 => x"C0C0C0BFB0B0F882",
 -3375 => x"C0C0C0BFB0B0F892",
 -3374 => x"C0C0C0BFB0B0F899",
 -3373 => x"C0C0C0BFB0B0F8B0",
 -3372 => x"C0C0C0BFB0B0F8A4",
 -3371 => x"C0C0C0BFB0B0F8F9",
 -3370 => x"C0C0C0BFB0B0F8C0",
 -3369 => x"C0C0C0BFB0B08290",
 -3368 => x"C0C0C0BFB0B08280",
 -3367 => x"C0C0C0BFB0B082F8",
 -3366 => x"C0C0C0BFB0B08282",
 -3365 => x"C0C0C0BFB0B08292",
 -3364 => x"C0C0C0BFB0B08299",
 -3363 => x"C0C0C0BFB0B082B0",
 -3362 => x"C0C0C0BFB0B082A4",
 -3361 => x"C0C0C0BFB0B082F9",
 -3360 => x"C0C0C0BFB0B082C0",
 -3359 => x"C0C0C0BFB0B09290",
 -3358 => x"C0C0C0BFB0B09280",
 -3357 => x"C0C0C0BFB0B092F8",
 -3356 => x"C0C0C0BFB0B09282",
 -3355 => x"C0C0C0BFB0B09292",
 -3354 => x"C0C0C0BFB0B09299",
 -3353 => x"C0C0C0BFB0B092B0",
 -3352 => x"C0C0C0BFB0B092A4",
 -3351 => x"C0C0C0BFB0B092F9",
 -3350 => x"C0C0C0BFB0B092C0",
 -3349 => x"C0C0C0BFB0B09990",
 -3348 => x"C0C0C0BFB0B09980",
 -3347 => x"C0C0C0BFB0B099F8",
 -3346 => x"C0C0C0BFB0B09982",
 -3345 => x"C0C0C0BFB0B09992",
 -3344 => x"C0C0C0BFB0B09999",
 -3343 => x"C0C0C0BFB0B099B0",
 -3342 => x"C0C0C0BFB0B099A4",
 -3341 => x"C0C0C0BFB0B099F9",
 -3340 => x"C0C0C0BFB0B099C0",
 -3339 => x"C0C0C0BFB0B0B090",
 -3338 => x"C0C0C0BFB0B0B080",
 -3337 => x"C0C0C0BFB0B0B0F8",
 -3336 => x"C0C0C0BFB0B0B082",
 -3335 => x"C0C0C0BFB0B0B092",
 -3334 => x"C0C0C0BFB0B0B099",
 -3333 => x"C0C0C0BFB0B0B0B0",
 -3332 => x"C0C0C0BFB0B0B0A4",
 -3331 => x"C0C0C0BFB0B0B0F9",
 -3330 => x"C0C0C0BFB0B0B0C0",
 -3329 => x"C0C0C0BFB0B0A490",
 -3328 => x"C0C0C0BFB0B0A480",
 -3327 => x"C0C0C0BFB0B0A4F8",
 -3326 => x"C0C0C0BFB0B0A482",
 -3325 => x"C0C0C0BFB0B0A492",
 -3324 => x"C0C0C0BFB0B0A499",
 -3323 => x"C0C0C0BFB0B0A4B0",
 -3322 => x"C0C0C0BFB0B0A4A4",
 -3321 => x"C0C0C0BFB0B0A4F9",
 -3320 => x"C0C0C0BFB0B0A4C0",
 -3319 => x"C0C0C0BFB0B0F990",
 -3318 => x"C0C0C0BFB0B0F980",
 -3317 => x"C0C0C0BFB0B0F9F8",
 -3316 => x"C0C0C0BFB0B0F982",
 -3315 => x"C0C0C0BFB0B0F992",
 -3314 => x"C0C0C0BFB0B0F999",
 -3313 => x"C0C0C0BFB0B0F9B0",
 -3312 => x"C0C0C0BFB0B0F9A4",
 -3311 => x"C0C0C0BFB0B0F9F9",
 -3310 => x"C0C0C0BFB0B0F9C0",
 -3309 => x"C0C0C0BFB0B0C090",
 -3308 => x"C0C0C0BFB0B0C080",
 -3307 => x"C0C0C0BFB0B0C0F8",
 -3306 => x"C0C0C0BFB0B0C082",
 -3305 => x"C0C0C0BFB0B0C092",
 -3304 => x"C0C0C0BFB0B0C099",
 -3303 => x"C0C0C0BFB0B0C0B0",
 -3302 => x"C0C0C0BFB0B0C0A4",
 -3301 => x"C0C0C0BFB0B0C0F9",
 -3300 => x"C0C0C0BFB0B0C0C0",
 -3299 => x"C0C0C0BFB0A49090",
 -3298 => x"C0C0C0BFB0A49080",
 -3297 => x"C0C0C0BFB0A490F8",
 -3296 => x"C0C0C0BFB0A49082",
 -3295 => x"C0C0C0BFB0A49092",
 -3294 => x"C0C0C0BFB0A49099",
 -3293 => x"C0C0C0BFB0A490B0",
 -3292 => x"C0C0C0BFB0A490A4",
 -3291 => x"C0C0C0BFB0A490F9",
 -3290 => x"C0C0C0BFB0A490C0",
 -3289 => x"C0C0C0BFB0A48090",
 -3288 => x"C0C0C0BFB0A48080",
 -3287 => x"C0C0C0BFB0A480F8",
 -3286 => x"C0C0C0BFB0A48082",
 -3285 => x"C0C0C0BFB0A48092",
 -3284 => x"C0C0C0BFB0A48099",
 -3283 => x"C0C0C0BFB0A480B0",
 -3282 => x"C0C0C0BFB0A480A4",
 -3281 => x"C0C0C0BFB0A480F9",
 -3280 => x"C0C0C0BFB0A480C0",
 -3279 => x"C0C0C0BFB0A4F890",
 -3278 => x"C0C0C0BFB0A4F880",
 -3277 => x"C0C0C0BFB0A4F8F8",
 -3276 => x"C0C0C0BFB0A4F882",
 -3275 => x"C0C0C0BFB0A4F892",
 -3274 => x"C0C0C0BFB0A4F899",
 -3273 => x"C0C0C0BFB0A4F8B0",
 -3272 => x"C0C0C0BFB0A4F8A4",
 -3271 => x"C0C0C0BFB0A4F8F9",
 -3270 => x"C0C0C0BFB0A4F8C0",
 -3269 => x"C0C0C0BFB0A48290",
 -3268 => x"C0C0C0BFB0A48280",
 -3267 => x"C0C0C0BFB0A482F8",
 -3266 => x"C0C0C0BFB0A48282",
 -3265 => x"C0C0C0BFB0A48292",
 -3264 => x"C0C0C0BFB0A48299",
 -3263 => x"C0C0C0BFB0A482B0",
 -3262 => x"C0C0C0BFB0A482A4",
 -3261 => x"C0C0C0BFB0A482F9",
 -3260 => x"C0C0C0BFB0A482C0",
 -3259 => x"C0C0C0BFB0A49290",
 -3258 => x"C0C0C0BFB0A49280",
 -3257 => x"C0C0C0BFB0A492F8",
 -3256 => x"C0C0C0BFB0A49282",
 -3255 => x"C0C0C0BFB0A49292",
 -3254 => x"C0C0C0BFB0A49299",
 -3253 => x"C0C0C0BFB0A492B0",
 -3252 => x"C0C0C0BFB0A492A4",
 -3251 => x"C0C0C0BFB0A492F9",
 -3250 => x"C0C0C0BFB0A492C0",
 -3249 => x"C0C0C0BFB0A49990",
 -3248 => x"C0C0C0BFB0A49980",
 -3247 => x"C0C0C0BFB0A499F8",
 -3246 => x"C0C0C0BFB0A49982",
 -3245 => x"C0C0C0BFB0A49992",
 -3244 => x"C0C0C0BFB0A49999",
 -3243 => x"C0C0C0BFB0A499B0",
 -3242 => x"C0C0C0BFB0A499A4",
 -3241 => x"C0C0C0BFB0A499F9",
 -3240 => x"C0C0C0BFB0A499C0",
 -3239 => x"C0C0C0BFB0A4B090",
 -3238 => x"C0C0C0BFB0A4B080",
 -3237 => x"C0C0C0BFB0A4B0F8",
 -3236 => x"C0C0C0BFB0A4B082",
 -3235 => x"C0C0C0BFB0A4B092",
 -3234 => x"C0C0C0BFB0A4B099",
 -3233 => x"C0C0C0BFB0A4B0B0",
 -3232 => x"C0C0C0BFB0A4B0A4",
 -3231 => x"C0C0C0BFB0A4B0F9",
 -3230 => x"C0C0C0BFB0A4B0C0",
 -3229 => x"C0C0C0BFB0A4A490",
 -3228 => x"C0C0C0BFB0A4A480",
 -3227 => x"C0C0C0BFB0A4A4F8",
 -3226 => x"C0C0C0BFB0A4A482",
 -3225 => x"C0C0C0BFB0A4A492",
 -3224 => x"C0C0C0BFB0A4A499",
 -3223 => x"C0C0C0BFB0A4A4B0",
 -3222 => x"C0C0C0BFB0A4A4A4",
 -3221 => x"C0C0C0BFB0A4A4F9",
 -3220 => x"C0C0C0BFB0A4A4C0",
 -3219 => x"C0C0C0BFB0A4F990",
 -3218 => x"C0C0C0BFB0A4F980",
 -3217 => x"C0C0C0BFB0A4F9F8",
 -3216 => x"C0C0C0BFB0A4F982",
 -3215 => x"C0C0C0BFB0A4F992",
 -3214 => x"C0C0C0BFB0A4F999",
 -3213 => x"C0C0C0BFB0A4F9B0",
 -3212 => x"C0C0C0BFB0A4F9A4",
 -3211 => x"C0C0C0BFB0A4F9F9",
 -3210 => x"C0C0C0BFB0A4F9C0",
 -3209 => x"C0C0C0BFB0A4C090",
 -3208 => x"C0C0C0BFB0A4C080",
 -3207 => x"C0C0C0BFB0A4C0F8",
 -3206 => x"C0C0C0BFB0A4C082",
 -3205 => x"C0C0C0BFB0A4C092",
 -3204 => x"C0C0C0BFB0A4C099",
 -3203 => x"C0C0C0BFB0A4C0B0",
 -3202 => x"C0C0C0BFB0A4C0A4",
 -3201 => x"C0C0C0BFB0A4C0F9",
 -3200 => x"C0C0C0BFB0A4C0C0",
 -3199 => x"C0C0C0BFB0F99090",
 -3198 => x"C0C0C0BFB0F99080",
 -3197 => x"C0C0C0BFB0F990F8",
 -3196 => x"C0C0C0BFB0F99082",
 -3195 => x"C0C0C0BFB0F99092",
 -3194 => x"C0C0C0BFB0F99099",
 -3193 => x"C0C0C0BFB0F990B0",
 -3192 => x"C0C0C0BFB0F990A4",
 -3191 => x"C0C0C0BFB0F990F9",
 -3190 => x"C0C0C0BFB0F990C0",
 -3189 => x"C0C0C0BFB0F98090",
 -3188 => x"C0C0C0BFB0F98080",
 -3187 => x"C0C0C0BFB0F980F8",
 -3186 => x"C0C0C0BFB0F98082",
 -3185 => x"C0C0C0BFB0F98092",
 -3184 => x"C0C0C0BFB0F98099",
 -3183 => x"C0C0C0BFB0F980B0",
 -3182 => x"C0C0C0BFB0F980A4",
 -3181 => x"C0C0C0BFB0F980F9",
 -3180 => x"C0C0C0BFB0F980C0",
 -3179 => x"C0C0C0BFB0F9F890",
 -3178 => x"C0C0C0BFB0F9F880",
 -3177 => x"C0C0C0BFB0F9F8F8",
 -3176 => x"C0C0C0BFB0F9F882",
 -3175 => x"C0C0C0BFB0F9F892",
 -3174 => x"C0C0C0BFB0F9F899",
 -3173 => x"C0C0C0BFB0F9F8B0",
 -3172 => x"C0C0C0BFB0F9F8A4",
 -3171 => x"C0C0C0BFB0F9F8F9",
 -3170 => x"C0C0C0BFB0F9F8C0",
 -3169 => x"C0C0C0BFB0F98290",
 -3168 => x"C0C0C0BFB0F98280",
 -3167 => x"C0C0C0BFB0F982F8",
 -3166 => x"C0C0C0BFB0F98282",
 -3165 => x"C0C0C0BFB0F98292",
 -3164 => x"C0C0C0BFB0F98299",
 -3163 => x"C0C0C0BFB0F982B0",
 -3162 => x"C0C0C0BFB0F982A4",
 -3161 => x"C0C0C0BFB0F982F9",
 -3160 => x"C0C0C0BFB0F982C0",
 -3159 => x"C0C0C0BFB0F99290",
 -3158 => x"C0C0C0BFB0F99280",
 -3157 => x"C0C0C0BFB0F992F8",
 -3156 => x"C0C0C0BFB0F99282",
 -3155 => x"C0C0C0BFB0F99292",
 -3154 => x"C0C0C0BFB0F99299",
 -3153 => x"C0C0C0BFB0F992B0",
 -3152 => x"C0C0C0BFB0F992A4",
 -3151 => x"C0C0C0BFB0F992F9",
 -3150 => x"C0C0C0BFB0F992C0",
 -3149 => x"C0C0C0BFB0F99990",
 -3148 => x"C0C0C0BFB0F99980",
 -3147 => x"C0C0C0BFB0F999F8",
 -3146 => x"C0C0C0BFB0F99982",
 -3145 => x"C0C0C0BFB0F99992",
 -3144 => x"C0C0C0BFB0F99999",
 -3143 => x"C0C0C0BFB0F999B0",
 -3142 => x"C0C0C0BFB0F999A4",
 -3141 => x"C0C0C0BFB0F999F9",
 -3140 => x"C0C0C0BFB0F999C0",
 -3139 => x"C0C0C0BFB0F9B090",
 -3138 => x"C0C0C0BFB0F9B080",
 -3137 => x"C0C0C0BFB0F9B0F8",
 -3136 => x"C0C0C0BFB0F9B082",
 -3135 => x"C0C0C0BFB0F9B092",
 -3134 => x"C0C0C0BFB0F9B099",
 -3133 => x"C0C0C0BFB0F9B0B0",
 -3132 => x"C0C0C0BFB0F9B0A4",
 -3131 => x"C0C0C0BFB0F9B0F9",
 -3130 => x"C0C0C0BFB0F9B0C0",
 -3129 => x"C0C0C0BFB0F9A490",
 -3128 => x"C0C0C0BFB0F9A480",
 -3127 => x"C0C0C0BFB0F9A4F8",
 -3126 => x"C0C0C0BFB0F9A482",
 -3125 => x"C0C0C0BFB0F9A492",
 -3124 => x"C0C0C0BFB0F9A499",
 -3123 => x"C0C0C0BFB0F9A4B0",
 -3122 => x"C0C0C0BFB0F9A4A4",
 -3121 => x"C0C0C0BFB0F9A4F9",
 -3120 => x"C0C0C0BFB0F9A4C0",
 -3119 => x"C0C0C0BFB0F9F990",
 -3118 => x"C0C0C0BFB0F9F980",
 -3117 => x"C0C0C0BFB0F9F9F8",
 -3116 => x"C0C0C0BFB0F9F982",
 -3115 => x"C0C0C0BFB0F9F992",
 -3114 => x"C0C0C0BFB0F9F999",
 -3113 => x"C0C0C0BFB0F9F9B0",
 -3112 => x"C0C0C0BFB0F9F9A4",
 -3111 => x"C0C0C0BFB0F9F9F9",
 -3110 => x"C0C0C0BFB0F9F9C0",
 -3109 => x"C0C0C0BFB0F9C090",
 -3108 => x"C0C0C0BFB0F9C080",
 -3107 => x"C0C0C0BFB0F9C0F8",
 -3106 => x"C0C0C0BFB0F9C082",
 -3105 => x"C0C0C0BFB0F9C092",
 -3104 => x"C0C0C0BFB0F9C099",
 -3103 => x"C0C0C0BFB0F9C0B0",
 -3102 => x"C0C0C0BFB0F9C0A4",
 -3101 => x"C0C0C0BFB0F9C0F9",
 -3100 => x"C0C0C0BFB0F9C0C0",
 -3099 => x"C0C0C0BFB0C09090",
 -3098 => x"C0C0C0BFB0C09080",
 -3097 => x"C0C0C0BFB0C090F8",
 -3096 => x"C0C0C0BFB0C09082",
 -3095 => x"C0C0C0BFB0C09092",
 -3094 => x"C0C0C0BFB0C09099",
 -3093 => x"C0C0C0BFB0C090B0",
 -3092 => x"C0C0C0BFB0C090A4",
 -3091 => x"C0C0C0BFB0C090F9",
 -3090 => x"C0C0C0BFB0C090C0",
 -3089 => x"C0C0C0BFB0C08090",
 -3088 => x"C0C0C0BFB0C08080",
 -3087 => x"C0C0C0BFB0C080F8",
 -3086 => x"C0C0C0BFB0C08082",
 -3085 => x"C0C0C0BFB0C08092",
 -3084 => x"C0C0C0BFB0C08099",
 -3083 => x"C0C0C0BFB0C080B0",
 -3082 => x"C0C0C0BFB0C080A4",
 -3081 => x"C0C0C0BFB0C080F9",
 -3080 => x"C0C0C0BFB0C080C0",
 -3079 => x"C0C0C0BFB0C0F890",
 -3078 => x"C0C0C0BFB0C0F880",
 -3077 => x"C0C0C0BFB0C0F8F8",
 -3076 => x"C0C0C0BFB0C0F882",
 -3075 => x"C0C0C0BFB0C0F892",
 -3074 => x"C0C0C0BFB0C0F899",
 -3073 => x"C0C0C0BFB0C0F8B0",
 -3072 => x"C0C0C0BFB0C0F8A4",
 -3071 => x"C0C0C0BFB0C0F8F9",
 -3070 => x"C0C0C0BFB0C0F8C0",
 -3069 => x"C0C0C0BFB0C08290",
 -3068 => x"C0C0C0BFB0C08280",
 -3067 => x"C0C0C0BFB0C082F8",
 -3066 => x"C0C0C0BFB0C08282",
 -3065 => x"C0C0C0BFB0C08292",
 -3064 => x"C0C0C0BFB0C08299",
 -3063 => x"C0C0C0BFB0C082B0",
 -3062 => x"C0C0C0BFB0C082A4",
 -3061 => x"C0C0C0BFB0C082F9",
 -3060 => x"C0C0C0BFB0C082C0",
 -3059 => x"C0C0C0BFB0C09290",
 -3058 => x"C0C0C0BFB0C09280",
 -3057 => x"C0C0C0BFB0C092F8",
 -3056 => x"C0C0C0BFB0C09282",
 -3055 => x"C0C0C0BFB0C09292",
 -3054 => x"C0C0C0BFB0C09299",
 -3053 => x"C0C0C0BFB0C092B0",
 -3052 => x"C0C0C0BFB0C092A4",
 -3051 => x"C0C0C0BFB0C092F9",
 -3050 => x"C0C0C0BFB0C092C0",
 -3049 => x"C0C0C0BFB0C09990",
 -3048 => x"C0C0C0BFB0C09980",
 -3047 => x"C0C0C0BFB0C099F8",
 -3046 => x"C0C0C0BFB0C09982",
 -3045 => x"C0C0C0BFB0C09992",
 -3044 => x"C0C0C0BFB0C09999",
 -3043 => x"C0C0C0BFB0C099B0",
 -3042 => x"C0C0C0BFB0C099A4",
 -3041 => x"C0C0C0BFB0C099F9",
 -3040 => x"C0C0C0BFB0C099C0",
 -3039 => x"C0C0C0BFB0C0B090",
 -3038 => x"C0C0C0BFB0C0B080",
 -3037 => x"C0C0C0BFB0C0B0F8",
 -3036 => x"C0C0C0BFB0C0B082",
 -3035 => x"C0C0C0BFB0C0B092",
 -3034 => x"C0C0C0BFB0C0B099",
 -3033 => x"C0C0C0BFB0C0B0B0",
 -3032 => x"C0C0C0BFB0C0B0A4",
 -3031 => x"C0C0C0BFB0C0B0F9",
 -3030 => x"C0C0C0BFB0C0B0C0",
 -3029 => x"C0C0C0BFB0C0A490",
 -3028 => x"C0C0C0BFB0C0A480",
 -3027 => x"C0C0C0BFB0C0A4F8",
 -3026 => x"C0C0C0BFB0C0A482",
 -3025 => x"C0C0C0BFB0C0A492",
 -3024 => x"C0C0C0BFB0C0A499",
 -3023 => x"C0C0C0BFB0C0A4B0",
 -3022 => x"C0C0C0BFB0C0A4A4",
 -3021 => x"C0C0C0BFB0C0A4F9",
 -3020 => x"C0C0C0BFB0C0A4C0",
 -3019 => x"C0C0C0BFB0C0F990",
 -3018 => x"C0C0C0BFB0C0F980",
 -3017 => x"C0C0C0BFB0C0F9F8",
 -3016 => x"C0C0C0BFB0C0F982",
 -3015 => x"C0C0C0BFB0C0F992",
 -3014 => x"C0C0C0BFB0C0F999",
 -3013 => x"C0C0C0BFB0C0F9B0",
 -3012 => x"C0C0C0BFB0C0F9A4",
 -3011 => x"C0C0C0BFB0C0F9F9",
 -3010 => x"C0C0C0BFB0C0F9C0",
 -3009 => x"C0C0C0BFB0C0C090",
 -3008 => x"C0C0C0BFB0C0C080",
 -3007 => x"C0C0C0BFB0C0C0F8",
 -3006 => x"C0C0C0BFB0C0C082",
 -3005 => x"C0C0C0BFB0C0C092",
 -3004 => x"C0C0C0BFB0C0C099",
 -3003 => x"C0C0C0BFB0C0C0B0",
 -3002 => x"C0C0C0BFB0C0C0A4",
 -3001 => x"C0C0C0BFB0C0C0F9",
 -3000 => x"C0C0C0BFB0C0C0C0",
 -2999 => x"C0C0C0BFA4909090",
 -2998 => x"C0C0C0BFA4909080",
 -2997 => x"C0C0C0BFA49090F8",
 -2996 => x"C0C0C0BFA4909082",
 -2995 => x"C0C0C0BFA4909092",
 -2994 => x"C0C0C0BFA4909099",
 -2993 => x"C0C0C0BFA49090B0",
 -2992 => x"C0C0C0BFA49090A4",
 -2991 => x"C0C0C0BFA49090F9",
 -2990 => x"C0C0C0BFA49090C0",
 -2989 => x"C0C0C0BFA4908090",
 -2988 => x"C0C0C0BFA4908080",
 -2987 => x"C0C0C0BFA49080F8",
 -2986 => x"C0C0C0BFA4908082",
 -2985 => x"C0C0C0BFA4908092",
 -2984 => x"C0C0C0BFA4908099",
 -2983 => x"C0C0C0BFA49080B0",
 -2982 => x"C0C0C0BFA49080A4",
 -2981 => x"C0C0C0BFA49080F9",
 -2980 => x"C0C0C0BFA49080C0",
 -2979 => x"C0C0C0BFA490F890",
 -2978 => x"C0C0C0BFA490F880",
 -2977 => x"C0C0C0BFA490F8F8",
 -2976 => x"C0C0C0BFA490F882",
 -2975 => x"C0C0C0BFA490F892",
 -2974 => x"C0C0C0BFA490F899",
 -2973 => x"C0C0C0BFA490F8B0",
 -2972 => x"C0C0C0BFA490F8A4",
 -2971 => x"C0C0C0BFA490F8F9",
 -2970 => x"C0C0C0BFA490F8C0",
 -2969 => x"C0C0C0BFA4908290",
 -2968 => x"C0C0C0BFA4908280",
 -2967 => x"C0C0C0BFA49082F8",
 -2966 => x"C0C0C0BFA4908282",
 -2965 => x"C0C0C0BFA4908292",
 -2964 => x"C0C0C0BFA4908299",
 -2963 => x"C0C0C0BFA49082B0",
 -2962 => x"C0C0C0BFA49082A4",
 -2961 => x"C0C0C0BFA49082F9",
 -2960 => x"C0C0C0BFA49082C0",
 -2959 => x"C0C0C0BFA4909290",
 -2958 => x"C0C0C0BFA4909280",
 -2957 => x"C0C0C0BFA49092F8",
 -2956 => x"C0C0C0BFA4909282",
 -2955 => x"C0C0C0BFA4909292",
 -2954 => x"C0C0C0BFA4909299",
 -2953 => x"C0C0C0BFA49092B0",
 -2952 => x"C0C0C0BFA49092A4",
 -2951 => x"C0C0C0BFA49092F9",
 -2950 => x"C0C0C0BFA49092C0",
 -2949 => x"C0C0C0BFA4909990",
 -2948 => x"C0C0C0BFA4909980",
 -2947 => x"C0C0C0BFA49099F8",
 -2946 => x"C0C0C0BFA4909982",
 -2945 => x"C0C0C0BFA4909992",
 -2944 => x"C0C0C0BFA4909999",
 -2943 => x"C0C0C0BFA49099B0",
 -2942 => x"C0C0C0BFA49099A4",
 -2941 => x"C0C0C0BFA49099F9",
 -2940 => x"C0C0C0BFA49099C0",
 -2939 => x"C0C0C0BFA490B090",
 -2938 => x"C0C0C0BFA490B080",
 -2937 => x"C0C0C0BFA490B0F8",
 -2936 => x"C0C0C0BFA490B082",
 -2935 => x"C0C0C0BFA490B092",
 -2934 => x"C0C0C0BFA490B099",
 -2933 => x"C0C0C0BFA490B0B0",
 -2932 => x"C0C0C0BFA490B0A4",
 -2931 => x"C0C0C0BFA490B0F9",
 -2930 => x"C0C0C0BFA490B0C0",
 -2929 => x"C0C0C0BFA490A490",
 -2928 => x"C0C0C0BFA490A480",
 -2927 => x"C0C0C0BFA490A4F8",
 -2926 => x"C0C0C0BFA490A482",
 -2925 => x"C0C0C0BFA490A492",
 -2924 => x"C0C0C0BFA490A499",
 -2923 => x"C0C0C0BFA490A4B0",
 -2922 => x"C0C0C0BFA490A4A4",
 -2921 => x"C0C0C0BFA490A4F9",
 -2920 => x"C0C0C0BFA490A4C0",
 -2919 => x"C0C0C0BFA490F990",
 -2918 => x"C0C0C0BFA490F980",
 -2917 => x"C0C0C0BFA490F9F8",
 -2916 => x"C0C0C0BFA490F982",
 -2915 => x"C0C0C0BFA490F992",
 -2914 => x"C0C0C0BFA490F999",
 -2913 => x"C0C0C0BFA490F9B0",
 -2912 => x"C0C0C0BFA490F9A4",
 -2911 => x"C0C0C0BFA490F9F9",
 -2910 => x"C0C0C0BFA490F9C0",
 -2909 => x"C0C0C0BFA490C090",
 -2908 => x"C0C0C0BFA490C080",
 -2907 => x"C0C0C0BFA490C0F8",
 -2906 => x"C0C0C0BFA490C082",
 -2905 => x"C0C0C0BFA490C092",
 -2904 => x"C0C0C0BFA490C099",
 -2903 => x"C0C0C0BFA490C0B0",
 -2902 => x"C0C0C0BFA490C0A4",
 -2901 => x"C0C0C0BFA490C0F9",
 -2900 => x"C0C0C0BFA490C0C0",
 -2899 => x"C0C0C0BFA4809090",
 -2898 => x"C0C0C0BFA4809080",
 -2897 => x"C0C0C0BFA48090F8",
 -2896 => x"C0C0C0BFA4809082",
 -2895 => x"C0C0C0BFA4809092",
 -2894 => x"C0C0C0BFA4809099",
 -2893 => x"C0C0C0BFA48090B0",
 -2892 => x"C0C0C0BFA48090A4",
 -2891 => x"C0C0C0BFA48090F9",
 -2890 => x"C0C0C0BFA48090C0",
 -2889 => x"C0C0C0BFA4808090",
 -2888 => x"C0C0C0BFA4808080",
 -2887 => x"C0C0C0BFA48080F8",
 -2886 => x"C0C0C0BFA4808082",
 -2885 => x"C0C0C0BFA4808092",
 -2884 => x"C0C0C0BFA4808099",
 -2883 => x"C0C0C0BFA48080B0",
 -2882 => x"C0C0C0BFA48080A4",
 -2881 => x"C0C0C0BFA48080F9",
 -2880 => x"C0C0C0BFA48080C0",
 -2879 => x"C0C0C0BFA480F890",
 -2878 => x"C0C0C0BFA480F880",
 -2877 => x"C0C0C0BFA480F8F8",
 -2876 => x"C0C0C0BFA480F882",
 -2875 => x"C0C0C0BFA480F892",
 -2874 => x"C0C0C0BFA480F899",
 -2873 => x"C0C0C0BFA480F8B0",
 -2872 => x"C0C0C0BFA480F8A4",
 -2871 => x"C0C0C0BFA480F8F9",
 -2870 => x"C0C0C0BFA480F8C0",
 -2869 => x"C0C0C0BFA4808290",
 -2868 => x"C0C0C0BFA4808280",
 -2867 => x"C0C0C0BFA48082F8",
 -2866 => x"C0C0C0BFA4808282",
 -2865 => x"C0C0C0BFA4808292",
 -2864 => x"C0C0C0BFA4808299",
 -2863 => x"C0C0C0BFA48082B0",
 -2862 => x"C0C0C0BFA48082A4",
 -2861 => x"C0C0C0BFA48082F9",
 -2860 => x"C0C0C0BFA48082C0",
 -2859 => x"C0C0C0BFA4809290",
 -2858 => x"C0C0C0BFA4809280",
 -2857 => x"C0C0C0BFA48092F8",
 -2856 => x"C0C0C0BFA4809282",
 -2855 => x"C0C0C0BFA4809292",
 -2854 => x"C0C0C0BFA4809299",
 -2853 => x"C0C0C0BFA48092B0",
 -2852 => x"C0C0C0BFA48092A4",
 -2851 => x"C0C0C0BFA48092F9",
 -2850 => x"C0C0C0BFA48092C0",
 -2849 => x"C0C0C0BFA4809990",
 -2848 => x"C0C0C0BFA4809980",
 -2847 => x"C0C0C0BFA48099F8",
 -2846 => x"C0C0C0BFA4809982",
 -2845 => x"C0C0C0BFA4809992",
 -2844 => x"C0C0C0BFA4809999",
 -2843 => x"C0C0C0BFA48099B0",
 -2842 => x"C0C0C0BFA48099A4",
 -2841 => x"C0C0C0BFA48099F9",
 -2840 => x"C0C0C0BFA48099C0",
 -2839 => x"C0C0C0BFA480B090",
 -2838 => x"C0C0C0BFA480B080",
 -2837 => x"C0C0C0BFA480B0F8",
 -2836 => x"C0C0C0BFA480B082",
 -2835 => x"C0C0C0BFA480B092",
 -2834 => x"C0C0C0BFA480B099",
 -2833 => x"C0C0C0BFA480B0B0",
 -2832 => x"C0C0C0BFA480B0A4",
 -2831 => x"C0C0C0BFA480B0F9",
 -2830 => x"C0C0C0BFA480B0C0",
 -2829 => x"C0C0C0BFA480A490",
 -2828 => x"C0C0C0BFA480A480",
 -2827 => x"C0C0C0BFA480A4F8",
 -2826 => x"C0C0C0BFA480A482",
 -2825 => x"C0C0C0BFA480A492",
 -2824 => x"C0C0C0BFA480A499",
 -2823 => x"C0C0C0BFA480A4B0",
 -2822 => x"C0C0C0BFA480A4A4",
 -2821 => x"C0C0C0BFA480A4F9",
 -2820 => x"C0C0C0BFA480A4C0",
 -2819 => x"C0C0C0BFA480F990",
 -2818 => x"C0C0C0BFA480F980",
 -2817 => x"C0C0C0BFA480F9F8",
 -2816 => x"C0C0C0BFA480F982",
 -2815 => x"C0C0C0BFA480F992",
 -2814 => x"C0C0C0BFA480F999",
 -2813 => x"C0C0C0BFA480F9B0",
 -2812 => x"C0C0C0BFA480F9A4",
 -2811 => x"C0C0C0BFA480F9F9",
 -2810 => x"C0C0C0BFA480F9C0",
 -2809 => x"C0C0C0BFA480C090",
 -2808 => x"C0C0C0BFA480C080",
 -2807 => x"C0C0C0BFA480C0F8",
 -2806 => x"C0C0C0BFA480C082",
 -2805 => x"C0C0C0BFA480C092",
 -2804 => x"C0C0C0BFA480C099",
 -2803 => x"C0C0C0BFA480C0B0",
 -2802 => x"C0C0C0BFA480C0A4",
 -2801 => x"C0C0C0BFA480C0F9",
 -2800 => x"C0C0C0BFA480C0C0",
 -2799 => x"C0C0C0BFA4F89090",
 -2798 => x"C0C0C0BFA4F89080",
 -2797 => x"C0C0C0BFA4F890F8",
 -2796 => x"C0C0C0BFA4F89082",
 -2795 => x"C0C0C0BFA4F89092",
 -2794 => x"C0C0C0BFA4F89099",
 -2793 => x"C0C0C0BFA4F890B0",
 -2792 => x"C0C0C0BFA4F890A4",
 -2791 => x"C0C0C0BFA4F890F9",
 -2790 => x"C0C0C0BFA4F890C0",
 -2789 => x"C0C0C0BFA4F88090",
 -2788 => x"C0C0C0BFA4F88080",
 -2787 => x"C0C0C0BFA4F880F8",
 -2786 => x"C0C0C0BFA4F88082",
 -2785 => x"C0C0C0BFA4F88092",
 -2784 => x"C0C0C0BFA4F88099",
 -2783 => x"C0C0C0BFA4F880B0",
 -2782 => x"C0C0C0BFA4F880A4",
 -2781 => x"C0C0C0BFA4F880F9",
 -2780 => x"C0C0C0BFA4F880C0",
 -2779 => x"C0C0C0BFA4F8F890",
 -2778 => x"C0C0C0BFA4F8F880",
 -2777 => x"C0C0C0BFA4F8F8F8",
 -2776 => x"C0C0C0BFA4F8F882",
 -2775 => x"C0C0C0BFA4F8F892",
 -2774 => x"C0C0C0BFA4F8F899",
 -2773 => x"C0C0C0BFA4F8F8B0",
 -2772 => x"C0C0C0BFA4F8F8A4",
 -2771 => x"C0C0C0BFA4F8F8F9",
 -2770 => x"C0C0C0BFA4F8F8C0",
 -2769 => x"C0C0C0BFA4F88290",
 -2768 => x"C0C0C0BFA4F88280",
 -2767 => x"C0C0C0BFA4F882F8",
 -2766 => x"C0C0C0BFA4F88282",
 -2765 => x"C0C0C0BFA4F88292",
 -2764 => x"C0C0C0BFA4F88299",
 -2763 => x"C0C0C0BFA4F882B0",
 -2762 => x"C0C0C0BFA4F882A4",
 -2761 => x"C0C0C0BFA4F882F9",
 -2760 => x"C0C0C0BFA4F882C0",
 -2759 => x"C0C0C0BFA4F89290",
 -2758 => x"C0C0C0BFA4F89280",
 -2757 => x"C0C0C0BFA4F892F8",
 -2756 => x"C0C0C0BFA4F89282",
 -2755 => x"C0C0C0BFA4F89292",
 -2754 => x"C0C0C0BFA4F89299",
 -2753 => x"C0C0C0BFA4F892B0",
 -2752 => x"C0C0C0BFA4F892A4",
 -2751 => x"C0C0C0BFA4F892F9",
 -2750 => x"C0C0C0BFA4F892C0",
 -2749 => x"C0C0C0BFA4F89990",
 -2748 => x"C0C0C0BFA4F89980",
 -2747 => x"C0C0C0BFA4F899F8",
 -2746 => x"C0C0C0BFA4F89982",
 -2745 => x"C0C0C0BFA4F89992",
 -2744 => x"C0C0C0BFA4F89999",
 -2743 => x"C0C0C0BFA4F899B0",
 -2742 => x"C0C0C0BFA4F899A4",
 -2741 => x"C0C0C0BFA4F899F9",
 -2740 => x"C0C0C0BFA4F899C0",
 -2739 => x"C0C0C0BFA4F8B090",
 -2738 => x"C0C0C0BFA4F8B080",
 -2737 => x"C0C0C0BFA4F8B0F8",
 -2736 => x"C0C0C0BFA4F8B082",
 -2735 => x"C0C0C0BFA4F8B092",
 -2734 => x"C0C0C0BFA4F8B099",
 -2733 => x"C0C0C0BFA4F8B0B0",
 -2732 => x"C0C0C0BFA4F8B0A4",
 -2731 => x"C0C0C0BFA4F8B0F9",
 -2730 => x"C0C0C0BFA4F8B0C0",
 -2729 => x"C0C0C0BFA4F8A490",
 -2728 => x"C0C0C0BFA4F8A480",
 -2727 => x"C0C0C0BFA4F8A4F8",
 -2726 => x"C0C0C0BFA4F8A482",
 -2725 => x"C0C0C0BFA4F8A492",
 -2724 => x"C0C0C0BFA4F8A499",
 -2723 => x"C0C0C0BFA4F8A4B0",
 -2722 => x"C0C0C0BFA4F8A4A4",
 -2721 => x"C0C0C0BFA4F8A4F9",
 -2720 => x"C0C0C0BFA4F8A4C0",
 -2719 => x"C0C0C0BFA4F8F990",
 -2718 => x"C0C0C0BFA4F8F980",
 -2717 => x"C0C0C0BFA4F8F9F8",
 -2716 => x"C0C0C0BFA4F8F982",
 -2715 => x"C0C0C0BFA4F8F992",
 -2714 => x"C0C0C0BFA4F8F999",
 -2713 => x"C0C0C0BFA4F8F9B0",
 -2712 => x"C0C0C0BFA4F8F9A4",
 -2711 => x"C0C0C0BFA4F8F9F9",
 -2710 => x"C0C0C0BFA4F8F9C0",
 -2709 => x"C0C0C0BFA4F8C090",
 -2708 => x"C0C0C0BFA4F8C080",
 -2707 => x"C0C0C0BFA4F8C0F8",
 -2706 => x"C0C0C0BFA4F8C082",
 -2705 => x"C0C0C0BFA4F8C092",
 -2704 => x"C0C0C0BFA4F8C099",
 -2703 => x"C0C0C0BFA4F8C0B0",
 -2702 => x"C0C0C0BFA4F8C0A4",
 -2701 => x"C0C0C0BFA4F8C0F9",
 -2700 => x"C0C0C0BFA4F8C0C0",
 -2699 => x"C0C0C0BFA4829090",
 -2698 => x"C0C0C0BFA4829080",
 -2697 => x"C0C0C0BFA48290F8",
 -2696 => x"C0C0C0BFA4829082",
 -2695 => x"C0C0C0BFA4829092",
 -2694 => x"C0C0C0BFA4829099",
 -2693 => x"C0C0C0BFA48290B0",
 -2692 => x"C0C0C0BFA48290A4",
 -2691 => x"C0C0C0BFA48290F9",
 -2690 => x"C0C0C0BFA48290C0",
 -2689 => x"C0C0C0BFA4828090",
 -2688 => x"C0C0C0BFA4828080",
 -2687 => x"C0C0C0BFA48280F8",
 -2686 => x"C0C0C0BFA4828082",
 -2685 => x"C0C0C0BFA4828092",
 -2684 => x"C0C0C0BFA4828099",
 -2683 => x"C0C0C0BFA48280B0",
 -2682 => x"C0C0C0BFA48280A4",
 -2681 => x"C0C0C0BFA48280F9",
 -2680 => x"C0C0C0BFA48280C0",
 -2679 => x"C0C0C0BFA482F890",
 -2678 => x"C0C0C0BFA482F880",
 -2677 => x"C0C0C0BFA482F8F8",
 -2676 => x"C0C0C0BFA482F882",
 -2675 => x"C0C0C0BFA482F892",
 -2674 => x"C0C0C0BFA482F899",
 -2673 => x"C0C0C0BFA482F8B0",
 -2672 => x"C0C0C0BFA482F8A4",
 -2671 => x"C0C0C0BFA482F8F9",
 -2670 => x"C0C0C0BFA482F8C0",
 -2669 => x"C0C0C0BFA4828290",
 -2668 => x"C0C0C0BFA4828280",
 -2667 => x"C0C0C0BFA48282F8",
 -2666 => x"C0C0C0BFA4828282",
 -2665 => x"C0C0C0BFA4828292",
 -2664 => x"C0C0C0BFA4828299",
 -2663 => x"C0C0C0BFA48282B0",
 -2662 => x"C0C0C0BFA48282A4",
 -2661 => x"C0C0C0BFA48282F9",
 -2660 => x"C0C0C0BFA48282C0",
 -2659 => x"C0C0C0BFA4829290",
 -2658 => x"C0C0C0BFA4829280",
 -2657 => x"C0C0C0BFA48292F8",
 -2656 => x"C0C0C0BFA4829282",
 -2655 => x"C0C0C0BFA4829292",
 -2654 => x"C0C0C0BFA4829299",
 -2653 => x"C0C0C0BFA48292B0",
 -2652 => x"C0C0C0BFA48292A4",
 -2651 => x"C0C0C0BFA48292F9",
 -2650 => x"C0C0C0BFA48292C0",
 -2649 => x"C0C0C0BFA4829990",
 -2648 => x"C0C0C0BFA4829980",
 -2647 => x"C0C0C0BFA48299F8",
 -2646 => x"C0C0C0BFA4829982",
 -2645 => x"C0C0C0BFA4829992",
 -2644 => x"C0C0C0BFA4829999",
 -2643 => x"C0C0C0BFA48299B0",
 -2642 => x"C0C0C0BFA48299A4",
 -2641 => x"C0C0C0BFA48299F9",
 -2640 => x"C0C0C0BFA48299C0",
 -2639 => x"C0C0C0BFA482B090",
 -2638 => x"C0C0C0BFA482B080",
 -2637 => x"C0C0C0BFA482B0F8",
 -2636 => x"C0C0C0BFA482B082",
 -2635 => x"C0C0C0BFA482B092",
 -2634 => x"C0C0C0BFA482B099",
 -2633 => x"C0C0C0BFA482B0B0",
 -2632 => x"C0C0C0BFA482B0A4",
 -2631 => x"C0C0C0BFA482B0F9",
 -2630 => x"C0C0C0BFA482B0C0",
 -2629 => x"C0C0C0BFA482A490",
 -2628 => x"C0C0C0BFA482A480",
 -2627 => x"C0C0C0BFA482A4F8",
 -2626 => x"C0C0C0BFA482A482",
 -2625 => x"C0C0C0BFA482A492",
 -2624 => x"C0C0C0BFA482A499",
 -2623 => x"C0C0C0BFA482A4B0",
 -2622 => x"C0C0C0BFA482A4A4",
 -2621 => x"C0C0C0BFA482A4F9",
 -2620 => x"C0C0C0BFA482A4C0",
 -2619 => x"C0C0C0BFA482F990",
 -2618 => x"C0C0C0BFA482F980",
 -2617 => x"C0C0C0BFA482F9F8",
 -2616 => x"C0C0C0BFA482F982",
 -2615 => x"C0C0C0BFA482F992",
 -2614 => x"C0C0C0BFA482F999",
 -2613 => x"C0C0C0BFA482F9B0",
 -2612 => x"C0C0C0BFA482F9A4",
 -2611 => x"C0C0C0BFA482F9F9",
 -2610 => x"C0C0C0BFA482F9C0",
 -2609 => x"C0C0C0BFA482C090",
 -2608 => x"C0C0C0BFA482C080",
 -2607 => x"C0C0C0BFA482C0F8",
 -2606 => x"C0C0C0BFA482C082",
 -2605 => x"C0C0C0BFA482C092",
 -2604 => x"C0C0C0BFA482C099",
 -2603 => x"C0C0C0BFA482C0B0",
 -2602 => x"C0C0C0BFA482C0A4",
 -2601 => x"C0C0C0BFA482C0F9",
 -2600 => x"C0C0C0BFA482C0C0",
 -2599 => x"C0C0C0BFA4929090",
 -2598 => x"C0C0C0BFA4929080",
 -2597 => x"C0C0C0BFA49290F8",
 -2596 => x"C0C0C0BFA4929082",
 -2595 => x"C0C0C0BFA4929092",
 -2594 => x"C0C0C0BFA4929099",
 -2593 => x"C0C0C0BFA49290B0",
 -2592 => x"C0C0C0BFA49290A4",
 -2591 => x"C0C0C0BFA49290F9",
 -2590 => x"C0C0C0BFA49290C0",
 -2589 => x"C0C0C0BFA4928090",
 -2588 => x"C0C0C0BFA4928080",
 -2587 => x"C0C0C0BFA49280F8",
 -2586 => x"C0C0C0BFA4928082",
 -2585 => x"C0C0C0BFA4928092",
 -2584 => x"C0C0C0BFA4928099",
 -2583 => x"C0C0C0BFA49280B0",
 -2582 => x"C0C0C0BFA49280A4",
 -2581 => x"C0C0C0BFA49280F9",
 -2580 => x"C0C0C0BFA49280C0",
 -2579 => x"C0C0C0BFA492F890",
 -2578 => x"C0C0C0BFA492F880",
 -2577 => x"C0C0C0BFA492F8F8",
 -2576 => x"C0C0C0BFA492F882",
 -2575 => x"C0C0C0BFA492F892",
 -2574 => x"C0C0C0BFA492F899",
 -2573 => x"C0C0C0BFA492F8B0",
 -2572 => x"C0C0C0BFA492F8A4",
 -2571 => x"C0C0C0BFA492F8F9",
 -2570 => x"C0C0C0BFA492F8C0",
 -2569 => x"C0C0C0BFA4928290",
 -2568 => x"C0C0C0BFA4928280",
 -2567 => x"C0C0C0BFA49282F8",
 -2566 => x"C0C0C0BFA4928282",
 -2565 => x"C0C0C0BFA4928292",
 -2564 => x"C0C0C0BFA4928299",
 -2563 => x"C0C0C0BFA49282B0",
 -2562 => x"C0C0C0BFA49282A4",
 -2561 => x"C0C0C0BFA49282F9",
 -2560 => x"C0C0C0BFA49282C0",
 -2559 => x"C0C0C0BFA4929290",
 -2558 => x"C0C0C0BFA4929280",
 -2557 => x"C0C0C0BFA49292F8",
 -2556 => x"C0C0C0BFA4929282",
 -2555 => x"C0C0C0BFA4929292",
 -2554 => x"C0C0C0BFA4929299",
 -2553 => x"C0C0C0BFA49292B0",
 -2552 => x"C0C0C0BFA49292A4",
 -2551 => x"C0C0C0BFA49292F9",
 -2550 => x"C0C0C0BFA49292C0",
 -2549 => x"C0C0C0BFA4929990",
 -2548 => x"C0C0C0BFA4929980",
 -2547 => x"C0C0C0BFA49299F8",
 -2546 => x"C0C0C0BFA4929982",
 -2545 => x"C0C0C0BFA4929992",
 -2544 => x"C0C0C0BFA4929999",
 -2543 => x"C0C0C0BFA49299B0",
 -2542 => x"C0C0C0BFA49299A4",
 -2541 => x"C0C0C0BFA49299F9",
 -2540 => x"C0C0C0BFA49299C0",
 -2539 => x"C0C0C0BFA492B090",
 -2538 => x"C0C0C0BFA492B080",
 -2537 => x"C0C0C0BFA492B0F8",
 -2536 => x"C0C0C0BFA492B082",
 -2535 => x"C0C0C0BFA492B092",
 -2534 => x"C0C0C0BFA492B099",
 -2533 => x"C0C0C0BFA492B0B0",
 -2532 => x"C0C0C0BFA492B0A4",
 -2531 => x"C0C0C0BFA492B0F9",
 -2530 => x"C0C0C0BFA492B0C0",
 -2529 => x"C0C0C0BFA492A490",
 -2528 => x"C0C0C0BFA492A480",
 -2527 => x"C0C0C0BFA492A4F8",
 -2526 => x"C0C0C0BFA492A482",
 -2525 => x"C0C0C0BFA492A492",
 -2524 => x"C0C0C0BFA492A499",
 -2523 => x"C0C0C0BFA492A4B0",
 -2522 => x"C0C0C0BFA492A4A4",
 -2521 => x"C0C0C0BFA492A4F9",
 -2520 => x"C0C0C0BFA492A4C0",
 -2519 => x"C0C0C0BFA492F990",
 -2518 => x"C0C0C0BFA492F980",
 -2517 => x"C0C0C0BFA492F9F8",
 -2516 => x"C0C0C0BFA492F982",
 -2515 => x"C0C0C0BFA492F992",
 -2514 => x"C0C0C0BFA492F999",
 -2513 => x"C0C0C0BFA492F9B0",
 -2512 => x"C0C0C0BFA492F9A4",
 -2511 => x"C0C0C0BFA492F9F9",
 -2510 => x"C0C0C0BFA492F9C0",
 -2509 => x"C0C0C0BFA492C090",
 -2508 => x"C0C0C0BFA492C080",
 -2507 => x"C0C0C0BFA492C0F8",
 -2506 => x"C0C0C0BFA492C082",
 -2505 => x"C0C0C0BFA492C092",
 -2504 => x"C0C0C0BFA492C099",
 -2503 => x"C0C0C0BFA492C0B0",
 -2502 => x"C0C0C0BFA492C0A4",
 -2501 => x"C0C0C0BFA492C0F9",
 -2500 => x"C0C0C0BFA492C0C0",
 -2499 => x"C0C0C0BFA4999090",
 -2498 => x"C0C0C0BFA4999080",
 -2497 => x"C0C0C0BFA49990F8",
 -2496 => x"C0C0C0BFA4999082",
 -2495 => x"C0C0C0BFA4999092",
 -2494 => x"C0C0C0BFA4999099",
 -2493 => x"C0C0C0BFA49990B0",
 -2492 => x"C0C0C0BFA49990A4",
 -2491 => x"C0C0C0BFA49990F9",
 -2490 => x"C0C0C0BFA49990C0",
 -2489 => x"C0C0C0BFA4998090",
 -2488 => x"C0C0C0BFA4998080",
 -2487 => x"C0C0C0BFA49980F8",
 -2486 => x"C0C0C0BFA4998082",
 -2485 => x"C0C0C0BFA4998092",
 -2484 => x"C0C0C0BFA4998099",
 -2483 => x"C0C0C0BFA49980B0",
 -2482 => x"C0C0C0BFA49980A4",
 -2481 => x"C0C0C0BFA49980F9",
 -2480 => x"C0C0C0BFA49980C0",
 -2479 => x"C0C0C0BFA499F890",
 -2478 => x"C0C0C0BFA499F880",
 -2477 => x"C0C0C0BFA499F8F8",
 -2476 => x"C0C0C0BFA499F882",
 -2475 => x"C0C0C0BFA499F892",
 -2474 => x"C0C0C0BFA499F899",
 -2473 => x"C0C0C0BFA499F8B0",
 -2472 => x"C0C0C0BFA499F8A4",
 -2471 => x"C0C0C0BFA499F8F9",
 -2470 => x"C0C0C0BFA499F8C0",
 -2469 => x"C0C0C0BFA4998290",
 -2468 => x"C0C0C0BFA4998280",
 -2467 => x"C0C0C0BFA49982F8",
 -2466 => x"C0C0C0BFA4998282",
 -2465 => x"C0C0C0BFA4998292",
 -2464 => x"C0C0C0BFA4998299",
 -2463 => x"C0C0C0BFA49982B0",
 -2462 => x"C0C0C0BFA49982A4",
 -2461 => x"C0C0C0BFA49982F9",
 -2460 => x"C0C0C0BFA49982C0",
 -2459 => x"C0C0C0BFA4999290",
 -2458 => x"C0C0C0BFA4999280",
 -2457 => x"C0C0C0BFA49992F8",
 -2456 => x"C0C0C0BFA4999282",
 -2455 => x"C0C0C0BFA4999292",
 -2454 => x"C0C0C0BFA4999299",
 -2453 => x"C0C0C0BFA49992B0",
 -2452 => x"C0C0C0BFA49992A4",
 -2451 => x"C0C0C0BFA49992F9",
 -2450 => x"C0C0C0BFA49992C0",
 -2449 => x"C0C0C0BFA4999990",
 -2448 => x"C0C0C0BFA4999980",
 -2447 => x"C0C0C0BFA49999F8",
 -2446 => x"C0C0C0BFA4999982",
 -2445 => x"C0C0C0BFA4999992",
 -2444 => x"C0C0C0BFA4999999",
 -2443 => x"C0C0C0BFA49999B0",
 -2442 => x"C0C0C0BFA49999A4",
 -2441 => x"C0C0C0BFA49999F9",
 -2440 => x"C0C0C0BFA49999C0",
 -2439 => x"C0C0C0BFA499B090",
 -2438 => x"C0C0C0BFA499B080",
 -2437 => x"C0C0C0BFA499B0F8",
 -2436 => x"C0C0C0BFA499B082",
 -2435 => x"C0C0C0BFA499B092",
 -2434 => x"C0C0C0BFA499B099",
 -2433 => x"C0C0C0BFA499B0B0",
 -2432 => x"C0C0C0BFA499B0A4",
 -2431 => x"C0C0C0BFA499B0F9",
 -2430 => x"C0C0C0BFA499B0C0",
 -2429 => x"C0C0C0BFA499A490",
 -2428 => x"C0C0C0BFA499A480",
 -2427 => x"C0C0C0BFA499A4F8",
 -2426 => x"C0C0C0BFA499A482",
 -2425 => x"C0C0C0BFA499A492",
 -2424 => x"C0C0C0BFA499A499",
 -2423 => x"C0C0C0BFA499A4B0",
 -2422 => x"C0C0C0BFA499A4A4",
 -2421 => x"C0C0C0BFA499A4F9",
 -2420 => x"C0C0C0BFA499A4C0",
 -2419 => x"C0C0C0BFA499F990",
 -2418 => x"C0C0C0BFA499F980",
 -2417 => x"C0C0C0BFA499F9F8",
 -2416 => x"C0C0C0BFA499F982",
 -2415 => x"C0C0C0BFA499F992",
 -2414 => x"C0C0C0BFA499F999",
 -2413 => x"C0C0C0BFA499F9B0",
 -2412 => x"C0C0C0BFA499F9A4",
 -2411 => x"C0C0C0BFA499F9F9",
 -2410 => x"C0C0C0BFA499F9C0",
 -2409 => x"C0C0C0BFA499C090",
 -2408 => x"C0C0C0BFA499C080",
 -2407 => x"C0C0C0BFA499C0F8",
 -2406 => x"C0C0C0BFA499C082",
 -2405 => x"C0C0C0BFA499C092",
 -2404 => x"C0C0C0BFA499C099",
 -2403 => x"C0C0C0BFA499C0B0",
 -2402 => x"C0C0C0BFA499C0A4",
 -2401 => x"C0C0C0BFA499C0F9",
 -2400 => x"C0C0C0BFA499C0C0",
 -2399 => x"C0C0C0BFA4B09090",
 -2398 => x"C0C0C0BFA4B09080",
 -2397 => x"C0C0C0BFA4B090F8",
 -2396 => x"C0C0C0BFA4B09082",
 -2395 => x"C0C0C0BFA4B09092",
 -2394 => x"C0C0C0BFA4B09099",
 -2393 => x"C0C0C0BFA4B090B0",
 -2392 => x"C0C0C0BFA4B090A4",
 -2391 => x"C0C0C0BFA4B090F9",
 -2390 => x"C0C0C0BFA4B090C0",
 -2389 => x"C0C0C0BFA4B08090",
 -2388 => x"C0C0C0BFA4B08080",
 -2387 => x"C0C0C0BFA4B080F8",
 -2386 => x"C0C0C0BFA4B08082",
 -2385 => x"C0C0C0BFA4B08092",
 -2384 => x"C0C0C0BFA4B08099",
 -2383 => x"C0C0C0BFA4B080B0",
 -2382 => x"C0C0C0BFA4B080A4",
 -2381 => x"C0C0C0BFA4B080F9",
 -2380 => x"C0C0C0BFA4B080C0",
 -2379 => x"C0C0C0BFA4B0F890",
 -2378 => x"C0C0C0BFA4B0F880",
 -2377 => x"C0C0C0BFA4B0F8F8",
 -2376 => x"C0C0C0BFA4B0F882",
 -2375 => x"C0C0C0BFA4B0F892",
 -2374 => x"C0C0C0BFA4B0F899",
 -2373 => x"C0C0C0BFA4B0F8B0",
 -2372 => x"C0C0C0BFA4B0F8A4",
 -2371 => x"C0C0C0BFA4B0F8F9",
 -2370 => x"C0C0C0BFA4B0F8C0",
 -2369 => x"C0C0C0BFA4B08290",
 -2368 => x"C0C0C0BFA4B08280",
 -2367 => x"C0C0C0BFA4B082F8",
 -2366 => x"C0C0C0BFA4B08282",
 -2365 => x"C0C0C0BFA4B08292",
 -2364 => x"C0C0C0BFA4B08299",
 -2363 => x"C0C0C0BFA4B082B0",
 -2362 => x"C0C0C0BFA4B082A4",
 -2361 => x"C0C0C0BFA4B082F9",
 -2360 => x"C0C0C0BFA4B082C0",
 -2359 => x"C0C0C0BFA4B09290",
 -2358 => x"C0C0C0BFA4B09280",
 -2357 => x"C0C0C0BFA4B092F8",
 -2356 => x"C0C0C0BFA4B09282",
 -2355 => x"C0C0C0BFA4B09292",
 -2354 => x"C0C0C0BFA4B09299",
 -2353 => x"C0C0C0BFA4B092B0",
 -2352 => x"C0C0C0BFA4B092A4",
 -2351 => x"C0C0C0BFA4B092F9",
 -2350 => x"C0C0C0BFA4B092C0",
 -2349 => x"C0C0C0BFA4B09990",
 -2348 => x"C0C0C0BFA4B09980",
 -2347 => x"C0C0C0BFA4B099F8",
 -2346 => x"C0C0C0BFA4B09982",
 -2345 => x"C0C0C0BFA4B09992",
 -2344 => x"C0C0C0BFA4B09999",
 -2343 => x"C0C0C0BFA4B099B0",
 -2342 => x"C0C0C0BFA4B099A4",
 -2341 => x"C0C0C0BFA4B099F9",
 -2340 => x"C0C0C0BFA4B099C0",
 -2339 => x"C0C0C0BFA4B0B090",
 -2338 => x"C0C0C0BFA4B0B080",
 -2337 => x"C0C0C0BFA4B0B0F8",
 -2336 => x"C0C0C0BFA4B0B082",
 -2335 => x"C0C0C0BFA4B0B092",
 -2334 => x"C0C0C0BFA4B0B099",
 -2333 => x"C0C0C0BFA4B0B0B0",
 -2332 => x"C0C0C0BFA4B0B0A4",
 -2331 => x"C0C0C0BFA4B0B0F9",
 -2330 => x"C0C0C0BFA4B0B0C0",
 -2329 => x"C0C0C0BFA4B0A490",
 -2328 => x"C0C0C0BFA4B0A480",
 -2327 => x"C0C0C0BFA4B0A4F8",
 -2326 => x"C0C0C0BFA4B0A482",
 -2325 => x"C0C0C0BFA4B0A492",
 -2324 => x"C0C0C0BFA4B0A499",
 -2323 => x"C0C0C0BFA4B0A4B0",
 -2322 => x"C0C0C0BFA4B0A4A4",
 -2321 => x"C0C0C0BFA4B0A4F9",
 -2320 => x"C0C0C0BFA4B0A4C0",
 -2319 => x"C0C0C0BFA4B0F990",
 -2318 => x"C0C0C0BFA4B0F980",
 -2317 => x"C0C0C0BFA4B0F9F8",
 -2316 => x"C0C0C0BFA4B0F982",
 -2315 => x"C0C0C0BFA4B0F992",
 -2314 => x"C0C0C0BFA4B0F999",
 -2313 => x"C0C0C0BFA4B0F9B0",
 -2312 => x"C0C0C0BFA4B0F9A4",
 -2311 => x"C0C0C0BFA4B0F9F9",
 -2310 => x"C0C0C0BFA4B0F9C0",
 -2309 => x"C0C0C0BFA4B0C090",
 -2308 => x"C0C0C0BFA4B0C080",
 -2307 => x"C0C0C0BFA4B0C0F8",
 -2306 => x"C0C0C0BFA4B0C082",
 -2305 => x"C0C0C0BFA4B0C092",
 -2304 => x"C0C0C0BFA4B0C099",
 -2303 => x"C0C0C0BFA4B0C0B0",
 -2302 => x"C0C0C0BFA4B0C0A4",
 -2301 => x"C0C0C0BFA4B0C0F9",
 -2300 => x"C0C0C0BFA4B0C0C0",
 -2299 => x"C0C0C0BFA4A49090",
 -2298 => x"C0C0C0BFA4A49080",
 -2297 => x"C0C0C0BFA4A490F8",
 -2296 => x"C0C0C0BFA4A49082",
 -2295 => x"C0C0C0BFA4A49092",
 -2294 => x"C0C0C0BFA4A49099",
 -2293 => x"C0C0C0BFA4A490B0",
 -2292 => x"C0C0C0BFA4A490A4",
 -2291 => x"C0C0C0BFA4A490F9",
 -2290 => x"C0C0C0BFA4A490C0",
 -2289 => x"C0C0C0BFA4A48090",
 -2288 => x"C0C0C0BFA4A48080",
 -2287 => x"C0C0C0BFA4A480F8",
 -2286 => x"C0C0C0BFA4A48082",
 -2285 => x"C0C0C0BFA4A48092",
 -2284 => x"C0C0C0BFA4A48099",
 -2283 => x"C0C0C0BFA4A480B0",
 -2282 => x"C0C0C0BFA4A480A4",
 -2281 => x"C0C0C0BFA4A480F9",
 -2280 => x"C0C0C0BFA4A480C0",
 -2279 => x"C0C0C0BFA4A4F890",
 -2278 => x"C0C0C0BFA4A4F880",
 -2277 => x"C0C0C0BFA4A4F8F8",
 -2276 => x"C0C0C0BFA4A4F882",
 -2275 => x"C0C0C0BFA4A4F892",
 -2274 => x"C0C0C0BFA4A4F899",
 -2273 => x"C0C0C0BFA4A4F8B0",
 -2272 => x"C0C0C0BFA4A4F8A4",
 -2271 => x"C0C0C0BFA4A4F8F9",
 -2270 => x"C0C0C0BFA4A4F8C0",
 -2269 => x"C0C0C0BFA4A48290",
 -2268 => x"C0C0C0BFA4A48280",
 -2267 => x"C0C0C0BFA4A482F8",
 -2266 => x"C0C0C0BFA4A48282",
 -2265 => x"C0C0C0BFA4A48292",
 -2264 => x"C0C0C0BFA4A48299",
 -2263 => x"C0C0C0BFA4A482B0",
 -2262 => x"C0C0C0BFA4A482A4",
 -2261 => x"C0C0C0BFA4A482F9",
 -2260 => x"C0C0C0BFA4A482C0",
 -2259 => x"C0C0C0BFA4A49290",
 -2258 => x"C0C0C0BFA4A49280",
 -2257 => x"C0C0C0BFA4A492F8",
 -2256 => x"C0C0C0BFA4A49282",
 -2255 => x"C0C0C0BFA4A49292",
 -2254 => x"C0C0C0BFA4A49299",
 -2253 => x"C0C0C0BFA4A492B0",
 -2252 => x"C0C0C0BFA4A492A4",
 -2251 => x"C0C0C0BFA4A492F9",
 -2250 => x"C0C0C0BFA4A492C0",
 -2249 => x"C0C0C0BFA4A49990",
 -2248 => x"C0C0C0BFA4A49980",
 -2247 => x"C0C0C0BFA4A499F8",
 -2246 => x"C0C0C0BFA4A49982",
 -2245 => x"C0C0C0BFA4A49992",
 -2244 => x"C0C0C0BFA4A49999",
 -2243 => x"C0C0C0BFA4A499B0",
 -2242 => x"C0C0C0BFA4A499A4",
 -2241 => x"C0C0C0BFA4A499F9",
 -2240 => x"C0C0C0BFA4A499C0",
 -2239 => x"C0C0C0BFA4A4B090",
 -2238 => x"C0C0C0BFA4A4B080",
 -2237 => x"C0C0C0BFA4A4B0F8",
 -2236 => x"C0C0C0BFA4A4B082",
 -2235 => x"C0C0C0BFA4A4B092",
 -2234 => x"C0C0C0BFA4A4B099",
 -2233 => x"C0C0C0BFA4A4B0B0",
 -2232 => x"C0C0C0BFA4A4B0A4",
 -2231 => x"C0C0C0BFA4A4B0F9",
 -2230 => x"C0C0C0BFA4A4B0C0",
 -2229 => x"C0C0C0BFA4A4A490",
 -2228 => x"C0C0C0BFA4A4A480",
 -2227 => x"C0C0C0BFA4A4A4F8",
 -2226 => x"C0C0C0BFA4A4A482",
 -2225 => x"C0C0C0BFA4A4A492",
 -2224 => x"C0C0C0BFA4A4A499",
 -2223 => x"C0C0C0BFA4A4A4B0",
 -2222 => x"C0C0C0BFA4A4A4A4",
 -2221 => x"C0C0C0BFA4A4A4F9",
 -2220 => x"C0C0C0BFA4A4A4C0",
 -2219 => x"C0C0C0BFA4A4F990",
 -2218 => x"C0C0C0BFA4A4F980",
 -2217 => x"C0C0C0BFA4A4F9F8",
 -2216 => x"C0C0C0BFA4A4F982",
 -2215 => x"C0C0C0BFA4A4F992",
 -2214 => x"C0C0C0BFA4A4F999",
 -2213 => x"C0C0C0BFA4A4F9B0",
 -2212 => x"C0C0C0BFA4A4F9A4",
 -2211 => x"C0C0C0BFA4A4F9F9",
 -2210 => x"C0C0C0BFA4A4F9C0",
 -2209 => x"C0C0C0BFA4A4C090",
 -2208 => x"C0C0C0BFA4A4C080",
 -2207 => x"C0C0C0BFA4A4C0F8",
 -2206 => x"C0C0C0BFA4A4C082",
 -2205 => x"C0C0C0BFA4A4C092",
 -2204 => x"C0C0C0BFA4A4C099",
 -2203 => x"C0C0C0BFA4A4C0B0",
 -2202 => x"C0C0C0BFA4A4C0A4",
 -2201 => x"C0C0C0BFA4A4C0F9",
 -2200 => x"C0C0C0BFA4A4C0C0",
 -2199 => x"C0C0C0BFA4F99090",
 -2198 => x"C0C0C0BFA4F99080",
 -2197 => x"C0C0C0BFA4F990F8",
 -2196 => x"C0C0C0BFA4F99082",
 -2195 => x"C0C0C0BFA4F99092",
 -2194 => x"C0C0C0BFA4F99099",
 -2193 => x"C0C0C0BFA4F990B0",
 -2192 => x"C0C0C0BFA4F990A4",
 -2191 => x"C0C0C0BFA4F990F9",
 -2190 => x"C0C0C0BFA4F990C0",
 -2189 => x"C0C0C0BFA4F98090",
 -2188 => x"C0C0C0BFA4F98080",
 -2187 => x"C0C0C0BFA4F980F8",
 -2186 => x"C0C0C0BFA4F98082",
 -2185 => x"C0C0C0BFA4F98092",
 -2184 => x"C0C0C0BFA4F98099",
 -2183 => x"C0C0C0BFA4F980B0",
 -2182 => x"C0C0C0BFA4F980A4",
 -2181 => x"C0C0C0BFA4F980F9",
 -2180 => x"C0C0C0BFA4F980C0",
 -2179 => x"C0C0C0BFA4F9F890",
 -2178 => x"C0C0C0BFA4F9F880",
 -2177 => x"C0C0C0BFA4F9F8F8",
 -2176 => x"C0C0C0BFA4F9F882",
 -2175 => x"C0C0C0BFA4F9F892",
 -2174 => x"C0C0C0BFA4F9F899",
 -2173 => x"C0C0C0BFA4F9F8B0",
 -2172 => x"C0C0C0BFA4F9F8A4",
 -2171 => x"C0C0C0BFA4F9F8F9",
 -2170 => x"C0C0C0BFA4F9F8C0",
 -2169 => x"C0C0C0BFA4F98290",
 -2168 => x"C0C0C0BFA4F98280",
 -2167 => x"C0C0C0BFA4F982F8",
 -2166 => x"C0C0C0BFA4F98282",
 -2165 => x"C0C0C0BFA4F98292",
 -2164 => x"C0C0C0BFA4F98299",
 -2163 => x"C0C0C0BFA4F982B0",
 -2162 => x"C0C0C0BFA4F982A4",
 -2161 => x"C0C0C0BFA4F982F9",
 -2160 => x"C0C0C0BFA4F982C0",
 -2159 => x"C0C0C0BFA4F99290",
 -2158 => x"C0C0C0BFA4F99280",
 -2157 => x"C0C0C0BFA4F992F8",
 -2156 => x"C0C0C0BFA4F99282",
 -2155 => x"C0C0C0BFA4F99292",
 -2154 => x"C0C0C0BFA4F99299",
 -2153 => x"C0C0C0BFA4F992B0",
 -2152 => x"C0C0C0BFA4F992A4",
 -2151 => x"C0C0C0BFA4F992F9",
 -2150 => x"C0C0C0BFA4F992C0",
 -2149 => x"C0C0C0BFA4F99990",
 -2148 => x"C0C0C0BFA4F99980",
 -2147 => x"C0C0C0BFA4F999F8",
 -2146 => x"C0C0C0BFA4F99982",
 -2145 => x"C0C0C0BFA4F99992",
 -2144 => x"C0C0C0BFA4F99999",
 -2143 => x"C0C0C0BFA4F999B0",
 -2142 => x"C0C0C0BFA4F999A4",
 -2141 => x"C0C0C0BFA4F999F9",
 -2140 => x"C0C0C0BFA4F999C0",
 -2139 => x"C0C0C0BFA4F9B090",
 -2138 => x"C0C0C0BFA4F9B080",
 -2137 => x"C0C0C0BFA4F9B0F8",
 -2136 => x"C0C0C0BFA4F9B082",
 -2135 => x"C0C0C0BFA4F9B092",
 -2134 => x"C0C0C0BFA4F9B099",
 -2133 => x"C0C0C0BFA4F9B0B0",
 -2132 => x"C0C0C0BFA4F9B0A4",
 -2131 => x"C0C0C0BFA4F9B0F9",
 -2130 => x"C0C0C0BFA4F9B0C0",
 -2129 => x"C0C0C0BFA4F9A490",
 -2128 => x"C0C0C0BFA4F9A480",
 -2127 => x"C0C0C0BFA4F9A4F8",
 -2126 => x"C0C0C0BFA4F9A482",
 -2125 => x"C0C0C0BFA4F9A492",
 -2124 => x"C0C0C0BFA4F9A499",
 -2123 => x"C0C0C0BFA4F9A4B0",
 -2122 => x"C0C0C0BFA4F9A4A4",
 -2121 => x"C0C0C0BFA4F9A4F9",
 -2120 => x"C0C0C0BFA4F9A4C0",
 -2119 => x"C0C0C0BFA4F9F990",
 -2118 => x"C0C0C0BFA4F9F980",
 -2117 => x"C0C0C0BFA4F9F9F8",
 -2116 => x"C0C0C0BFA4F9F982",
 -2115 => x"C0C0C0BFA4F9F992",
 -2114 => x"C0C0C0BFA4F9F999",
 -2113 => x"C0C0C0BFA4F9F9B0",
 -2112 => x"C0C0C0BFA4F9F9A4",
 -2111 => x"C0C0C0BFA4F9F9F9",
 -2110 => x"C0C0C0BFA4F9F9C0",
 -2109 => x"C0C0C0BFA4F9C090",
 -2108 => x"C0C0C0BFA4F9C080",
 -2107 => x"C0C0C0BFA4F9C0F8",
 -2106 => x"C0C0C0BFA4F9C082",
 -2105 => x"C0C0C0BFA4F9C092",
 -2104 => x"C0C0C0BFA4F9C099",
 -2103 => x"C0C0C0BFA4F9C0B0",
 -2102 => x"C0C0C0BFA4F9C0A4",
 -2101 => x"C0C0C0BFA4F9C0F9",
 -2100 => x"C0C0C0BFA4F9C0C0",
 -2099 => x"C0C0C0BFA4C09090",
 -2098 => x"C0C0C0BFA4C09080",
 -2097 => x"C0C0C0BFA4C090F8",
 -2096 => x"C0C0C0BFA4C09082",
 -2095 => x"C0C0C0BFA4C09092",
 -2094 => x"C0C0C0BFA4C09099",
 -2093 => x"C0C0C0BFA4C090B0",
 -2092 => x"C0C0C0BFA4C090A4",
 -2091 => x"C0C0C0BFA4C090F9",
 -2090 => x"C0C0C0BFA4C090C0",
 -2089 => x"C0C0C0BFA4C08090",
 -2088 => x"C0C0C0BFA4C08080",
 -2087 => x"C0C0C0BFA4C080F8",
 -2086 => x"C0C0C0BFA4C08082",
 -2085 => x"C0C0C0BFA4C08092",
 -2084 => x"C0C0C0BFA4C08099",
 -2083 => x"C0C0C0BFA4C080B0",
 -2082 => x"C0C0C0BFA4C080A4",
 -2081 => x"C0C0C0BFA4C080F9",
 -2080 => x"C0C0C0BFA4C080C0",
 -2079 => x"C0C0C0BFA4C0F890",
 -2078 => x"C0C0C0BFA4C0F880",
 -2077 => x"C0C0C0BFA4C0F8F8",
 -2076 => x"C0C0C0BFA4C0F882",
 -2075 => x"C0C0C0BFA4C0F892",
 -2074 => x"C0C0C0BFA4C0F899",
 -2073 => x"C0C0C0BFA4C0F8B0",
 -2072 => x"C0C0C0BFA4C0F8A4",
 -2071 => x"C0C0C0BFA4C0F8F9",
 -2070 => x"C0C0C0BFA4C0F8C0",
 -2069 => x"C0C0C0BFA4C08290",
 -2068 => x"C0C0C0BFA4C08280",
 -2067 => x"C0C0C0BFA4C082F8",
 -2066 => x"C0C0C0BFA4C08282",
 -2065 => x"C0C0C0BFA4C08292",
 -2064 => x"C0C0C0BFA4C08299",
 -2063 => x"C0C0C0BFA4C082B0",
 -2062 => x"C0C0C0BFA4C082A4",
 -2061 => x"C0C0C0BFA4C082F9",
 -2060 => x"C0C0C0BFA4C082C0",
 -2059 => x"C0C0C0BFA4C09290",
 -2058 => x"C0C0C0BFA4C09280",
 -2057 => x"C0C0C0BFA4C092F8",
 -2056 => x"C0C0C0BFA4C09282",
 -2055 => x"C0C0C0BFA4C09292",
 -2054 => x"C0C0C0BFA4C09299",
 -2053 => x"C0C0C0BFA4C092B0",
 -2052 => x"C0C0C0BFA4C092A4",
 -2051 => x"C0C0C0BFA4C092F9",
 -2050 => x"C0C0C0BFA4C092C0",
 -2049 => x"C0C0C0BFA4C09990",
 -2048 => x"C0C0C0BFA4C09980",
 -2047 => x"C0C0C0BFA4C099F8",
 -2046 => x"C0C0C0BFA4C09982",
 -2045 => x"C0C0C0BFA4C09992",
 -2044 => x"C0C0C0BFA4C09999",
 -2043 => x"C0C0C0BFA4C099B0",
 -2042 => x"C0C0C0BFA4C099A4",
 -2041 => x"C0C0C0BFA4C099F9",
 -2040 => x"C0C0C0BFA4C099C0",
 -2039 => x"C0C0C0BFA4C0B090",
 -2038 => x"C0C0C0BFA4C0B080",
 -2037 => x"C0C0C0BFA4C0B0F8",
 -2036 => x"C0C0C0BFA4C0B082",
 -2035 => x"C0C0C0BFA4C0B092",
 -2034 => x"C0C0C0BFA4C0B099",
 -2033 => x"C0C0C0BFA4C0B0B0",
 -2032 => x"C0C0C0BFA4C0B0A4",
 -2031 => x"C0C0C0BFA4C0B0F9",
 -2030 => x"C0C0C0BFA4C0B0C0",
 -2029 => x"C0C0C0BFA4C0A490",
 -2028 => x"C0C0C0BFA4C0A480",
 -2027 => x"C0C0C0BFA4C0A4F8",
 -2026 => x"C0C0C0BFA4C0A482",
 -2025 => x"C0C0C0BFA4C0A492",
 -2024 => x"C0C0C0BFA4C0A499",
 -2023 => x"C0C0C0BFA4C0A4B0",
 -2022 => x"C0C0C0BFA4C0A4A4",
 -2021 => x"C0C0C0BFA4C0A4F9",
 -2020 => x"C0C0C0BFA4C0A4C0",
 -2019 => x"C0C0C0BFA4C0F990",
 -2018 => x"C0C0C0BFA4C0F980",
 -2017 => x"C0C0C0BFA4C0F9F8",
 -2016 => x"C0C0C0BFA4C0F982",
 -2015 => x"C0C0C0BFA4C0F992",
 -2014 => x"C0C0C0BFA4C0F999",
 -2013 => x"C0C0C0BFA4C0F9B0",
 -2012 => x"C0C0C0BFA4C0F9A4",
 -2011 => x"C0C0C0BFA4C0F9F9",
 -2010 => x"C0C0C0BFA4C0F9C0",
 -2009 => x"C0C0C0BFA4C0C090",
 -2008 => x"C0C0C0BFA4C0C080",
 -2007 => x"C0C0C0BFA4C0C0F8",
 -2006 => x"C0C0C0BFA4C0C082",
 -2005 => x"C0C0C0BFA4C0C092",
 -2004 => x"C0C0C0BFA4C0C099",
 -2003 => x"C0C0C0BFA4C0C0B0",
 -2002 => x"C0C0C0BFA4C0C0A4",
 -2001 => x"C0C0C0BFA4C0C0F9",
 -2000 => x"C0C0C0BFA4C0C0C0",
 -1999 => x"C0C0C0BFF9909090",
 -1998 => x"C0C0C0BFF9909080",
 -1997 => x"C0C0C0BFF99090F8",
 -1996 => x"C0C0C0BFF9909082",
 -1995 => x"C0C0C0BFF9909092",
 -1994 => x"C0C0C0BFF9909099",
 -1993 => x"C0C0C0BFF99090B0",
 -1992 => x"C0C0C0BFF99090A4",
 -1991 => x"C0C0C0BFF99090F9",
 -1990 => x"C0C0C0BFF99090C0",
 -1989 => x"C0C0C0BFF9908090",
 -1988 => x"C0C0C0BFF9908080",
 -1987 => x"C0C0C0BFF99080F8",
 -1986 => x"C0C0C0BFF9908082",
 -1985 => x"C0C0C0BFF9908092",
 -1984 => x"C0C0C0BFF9908099",
 -1983 => x"C0C0C0BFF99080B0",
 -1982 => x"C0C0C0BFF99080A4",
 -1981 => x"C0C0C0BFF99080F9",
 -1980 => x"C0C0C0BFF99080C0",
 -1979 => x"C0C0C0BFF990F890",
 -1978 => x"C0C0C0BFF990F880",
 -1977 => x"C0C0C0BFF990F8F8",
 -1976 => x"C0C0C0BFF990F882",
 -1975 => x"C0C0C0BFF990F892",
 -1974 => x"C0C0C0BFF990F899",
 -1973 => x"C0C0C0BFF990F8B0",
 -1972 => x"C0C0C0BFF990F8A4",
 -1971 => x"C0C0C0BFF990F8F9",
 -1970 => x"C0C0C0BFF990F8C0",
 -1969 => x"C0C0C0BFF9908290",
 -1968 => x"C0C0C0BFF9908280",
 -1967 => x"C0C0C0BFF99082F8",
 -1966 => x"C0C0C0BFF9908282",
 -1965 => x"C0C0C0BFF9908292",
 -1964 => x"C0C0C0BFF9908299",
 -1963 => x"C0C0C0BFF99082B0",
 -1962 => x"C0C0C0BFF99082A4",
 -1961 => x"C0C0C0BFF99082F9",
 -1960 => x"C0C0C0BFF99082C0",
 -1959 => x"C0C0C0BFF9909290",
 -1958 => x"C0C0C0BFF9909280",
 -1957 => x"C0C0C0BFF99092F8",
 -1956 => x"C0C0C0BFF9909282",
 -1955 => x"C0C0C0BFF9909292",
 -1954 => x"C0C0C0BFF9909299",
 -1953 => x"C0C0C0BFF99092B0",
 -1952 => x"C0C0C0BFF99092A4",
 -1951 => x"C0C0C0BFF99092F9",
 -1950 => x"C0C0C0BFF99092C0",
 -1949 => x"C0C0C0BFF9909990",
 -1948 => x"C0C0C0BFF9909980",
 -1947 => x"C0C0C0BFF99099F8",
 -1946 => x"C0C0C0BFF9909982",
 -1945 => x"C0C0C0BFF9909992",
 -1944 => x"C0C0C0BFF9909999",
 -1943 => x"C0C0C0BFF99099B0",
 -1942 => x"C0C0C0BFF99099A4",
 -1941 => x"C0C0C0BFF99099F9",
 -1940 => x"C0C0C0BFF99099C0",
 -1939 => x"C0C0C0BFF990B090",
 -1938 => x"C0C0C0BFF990B080",
 -1937 => x"C0C0C0BFF990B0F8",
 -1936 => x"C0C0C0BFF990B082",
 -1935 => x"C0C0C0BFF990B092",
 -1934 => x"C0C0C0BFF990B099",
 -1933 => x"C0C0C0BFF990B0B0",
 -1932 => x"C0C0C0BFF990B0A4",
 -1931 => x"C0C0C0BFF990B0F9",
 -1930 => x"C0C0C0BFF990B0C0",
 -1929 => x"C0C0C0BFF990A490",
 -1928 => x"C0C0C0BFF990A480",
 -1927 => x"C0C0C0BFF990A4F8",
 -1926 => x"C0C0C0BFF990A482",
 -1925 => x"C0C0C0BFF990A492",
 -1924 => x"C0C0C0BFF990A499",
 -1923 => x"C0C0C0BFF990A4B0",
 -1922 => x"C0C0C0BFF990A4A4",
 -1921 => x"C0C0C0BFF990A4F9",
 -1920 => x"C0C0C0BFF990A4C0",
 -1919 => x"C0C0C0BFF990F990",
 -1918 => x"C0C0C0BFF990F980",
 -1917 => x"C0C0C0BFF990F9F8",
 -1916 => x"C0C0C0BFF990F982",
 -1915 => x"C0C0C0BFF990F992",
 -1914 => x"C0C0C0BFF990F999",
 -1913 => x"C0C0C0BFF990F9B0",
 -1912 => x"C0C0C0BFF990F9A4",
 -1911 => x"C0C0C0BFF990F9F9",
 -1910 => x"C0C0C0BFF990F9C0",
 -1909 => x"C0C0C0BFF990C090",
 -1908 => x"C0C0C0BFF990C080",
 -1907 => x"C0C0C0BFF990C0F8",
 -1906 => x"C0C0C0BFF990C082",
 -1905 => x"C0C0C0BFF990C092",
 -1904 => x"C0C0C0BFF990C099",
 -1903 => x"C0C0C0BFF990C0B0",
 -1902 => x"C0C0C0BFF990C0A4",
 -1901 => x"C0C0C0BFF990C0F9",
 -1900 => x"C0C0C0BFF990C0C0",
 -1899 => x"C0C0C0BFF9809090",
 -1898 => x"C0C0C0BFF9809080",
 -1897 => x"C0C0C0BFF98090F8",
 -1896 => x"C0C0C0BFF9809082",
 -1895 => x"C0C0C0BFF9809092",
 -1894 => x"C0C0C0BFF9809099",
 -1893 => x"C0C0C0BFF98090B0",
 -1892 => x"C0C0C0BFF98090A4",
 -1891 => x"C0C0C0BFF98090F9",
 -1890 => x"C0C0C0BFF98090C0",
 -1889 => x"C0C0C0BFF9808090",
 -1888 => x"C0C0C0BFF9808080",
 -1887 => x"C0C0C0BFF98080F8",
 -1886 => x"C0C0C0BFF9808082",
 -1885 => x"C0C0C0BFF9808092",
 -1884 => x"C0C0C0BFF9808099",
 -1883 => x"C0C0C0BFF98080B0",
 -1882 => x"C0C0C0BFF98080A4",
 -1881 => x"C0C0C0BFF98080F9",
 -1880 => x"C0C0C0BFF98080C0",
 -1879 => x"C0C0C0BFF980F890",
 -1878 => x"C0C0C0BFF980F880",
 -1877 => x"C0C0C0BFF980F8F8",
 -1876 => x"C0C0C0BFF980F882",
 -1875 => x"C0C0C0BFF980F892",
 -1874 => x"C0C0C0BFF980F899",
 -1873 => x"C0C0C0BFF980F8B0",
 -1872 => x"C0C0C0BFF980F8A4",
 -1871 => x"C0C0C0BFF980F8F9",
 -1870 => x"C0C0C0BFF980F8C0",
 -1869 => x"C0C0C0BFF9808290",
 -1868 => x"C0C0C0BFF9808280",
 -1867 => x"C0C0C0BFF98082F8",
 -1866 => x"C0C0C0BFF9808282",
 -1865 => x"C0C0C0BFF9808292",
 -1864 => x"C0C0C0BFF9808299",
 -1863 => x"C0C0C0BFF98082B0",
 -1862 => x"C0C0C0BFF98082A4",
 -1861 => x"C0C0C0BFF98082F9",
 -1860 => x"C0C0C0BFF98082C0",
 -1859 => x"C0C0C0BFF9809290",
 -1858 => x"C0C0C0BFF9809280",
 -1857 => x"C0C0C0BFF98092F8",
 -1856 => x"C0C0C0BFF9809282",
 -1855 => x"C0C0C0BFF9809292",
 -1854 => x"C0C0C0BFF9809299",
 -1853 => x"C0C0C0BFF98092B0",
 -1852 => x"C0C0C0BFF98092A4",
 -1851 => x"C0C0C0BFF98092F9",
 -1850 => x"C0C0C0BFF98092C0",
 -1849 => x"C0C0C0BFF9809990",
 -1848 => x"C0C0C0BFF9809980",
 -1847 => x"C0C0C0BFF98099F8",
 -1846 => x"C0C0C0BFF9809982",
 -1845 => x"C0C0C0BFF9809992",
 -1844 => x"C0C0C0BFF9809999",
 -1843 => x"C0C0C0BFF98099B0",
 -1842 => x"C0C0C0BFF98099A4",
 -1841 => x"C0C0C0BFF98099F9",
 -1840 => x"C0C0C0BFF98099C0",
 -1839 => x"C0C0C0BFF980B090",
 -1838 => x"C0C0C0BFF980B080",
 -1837 => x"C0C0C0BFF980B0F8",
 -1836 => x"C0C0C0BFF980B082",
 -1835 => x"C0C0C0BFF980B092",
 -1834 => x"C0C0C0BFF980B099",
 -1833 => x"C0C0C0BFF980B0B0",
 -1832 => x"C0C0C0BFF980B0A4",
 -1831 => x"C0C0C0BFF980B0F9",
 -1830 => x"C0C0C0BFF980B0C0",
 -1829 => x"C0C0C0BFF980A490",
 -1828 => x"C0C0C0BFF980A480",
 -1827 => x"C0C0C0BFF980A4F8",
 -1826 => x"C0C0C0BFF980A482",
 -1825 => x"C0C0C0BFF980A492",
 -1824 => x"C0C0C0BFF980A499",
 -1823 => x"C0C0C0BFF980A4B0",
 -1822 => x"C0C0C0BFF980A4A4",
 -1821 => x"C0C0C0BFF980A4F9",
 -1820 => x"C0C0C0BFF980A4C0",
 -1819 => x"C0C0C0BFF980F990",
 -1818 => x"C0C0C0BFF980F980",
 -1817 => x"C0C0C0BFF980F9F8",
 -1816 => x"C0C0C0BFF980F982",
 -1815 => x"C0C0C0BFF980F992",
 -1814 => x"C0C0C0BFF980F999",
 -1813 => x"C0C0C0BFF980F9B0",
 -1812 => x"C0C0C0BFF980F9A4",
 -1811 => x"C0C0C0BFF980F9F9",
 -1810 => x"C0C0C0BFF980F9C0",
 -1809 => x"C0C0C0BFF980C090",
 -1808 => x"C0C0C0BFF980C080",
 -1807 => x"C0C0C0BFF980C0F8",
 -1806 => x"C0C0C0BFF980C082",
 -1805 => x"C0C0C0BFF980C092",
 -1804 => x"C0C0C0BFF980C099",
 -1803 => x"C0C0C0BFF980C0B0",
 -1802 => x"C0C0C0BFF980C0A4",
 -1801 => x"C0C0C0BFF980C0F9",
 -1800 => x"C0C0C0BFF980C0C0",
 -1799 => x"C0C0C0BFF9F89090",
 -1798 => x"C0C0C0BFF9F89080",
 -1797 => x"C0C0C0BFF9F890F8",
 -1796 => x"C0C0C0BFF9F89082",
 -1795 => x"C0C0C0BFF9F89092",
 -1794 => x"C0C0C0BFF9F89099",
 -1793 => x"C0C0C0BFF9F890B0",
 -1792 => x"C0C0C0BFF9F890A4",
 -1791 => x"C0C0C0BFF9F890F9",
 -1790 => x"C0C0C0BFF9F890C0",
 -1789 => x"C0C0C0BFF9F88090",
 -1788 => x"C0C0C0BFF9F88080",
 -1787 => x"C0C0C0BFF9F880F8",
 -1786 => x"C0C0C0BFF9F88082",
 -1785 => x"C0C0C0BFF9F88092",
 -1784 => x"C0C0C0BFF9F88099",
 -1783 => x"C0C0C0BFF9F880B0",
 -1782 => x"C0C0C0BFF9F880A4",
 -1781 => x"C0C0C0BFF9F880F9",
 -1780 => x"C0C0C0BFF9F880C0",
 -1779 => x"C0C0C0BFF9F8F890",
 -1778 => x"C0C0C0BFF9F8F880",
 -1777 => x"C0C0C0BFF9F8F8F8",
 -1776 => x"C0C0C0BFF9F8F882",
 -1775 => x"C0C0C0BFF9F8F892",
 -1774 => x"C0C0C0BFF9F8F899",
 -1773 => x"C0C0C0BFF9F8F8B0",
 -1772 => x"C0C0C0BFF9F8F8A4",
 -1771 => x"C0C0C0BFF9F8F8F9",
 -1770 => x"C0C0C0BFF9F8F8C0",
 -1769 => x"C0C0C0BFF9F88290",
 -1768 => x"C0C0C0BFF9F88280",
 -1767 => x"C0C0C0BFF9F882F8",
 -1766 => x"C0C0C0BFF9F88282",
 -1765 => x"C0C0C0BFF9F88292",
 -1764 => x"C0C0C0BFF9F88299",
 -1763 => x"C0C0C0BFF9F882B0",
 -1762 => x"C0C0C0BFF9F882A4",
 -1761 => x"C0C0C0BFF9F882F9",
 -1760 => x"C0C0C0BFF9F882C0",
 -1759 => x"C0C0C0BFF9F89290",
 -1758 => x"C0C0C0BFF9F89280",
 -1757 => x"C0C0C0BFF9F892F8",
 -1756 => x"C0C0C0BFF9F89282",
 -1755 => x"C0C0C0BFF9F89292",
 -1754 => x"C0C0C0BFF9F89299",
 -1753 => x"C0C0C0BFF9F892B0",
 -1752 => x"C0C0C0BFF9F892A4",
 -1751 => x"C0C0C0BFF9F892F9",
 -1750 => x"C0C0C0BFF9F892C0",
 -1749 => x"C0C0C0BFF9F89990",
 -1748 => x"C0C0C0BFF9F89980",
 -1747 => x"C0C0C0BFF9F899F8",
 -1746 => x"C0C0C0BFF9F89982",
 -1745 => x"C0C0C0BFF9F89992",
 -1744 => x"C0C0C0BFF9F89999",
 -1743 => x"C0C0C0BFF9F899B0",
 -1742 => x"C0C0C0BFF9F899A4",
 -1741 => x"C0C0C0BFF9F899F9",
 -1740 => x"C0C0C0BFF9F899C0",
 -1739 => x"C0C0C0BFF9F8B090",
 -1738 => x"C0C0C0BFF9F8B080",
 -1737 => x"C0C0C0BFF9F8B0F8",
 -1736 => x"C0C0C0BFF9F8B082",
 -1735 => x"C0C0C0BFF9F8B092",
 -1734 => x"C0C0C0BFF9F8B099",
 -1733 => x"C0C0C0BFF9F8B0B0",
 -1732 => x"C0C0C0BFF9F8B0A4",
 -1731 => x"C0C0C0BFF9F8B0F9",
 -1730 => x"C0C0C0BFF9F8B0C0",
 -1729 => x"C0C0C0BFF9F8A490",
 -1728 => x"C0C0C0BFF9F8A480",
 -1727 => x"C0C0C0BFF9F8A4F8",
 -1726 => x"C0C0C0BFF9F8A482",
 -1725 => x"C0C0C0BFF9F8A492",
 -1724 => x"C0C0C0BFF9F8A499",
 -1723 => x"C0C0C0BFF9F8A4B0",
 -1722 => x"C0C0C0BFF9F8A4A4",
 -1721 => x"C0C0C0BFF9F8A4F9",
 -1720 => x"C0C0C0BFF9F8A4C0",
 -1719 => x"C0C0C0BFF9F8F990",
 -1718 => x"C0C0C0BFF9F8F980",
 -1717 => x"C0C0C0BFF9F8F9F8",
 -1716 => x"C0C0C0BFF9F8F982",
 -1715 => x"C0C0C0BFF9F8F992",
 -1714 => x"C0C0C0BFF9F8F999",
 -1713 => x"C0C0C0BFF9F8F9B0",
 -1712 => x"C0C0C0BFF9F8F9A4",
 -1711 => x"C0C0C0BFF9F8F9F9",
 -1710 => x"C0C0C0BFF9F8F9C0",
 -1709 => x"C0C0C0BFF9F8C090",
 -1708 => x"C0C0C0BFF9F8C080",
 -1707 => x"C0C0C0BFF9F8C0F8",
 -1706 => x"C0C0C0BFF9F8C082",
 -1705 => x"C0C0C0BFF9F8C092",
 -1704 => x"C0C0C0BFF9F8C099",
 -1703 => x"C0C0C0BFF9F8C0B0",
 -1702 => x"C0C0C0BFF9F8C0A4",
 -1701 => x"C0C0C0BFF9F8C0F9",
 -1700 => x"C0C0C0BFF9F8C0C0",
 -1699 => x"C0C0C0BFF9829090",
 -1698 => x"C0C0C0BFF9829080",
 -1697 => x"C0C0C0BFF98290F8",
 -1696 => x"C0C0C0BFF9829082",
 -1695 => x"C0C0C0BFF9829092",
 -1694 => x"C0C0C0BFF9829099",
 -1693 => x"C0C0C0BFF98290B0",
 -1692 => x"C0C0C0BFF98290A4",
 -1691 => x"C0C0C0BFF98290F9",
 -1690 => x"C0C0C0BFF98290C0",
 -1689 => x"C0C0C0BFF9828090",
 -1688 => x"C0C0C0BFF9828080",
 -1687 => x"C0C0C0BFF98280F8",
 -1686 => x"C0C0C0BFF9828082",
 -1685 => x"C0C0C0BFF9828092",
 -1684 => x"C0C0C0BFF9828099",
 -1683 => x"C0C0C0BFF98280B0",
 -1682 => x"C0C0C0BFF98280A4",
 -1681 => x"C0C0C0BFF98280F9",
 -1680 => x"C0C0C0BFF98280C0",
 -1679 => x"C0C0C0BFF982F890",
 -1678 => x"C0C0C0BFF982F880",
 -1677 => x"C0C0C0BFF982F8F8",
 -1676 => x"C0C0C0BFF982F882",
 -1675 => x"C0C0C0BFF982F892",
 -1674 => x"C0C0C0BFF982F899",
 -1673 => x"C0C0C0BFF982F8B0",
 -1672 => x"C0C0C0BFF982F8A4",
 -1671 => x"C0C0C0BFF982F8F9",
 -1670 => x"C0C0C0BFF982F8C0",
 -1669 => x"C0C0C0BFF9828290",
 -1668 => x"C0C0C0BFF9828280",
 -1667 => x"C0C0C0BFF98282F8",
 -1666 => x"C0C0C0BFF9828282",
 -1665 => x"C0C0C0BFF9828292",
 -1664 => x"C0C0C0BFF9828299",
 -1663 => x"C0C0C0BFF98282B0",
 -1662 => x"C0C0C0BFF98282A4",
 -1661 => x"C0C0C0BFF98282F9",
 -1660 => x"C0C0C0BFF98282C0",
 -1659 => x"C0C0C0BFF9829290",
 -1658 => x"C0C0C0BFF9829280",
 -1657 => x"C0C0C0BFF98292F8",
 -1656 => x"C0C0C0BFF9829282",
 -1655 => x"C0C0C0BFF9829292",
 -1654 => x"C0C0C0BFF9829299",
 -1653 => x"C0C0C0BFF98292B0",
 -1652 => x"C0C0C0BFF98292A4",
 -1651 => x"C0C0C0BFF98292F9",
 -1650 => x"C0C0C0BFF98292C0",
 -1649 => x"C0C0C0BFF9829990",
 -1648 => x"C0C0C0BFF9829980",
 -1647 => x"C0C0C0BFF98299F8",
 -1646 => x"C0C0C0BFF9829982",
 -1645 => x"C0C0C0BFF9829992",
 -1644 => x"C0C0C0BFF9829999",
 -1643 => x"C0C0C0BFF98299B0",
 -1642 => x"C0C0C0BFF98299A4",
 -1641 => x"C0C0C0BFF98299F9",
 -1640 => x"C0C0C0BFF98299C0",
 -1639 => x"C0C0C0BFF982B090",
 -1638 => x"C0C0C0BFF982B080",
 -1637 => x"C0C0C0BFF982B0F8",
 -1636 => x"C0C0C0BFF982B082",
 -1635 => x"C0C0C0BFF982B092",
 -1634 => x"C0C0C0BFF982B099",
 -1633 => x"C0C0C0BFF982B0B0",
 -1632 => x"C0C0C0BFF982B0A4",
 -1631 => x"C0C0C0BFF982B0F9",
 -1630 => x"C0C0C0BFF982B0C0",
 -1629 => x"C0C0C0BFF982A490",
 -1628 => x"C0C0C0BFF982A480",
 -1627 => x"C0C0C0BFF982A4F8",
 -1626 => x"C0C0C0BFF982A482",
 -1625 => x"C0C0C0BFF982A492",
 -1624 => x"C0C0C0BFF982A499",
 -1623 => x"C0C0C0BFF982A4B0",
 -1622 => x"C0C0C0BFF982A4A4",
 -1621 => x"C0C0C0BFF982A4F9",
 -1620 => x"C0C0C0BFF982A4C0",
 -1619 => x"C0C0C0BFF982F990",
 -1618 => x"C0C0C0BFF982F980",
 -1617 => x"C0C0C0BFF982F9F8",
 -1616 => x"C0C0C0BFF982F982",
 -1615 => x"C0C0C0BFF982F992",
 -1614 => x"C0C0C0BFF982F999",
 -1613 => x"C0C0C0BFF982F9B0",
 -1612 => x"C0C0C0BFF982F9A4",
 -1611 => x"C0C0C0BFF982F9F9",
 -1610 => x"C0C0C0BFF982F9C0",
 -1609 => x"C0C0C0BFF982C090",
 -1608 => x"C0C0C0BFF982C080",
 -1607 => x"C0C0C0BFF982C0F8",
 -1606 => x"C0C0C0BFF982C082",
 -1605 => x"C0C0C0BFF982C092",
 -1604 => x"C0C0C0BFF982C099",
 -1603 => x"C0C0C0BFF982C0B0",
 -1602 => x"C0C0C0BFF982C0A4",
 -1601 => x"C0C0C0BFF982C0F9",
 -1600 => x"C0C0C0BFF982C0C0",
 -1599 => x"C0C0C0BFF9929090",
 -1598 => x"C0C0C0BFF9929080",
 -1597 => x"C0C0C0BFF99290F8",
 -1596 => x"C0C0C0BFF9929082",
 -1595 => x"C0C0C0BFF9929092",
 -1594 => x"C0C0C0BFF9929099",
 -1593 => x"C0C0C0BFF99290B0",
 -1592 => x"C0C0C0BFF99290A4",
 -1591 => x"C0C0C0BFF99290F9",
 -1590 => x"C0C0C0BFF99290C0",
 -1589 => x"C0C0C0BFF9928090",
 -1588 => x"C0C0C0BFF9928080",
 -1587 => x"C0C0C0BFF99280F8",
 -1586 => x"C0C0C0BFF9928082",
 -1585 => x"C0C0C0BFF9928092",
 -1584 => x"C0C0C0BFF9928099",
 -1583 => x"C0C0C0BFF99280B0",
 -1582 => x"C0C0C0BFF99280A4",
 -1581 => x"C0C0C0BFF99280F9",
 -1580 => x"C0C0C0BFF99280C0",
 -1579 => x"C0C0C0BFF992F890",
 -1578 => x"C0C0C0BFF992F880",
 -1577 => x"C0C0C0BFF992F8F8",
 -1576 => x"C0C0C0BFF992F882",
 -1575 => x"C0C0C0BFF992F892",
 -1574 => x"C0C0C0BFF992F899",
 -1573 => x"C0C0C0BFF992F8B0",
 -1572 => x"C0C0C0BFF992F8A4",
 -1571 => x"C0C0C0BFF992F8F9",
 -1570 => x"C0C0C0BFF992F8C0",
 -1569 => x"C0C0C0BFF9928290",
 -1568 => x"C0C0C0BFF9928280",
 -1567 => x"C0C0C0BFF99282F8",
 -1566 => x"C0C0C0BFF9928282",
 -1565 => x"C0C0C0BFF9928292",
 -1564 => x"C0C0C0BFF9928299",
 -1563 => x"C0C0C0BFF99282B0",
 -1562 => x"C0C0C0BFF99282A4",
 -1561 => x"C0C0C0BFF99282F9",
 -1560 => x"C0C0C0BFF99282C0",
 -1559 => x"C0C0C0BFF9929290",
 -1558 => x"C0C0C0BFF9929280",
 -1557 => x"C0C0C0BFF99292F8",
 -1556 => x"C0C0C0BFF9929282",
 -1555 => x"C0C0C0BFF9929292",
 -1554 => x"C0C0C0BFF9929299",
 -1553 => x"C0C0C0BFF99292B0",
 -1552 => x"C0C0C0BFF99292A4",
 -1551 => x"C0C0C0BFF99292F9",
 -1550 => x"C0C0C0BFF99292C0",
 -1549 => x"C0C0C0BFF9929990",
 -1548 => x"C0C0C0BFF9929980",
 -1547 => x"C0C0C0BFF99299F8",
 -1546 => x"C0C0C0BFF9929982",
 -1545 => x"C0C0C0BFF9929992",
 -1544 => x"C0C0C0BFF9929999",
 -1543 => x"C0C0C0BFF99299B0",
 -1542 => x"C0C0C0BFF99299A4",
 -1541 => x"C0C0C0BFF99299F9",
 -1540 => x"C0C0C0BFF99299C0",
 -1539 => x"C0C0C0BFF992B090",
 -1538 => x"C0C0C0BFF992B080",
 -1537 => x"C0C0C0BFF992B0F8",
 -1536 => x"C0C0C0BFF992B082",
 -1535 => x"C0C0C0BFF992B092",
 -1534 => x"C0C0C0BFF992B099",
 -1533 => x"C0C0C0BFF992B0B0",
 -1532 => x"C0C0C0BFF992B0A4",
 -1531 => x"C0C0C0BFF992B0F9",
 -1530 => x"C0C0C0BFF992B0C0",
 -1529 => x"C0C0C0BFF992A490",
 -1528 => x"C0C0C0BFF992A480",
 -1527 => x"C0C0C0BFF992A4F8",
 -1526 => x"C0C0C0BFF992A482",
 -1525 => x"C0C0C0BFF992A492",
 -1524 => x"C0C0C0BFF992A499",
 -1523 => x"C0C0C0BFF992A4B0",
 -1522 => x"C0C0C0BFF992A4A4",
 -1521 => x"C0C0C0BFF992A4F9",
 -1520 => x"C0C0C0BFF992A4C0",
 -1519 => x"C0C0C0BFF992F990",
 -1518 => x"C0C0C0BFF992F980",
 -1517 => x"C0C0C0BFF992F9F8",
 -1516 => x"C0C0C0BFF992F982",
 -1515 => x"C0C0C0BFF992F992",
 -1514 => x"C0C0C0BFF992F999",
 -1513 => x"C0C0C0BFF992F9B0",
 -1512 => x"C0C0C0BFF992F9A4",
 -1511 => x"C0C0C0BFF992F9F9",
 -1510 => x"C0C0C0BFF992F9C0",
 -1509 => x"C0C0C0BFF992C090",
 -1508 => x"C0C0C0BFF992C080",
 -1507 => x"C0C0C0BFF992C0F8",
 -1506 => x"C0C0C0BFF992C082",
 -1505 => x"C0C0C0BFF992C092",
 -1504 => x"C0C0C0BFF992C099",
 -1503 => x"C0C0C0BFF992C0B0",
 -1502 => x"C0C0C0BFF992C0A4",
 -1501 => x"C0C0C0BFF992C0F9",
 -1500 => x"C0C0C0BFF992C0C0",
 -1499 => x"C0C0C0BFF9999090",
 -1498 => x"C0C0C0BFF9999080",
 -1497 => x"C0C0C0BFF99990F8",
 -1496 => x"C0C0C0BFF9999082",
 -1495 => x"C0C0C0BFF9999092",
 -1494 => x"C0C0C0BFF9999099",
 -1493 => x"C0C0C0BFF99990B0",
 -1492 => x"C0C0C0BFF99990A4",
 -1491 => x"C0C0C0BFF99990F9",
 -1490 => x"C0C0C0BFF99990C0",
 -1489 => x"C0C0C0BFF9998090",
 -1488 => x"C0C0C0BFF9998080",
 -1487 => x"C0C0C0BFF99980F8",
 -1486 => x"C0C0C0BFF9998082",
 -1485 => x"C0C0C0BFF9998092",
 -1484 => x"C0C0C0BFF9998099",
 -1483 => x"C0C0C0BFF99980B0",
 -1482 => x"C0C0C0BFF99980A4",
 -1481 => x"C0C0C0BFF99980F9",
 -1480 => x"C0C0C0BFF99980C0",
 -1479 => x"C0C0C0BFF999F890",
 -1478 => x"C0C0C0BFF999F880",
 -1477 => x"C0C0C0BFF999F8F8",
 -1476 => x"C0C0C0BFF999F882",
 -1475 => x"C0C0C0BFF999F892",
 -1474 => x"C0C0C0BFF999F899",
 -1473 => x"C0C0C0BFF999F8B0",
 -1472 => x"C0C0C0BFF999F8A4",
 -1471 => x"C0C0C0BFF999F8F9",
 -1470 => x"C0C0C0BFF999F8C0",
 -1469 => x"C0C0C0BFF9998290",
 -1468 => x"C0C0C0BFF9998280",
 -1467 => x"C0C0C0BFF99982F8",
 -1466 => x"C0C0C0BFF9998282",
 -1465 => x"C0C0C0BFF9998292",
 -1464 => x"C0C0C0BFF9998299",
 -1463 => x"C0C0C0BFF99982B0",
 -1462 => x"C0C0C0BFF99982A4",
 -1461 => x"C0C0C0BFF99982F9",
 -1460 => x"C0C0C0BFF99982C0",
 -1459 => x"C0C0C0BFF9999290",
 -1458 => x"C0C0C0BFF9999280",
 -1457 => x"C0C0C0BFF99992F8",
 -1456 => x"C0C0C0BFF9999282",
 -1455 => x"C0C0C0BFF9999292",
 -1454 => x"C0C0C0BFF9999299",
 -1453 => x"C0C0C0BFF99992B0",
 -1452 => x"C0C0C0BFF99992A4",
 -1451 => x"C0C0C0BFF99992F9",
 -1450 => x"C0C0C0BFF99992C0",
 -1449 => x"C0C0C0BFF9999990",
 -1448 => x"C0C0C0BFF9999980",
 -1447 => x"C0C0C0BFF99999F8",
 -1446 => x"C0C0C0BFF9999982",
 -1445 => x"C0C0C0BFF9999992",
 -1444 => x"C0C0C0BFF9999999",
 -1443 => x"C0C0C0BFF99999B0",
 -1442 => x"C0C0C0BFF99999A4",
 -1441 => x"C0C0C0BFF99999F9",
 -1440 => x"C0C0C0BFF99999C0",
 -1439 => x"C0C0C0BFF999B090",
 -1438 => x"C0C0C0BFF999B080",
 -1437 => x"C0C0C0BFF999B0F8",
 -1436 => x"C0C0C0BFF999B082",
 -1435 => x"C0C0C0BFF999B092",
 -1434 => x"C0C0C0BFF999B099",
 -1433 => x"C0C0C0BFF999B0B0",
 -1432 => x"C0C0C0BFF999B0A4",
 -1431 => x"C0C0C0BFF999B0F9",
 -1430 => x"C0C0C0BFF999B0C0",
 -1429 => x"C0C0C0BFF999A490",
 -1428 => x"C0C0C0BFF999A480",
 -1427 => x"C0C0C0BFF999A4F8",
 -1426 => x"C0C0C0BFF999A482",
 -1425 => x"C0C0C0BFF999A492",
 -1424 => x"C0C0C0BFF999A499",
 -1423 => x"C0C0C0BFF999A4B0",
 -1422 => x"C0C0C0BFF999A4A4",
 -1421 => x"C0C0C0BFF999A4F9",
 -1420 => x"C0C0C0BFF999A4C0",
 -1419 => x"C0C0C0BFF999F990",
 -1418 => x"C0C0C0BFF999F980",
 -1417 => x"C0C0C0BFF999F9F8",
 -1416 => x"C0C0C0BFF999F982",
 -1415 => x"C0C0C0BFF999F992",
 -1414 => x"C0C0C0BFF999F999",
 -1413 => x"C0C0C0BFF999F9B0",
 -1412 => x"C0C0C0BFF999F9A4",
 -1411 => x"C0C0C0BFF999F9F9",
 -1410 => x"C0C0C0BFF999F9C0",
 -1409 => x"C0C0C0BFF999C090",
 -1408 => x"C0C0C0BFF999C080",
 -1407 => x"C0C0C0BFF999C0F8",
 -1406 => x"C0C0C0BFF999C082",
 -1405 => x"C0C0C0BFF999C092",
 -1404 => x"C0C0C0BFF999C099",
 -1403 => x"C0C0C0BFF999C0B0",
 -1402 => x"C0C0C0BFF999C0A4",
 -1401 => x"C0C0C0BFF999C0F9",
 -1400 => x"C0C0C0BFF999C0C0",
 -1399 => x"C0C0C0BFF9B09090",
 -1398 => x"C0C0C0BFF9B09080",
 -1397 => x"C0C0C0BFF9B090F8",
 -1396 => x"C0C0C0BFF9B09082",
 -1395 => x"C0C0C0BFF9B09092",
 -1394 => x"C0C0C0BFF9B09099",
 -1393 => x"C0C0C0BFF9B090B0",
 -1392 => x"C0C0C0BFF9B090A4",
 -1391 => x"C0C0C0BFF9B090F9",
 -1390 => x"C0C0C0BFF9B090C0",
 -1389 => x"C0C0C0BFF9B08090",
 -1388 => x"C0C0C0BFF9B08080",
 -1387 => x"C0C0C0BFF9B080F8",
 -1386 => x"C0C0C0BFF9B08082",
 -1385 => x"C0C0C0BFF9B08092",
 -1384 => x"C0C0C0BFF9B08099",
 -1383 => x"C0C0C0BFF9B080B0",
 -1382 => x"C0C0C0BFF9B080A4",
 -1381 => x"C0C0C0BFF9B080F9",
 -1380 => x"C0C0C0BFF9B080C0",
 -1379 => x"C0C0C0BFF9B0F890",
 -1378 => x"C0C0C0BFF9B0F880",
 -1377 => x"C0C0C0BFF9B0F8F8",
 -1376 => x"C0C0C0BFF9B0F882",
 -1375 => x"C0C0C0BFF9B0F892",
 -1374 => x"C0C0C0BFF9B0F899",
 -1373 => x"C0C0C0BFF9B0F8B0",
 -1372 => x"C0C0C0BFF9B0F8A4",
 -1371 => x"C0C0C0BFF9B0F8F9",
 -1370 => x"C0C0C0BFF9B0F8C0",
 -1369 => x"C0C0C0BFF9B08290",
 -1368 => x"C0C0C0BFF9B08280",
 -1367 => x"C0C0C0BFF9B082F8",
 -1366 => x"C0C0C0BFF9B08282",
 -1365 => x"C0C0C0BFF9B08292",
 -1364 => x"C0C0C0BFF9B08299",
 -1363 => x"C0C0C0BFF9B082B0",
 -1362 => x"C0C0C0BFF9B082A4",
 -1361 => x"C0C0C0BFF9B082F9",
 -1360 => x"C0C0C0BFF9B082C0",
 -1359 => x"C0C0C0BFF9B09290",
 -1358 => x"C0C0C0BFF9B09280",
 -1357 => x"C0C0C0BFF9B092F8",
 -1356 => x"C0C0C0BFF9B09282",
 -1355 => x"C0C0C0BFF9B09292",
 -1354 => x"C0C0C0BFF9B09299",
 -1353 => x"C0C0C0BFF9B092B0",
 -1352 => x"C0C0C0BFF9B092A4",
 -1351 => x"C0C0C0BFF9B092F9",
 -1350 => x"C0C0C0BFF9B092C0",
 -1349 => x"C0C0C0BFF9B09990",
 -1348 => x"C0C0C0BFF9B09980",
 -1347 => x"C0C0C0BFF9B099F8",
 -1346 => x"C0C0C0BFF9B09982",
 -1345 => x"C0C0C0BFF9B09992",
 -1344 => x"C0C0C0BFF9B09999",
 -1343 => x"C0C0C0BFF9B099B0",
 -1342 => x"C0C0C0BFF9B099A4",
 -1341 => x"C0C0C0BFF9B099F9",
 -1340 => x"C0C0C0BFF9B099C0",
 -1339 => x"C0C0C0BFF9B0B090",
 -1338 => x"C0C0C0BFF9B0B080",
 -1337 => x"C0C0C0BFF9B0B0F8",
 -1336 => x"C0C0C0BFF9B0B082",
 -1335 => x"C0C0C0BFF9B0B092",
 -1334 => x"C0C0C0BFF9B0B099",
 -1333 => x"C0C0C0BFF9B0B0B0",
 -1332 => x"C0C0C0BFF9B0B0A4",
 -1331 => x"C0C0C0BFF9B0B0F9",
 -1330 => x"C0C0C0BFF9B0B0C0",
 -1329 => x"C0C0C0BFF9B0A490",
 -1328 => x"C0C0C0BFF9B0A480",
 -1327 => x"C0C0C0BFF9B0A4F8",
 -1326 => x"C0C0C0BFF9B0A482",
 -1325 => x"C0C0C0BFF9B0A492",
 -1324 => x"C0C0C0BFF9B0A499",
 -1323 => x"C0C0C0BFF9B0A4B0",
 -1322 => x"C0C0C0BFF9B0A4A4",
 -1321 => x"C0C0C0BFF9B0A4F9",
 -1320 => x"C0C0C0BFF9B0A4C0",
 -1319 => x"C0C0C0BFF9B0F990",
 -1318 => x"C0C0C0BFF9B0F980",
 -1317 => x"C0C0C0BFF9B0F9F8",
 -1316 => x"C0C0C0BFF9B0F982",
 -1315 => x"C0C0C0BFF9B0F992",
 -1314 => x"C0C0C0BFF9B0F999",
 -1313 => x"C0C0C0BFF9B0F9B0",
 -1312 => x"C0C0C0BFF9B0F9A4",
 -1311 => x"C0C0C0BFF9B0F9F9",
 -1310 => x"C0C0C0BFF9B0F9C0",
 -1309 => x"C0C0C0BFF9B0C090",
 -1308 => x"C0C0C0BFF9B0C080",
 -1307 => x"C0C0C0BFF9B0C0F8",
 -1306 => x"C0C0C0BFF9B0C082",
 -1305 => x"C0C0C0BFF9B0C092",
 -1304 => x"C0C0C0BFF9B0C099",
 -1303 => x"C0C0C0BFF9B0C0B0",
 -1302 => x"C0C0C0BFF9B0C0A4",
 -1301 => x"C0C0C0BFF9B0C0F9",
 -1300 => x"C0C0C0BFF9B0C0C0",
 -1299 => x"C0C0C0BFF9A49090",
 -1298 => x"C0C0C0BFF9A49080",
 -1297 => x"C0C0C0BFF9A490F8",
 -1296 => x"C0C0C0BFF9A49082",
 -1295 => x"C0C0C0BFF9A49092",
 -1294 => x"C0C0C0BFF9A49099",
 -1293 => x"C0C0C0BFF9A490B0",
 -1292 => x"C0C0C0BFF9A490A4",
 -1291 => x"C0C0C0BFF9A490F9",
 -1290 => x"C0C0C0BFF9A490C0",
 -1289 => x"C0C0C0BFF9A48090",
 -1288 => x"C0C0C0BFF9A48080",
 -1287 => x"C0C0C0BFF9A480F8",
 -1286 => x"C0C0C0BFF9A48082",
 -1285 => x"C0C0C0BFF9A48092",
 -1284 => x"C0C0C0BFF9A48099",
 -1283 => x"C0C0C0BFF9A480B0",
 -1282 => x"C0C0C0BFF9A480A4",
 -1281 => x"C0C0C0BFF9A480F9",
 -1280 => x"C0C0C0BFF9A480C0",
 -1279 => x"C0C0C0BFF9A4F890",
 -1278 => x"C0C0C0BFF9A4F880",
 -1277 => x"C0C0C0BFF9A4F8F8",
 -1276 => x"C0C0C0BFF9A4F882",
 -1275 => x"C0C0C0BFF9A4F892",
 -1274 => x"C0C0C0BFF9A4F899",
 -1273 => x"C0C0C0BFF9A4F8B0",
 -1272 => x"C0C0C0BFF9A4F8A4",
 -1271 => x"C0C0C0BFF9A4F8F9",
 -1270 => x"C0C0C0BFF9A4F8C0",
 -1269 => x"C0C0C0BFF9A48290",
 -1268 => x"C0C0C0BFF9A48280",
 -1267 => x"C0C0C0BFF9A482F8",
 -1266 => x"C0C0C0BFF9A48282",
 -1265 => x"C0C0C0BFF9A48292",
 -1264 => x"C0C0C0BFF9A48299",
 -1263 => x"C0C0C0BFF9A482B0",
 -1262 => x"C0C0C0BFF9A482A4",
 -1261 => x"C0C0C0BFF9A482F9",
 -1260 => x"C0C0C0BFF9A482C0",
 -1259 => x"C0C0C0BFF9A49290",
 -1258 => x"C0C0C0BFF9A49280",
 -1257 => x"C0C0C0BFF9A492F8",
 -1256 => x"C0C0C0BFF9A49282",
 -1255 => x"C0C0C0BFF9A49292",
 -1254 => x"C0C0C0BFF9A49299",
 -1253 => x"C0C0C0BFF9A492B0",
 -1252 => x"C0C0C0BFF9A492A4",
 -1251 => x"C0C0C0BFF9A492F9",
 -1250 => x"C0C0C0BFF9A492C0",
 -1249 => x"C0C0C0BFF9A49990",
 -1248 => x"C0C0C0BFF9A49980",
 -1247 => x"C0C0C0BFF9A499F8",
 -1246 => x"C0C0C0BFF9A49982",
 -1245 => x"C0C0C0BFF9A49992",
 -1244 => x"C0C0C0BFF9A49999",
 -1243 => x"C0C0C0BFF9A499B0",
 -1242 => x"C0C0C0BFF9A499A4",
 -1241 => x"C0C0C0BFF9A499F9",
 -1240 => x"C0C0C0BFF9A499C0",
 -1239 => x"C0C0C0BFF9A4B090",
 -1238 => x"C0C0C0BFF9A4B080",
 -1237 => x"C0C0C0BFF9A4B0F8",
 -1236 => x"C0C0C0BFF9A4B082",
 -1235 => x"C0C0C0BFF9A4B092",
 -1234 => x"C0C0C0BFF9A4B099",
 -1233 => x"C0C0C0BFF9A4B0B0",
 -1232 => x"C0C0C0BFF9A4B0A4",
 -1231 => x"C0C0C0BFF9A4B0F9",
 -1230 => x"C0C0C0BFF9A4B0C0",
 -1229 => x"C0C0C0BFF9A4A490",
 -1228 => x"C0C0C0BFF9A4A480",
 -1227 => x"C0C0C0BFF9A4A4F8",
 -1226 => x"C0C0C0BFF9A4A482",
 -1225 => x"C0C0C0BFF9A4A492",
 -1224 => x"C0C0C0BFF9A4A499",
 -1223 => x"C0C0C0BFF9A4A4B0",
 -1222 => x"C0C0C0BFF9A4A4A4",
 -1221 => x"C0C0C0BFF9A4A4F9",
 -1220 => x"C0C0C0BFF9A4A4C0",
 -1219 => x"C0C0C0BFF9A4F990",
 -1218 => x"C0C0C0BFF9A4F980",
 -1217 => x"C0C0C0BFF9A4F9F8",
 -1216 => x"C0C0C0BFF9A4F982",
 -1215 => x"C0C0C0BFF9A4F992",
 -1214 => x"C0C0C0BFF9A4F999",
 -1213 => x"C0C0C0BFF9A4F9B0",
 -1212 => x"C0C0C0BFF9A4F9A4",
 -1211 => x"C0C0C0BFF9A4F9F9",
 -1210 => x"C0C0C0BFF9A4F9C0",
 -1209 => x"C0C0C0BFF9A4C090",
 -1208 => x"C0C0C0BFF9A4C080",
 -1207 => x"C0C0C0BFF9A4C0F8",
 -1206 => x"C0C0C0BFF9A4C082",
 -1205 => x"C0C0C0BFF9A4C092",
 -1204 => x"C0C0C0BFF9A4C099",
 -1203 => x"C0C0C0BFF9A4C0B0",
 -1202 => x"C0C0C0BFF9A4C0A4",
 -1201 => x"C0C0C0BFF9A4C0F9",
 -1200 => x"C0C0C0BFF9A4C0C0",
 -1199 => x"C0C0C0BFF9F99090",
 -1198 => x"C0C0C0BFF9F99080",
 -1197 => x"C0C0C0BFF9F990F8",
 -1196 => x"C0C0C0BFF9F99082",
 -1195 => x"C0C0C0BFF9F99092",
 -1194 => x"C0C0C0BFF9F99099",
 -1193 => x"C0C0C0BFF9F990B0",
 -1192 => x"C0C0C0BFF9F990A4",
 -1191 => x"C0C0C0BFF9F990F9",
 -1190 => x"C0C0C0BFF9F990C0",
 -1189 => x"C0C0C0BFF9F98090",
 -1188 => x"C0C0C0BFF9F98080",
 -1187 => x"C0C0C0BFF9F980F8",
 -1186 => x"C0C0C0BFF9F98082",
 -1185 => x"C0C0C0BFF9F98092",
 -1184 => x"C0C0C0BFF9F98099",
 -1183 => x"C0C0C0BFF9F980B0",
 -1182 => x"C0C0C0BFF9F980A4",
 -1181 => x"C0C0C0BFF9F980F9",
 -1180 => x"C0C0C0BFF9F980C0",
 -1179 => x"C0C0C0BFF9F9F890",
 -1178 => x"C0C0C0BFF9F9F880",
 -1177 => x"C0C0C0BFF9F9F8F8",
 -1176 => x"C0C0C0BFF9F9F882",
 -1175 => x"C0C0C0BFF9F9F892",
 -1174 => x"C0C0C0BFF9F9F899",
 -1173 => x"C0C0C0BFF9F9F8B0",
 -1172 => x"C0C0C0BFF9F9F8A4",
 -1171 => x"C0C0C0BFF9F9F8F9",
 -1170 => x"C0C0C0BFF9F9F8C0",
 -1169 => x"C0C0C0BFF9F98290",
 -1168 => x"C0C0C0BFF9F98280",
 -1167 => x"C0C0C0BFF9F982F8",
 -1166 => x"C0C0C0BFF9F98282",
 -1165 => x"C0C0C0BFF9F98292",
 -1164 => x"C0C0C0BFF9F98299",
 -1163 => x"C0C0C0BFF9F982B0",
 -1162 => x"C0C0C0BFF9F982A4",
 -1161 => x"C0C0C0BFF9F982F9",
 -1160 => x"C0C0C0BFF9F982C0",
 -1159 => x"C0C0C0BFF9F99290",
 -1158 => x"C0C0C0BFF9F99280",
 -1157 => x"C0C0C0BFF9F992F8",
 -1156 => x"C0C0C0BFF9F99282",
 -1155 => x"C0C0C0BFF9F99292",
 -1154 => x"C0C0C0BFF9F99299",
 -1153 => x"C0C0C0BFF9F992B0",
 -1152 => x"C0C0C0BFF9F992A4",
 -1151 => x"C0C0C0BFF9F992F9",
 -1150 => x"C0C0C0BFF9F992C0",
 -1149 => x"C0C0C0BFF9F99990",
 -1148 => x"C0C0C0BFF9F99980",
 -1147 => x"C0C0C0BFF9F999F8",
 -1146 => x"C0C0C0BFF9F99982",
 -1145 => x"C0C0C0BFF9F99992",
 -1144 => x"C0C0C0BFF9F99999",
 -1143 => x"C0C0C0BFF9F999B0",
 -1142 => x"C0C0C0BFF9F999A4",
 -1141 => x"C0C0C0BFF9F999F9",
 -1140 => x"C0C0C0BFF9F999C0",
 -1139 => x"C0C0C0BFF9F9B090",
 -1138 => x"C0C0C0BFF9F9B080",
 -1137 => x"C0C0C0BFF9F9B0F8",
 -1136 => x"C0C0C0BFF9F9B082",
 -1135 => x"C0C0C0BFF9F9B092",
 -1134 => x"C0C0C0BFF9F9B099",
 -1133 => x"C0C0C0BFF9F9B0B0",
 -1132 => x"C0C0C0BFF9F9B0A4",
 -1131 => x"C0C0C0BFF9F9B0F9",
 -1130 => x"C0C0C0BFF9F9B0C0",
 -1129 => x"C0C0C0BFF9F9A490",
 -1128 => x"C0C0C0BFF9F9A480",
 -1127 => x"C0C0C0BFF9F9A4F8",
 -1126 => x"C0C0C0BFF9F9A482",
 -1125 => x"C0C0C0BFF9F9A492",
 -1124 => x"C0C0C0BFF9F9A499",
 -1123 => x"C0C0C0BFF9F9A4B0",
 -1122 => x"C0C0C0BFF9F9A4A4",
 -1121 => x"C0C0C0BFF9F9A4F9",
 -1120 => x"C0C0C0BFF9F9A4C0",
 -1119 => x"C0C0C0BFF9F9F990",
 -1118 => x"C0C0C0BFF9F9F980",
 -1117 => x"C0C0C0BFF9F9F9F8",
 -1116 => x"C0C0C0BFF9F9F982",
 -1115 => x"C0C0C0BFF9F9F992",
 -1114 => x"C0C0C0BFF9F9F999",
 -1113 => x"C0C0C0BFF9F9F9B0",
 -1112 => x"C0C0C0BFF9F9F9A4",
 -1111 => x"C0C0C0BFF9F9F9F9",
 -1110 => x"C0C0C0BFF9F9F9C0",
 -1109 => x"C0C0C0BFF9F9C090",
 -1108 => x"C0C0C0BFF9F9C080",
 -1107 => x"C0C0C0BFF9F9C0F8",
 -1106 => x"C0C0C0BFF9F9C082",
 -1105 => x"C0C0C0BFF9F9C092",
 -1104 => x"C0C0C0BFF9F9C099",
 -1103 => x"C0C0C0BFF9F9C0B0",
 -1102 => x"C0C0C0BFF9F9C0A4",
 -1101 => x"C0C0C0BFF9F9C0F9",
 -1100 => x"C0C0C0BFF9F9C0C0",
 -1099 => x"C0C0C0BFF9C09090",
 -1098 => x"C0C0C0BFF9C09080",
 -1097 => x"C0C0C0BFF9C090F8",
 -1096 => x"C0C0C0BFF9C09082",
 -1095 => x"C0C0C0BFF9C09092",
 -1094 => x"C0C0C0BFF9C09099",
 -1093 => x"C0C0C0BFF9C090B0",
 -1092 => x"C0C0C0BFF9C090A4",
 -1091 => x"C0C0C0BFF9C090F9",
 -1090 => x"C0C0C0BFF9C090C0",
 -1089 => x"C0C0C0BFF9C08090",
 -1088 => x"C0C0C0BFF9C08080",
 -1087 => x"C0C0C0BFF9C080F8",
 -1086 => x"C0C0C0BFF9C08082",
 -1085 => x"C0C0C0BFF9C08092",
 -1084 => x"C0C0C0BFF9C08099",
 -1083 => x"C0C0C0BFF9C080B0",
 -1082 => x"C0C0C0BFF9C080A4",
 -1081 => x"C0C0C0BFF9C080F9",
 -1080 => x"C0C0C0BFF9C080C0",
 -1079 => x"C0C0C0BFF9C0F890",
 -1078 => x"C0C0C0BFF9C0F880",
 -1077 => x"C0C0C0BFF9C0F8F8",
 -1076 => x"C0C0C0BFF9C0F882",
 -1075 => x"C0C0C0BFF9C0F892",
 -1074 => x"C0C0C0BFF9C0F899",
 -1073 => x"C0C0C0BFF9C0F8B0",
 -1072 => x"C0C0C0BFF9C0F8A4",
 -1071 => x"C0C0C0BFF9C0F8F9",
 -1070 => x"C0C0C0BFF9C0F8C0",
 -1069 => x"C0C0C0BFF9C08290",
 -1068 => x"C0C0C0BFF9C08280",
 -1067 => x"C0C0C0BFF9C082F8",
 -1066 => x"C0C0C0BFF9C08282",
 -1065 => x"C0C0C0BFF9C08292",
 -1064 => x"C0C0C0BFF9C08299",
 -1063 => x"C0C0C0BFF9C082B0",
 -1062 => x"C0C0C0BFF9C082A4",
 -1061 => x"C0C0C0BFF9C082F9",
 -1060 => x"C0C0C0BFF9C082C0",
 -1059 => x"C0C0C0BFF9C09290",
 -1058 => x"C0C0C0BFF9C09280",
 -1057 => x"C0C0C0BFF9C092F8",
 -1056 => x"C0C0C0BFF9C09282",
 -1055 => x"C0C0C0BFF9C09292",
 -1054 => x"C0C0C0BFF9C09299",
 -1053 => x"C0C0C0BFF9C092B0",
 -1052 => x"C0C0C0BFF9C092A4",
 -1051 => x"C0C0C0BFF9C092F9",
 -1050 => x"C0C0C0BFF9C092C0",
 -1049 => x"C0C0C0BFF9C09990",
 -1048 => x"C0C0C0BFF9C09980",
 -1047 => x"C0C0C0BFF9C099F8",
 -1046 => x"C0C0C0BFF9C09982",
 -1045 => x"C0C0C0BFF9C09992",
 -1044 => x"C0C0C0BFF9C09999",
 -1043 => x"C0C0C0BFF9C099B0",
 -1042 => x"C0C0C0BFF9C099A4",
 -1041 => x"C0C0C0BFF9C099F9",
 -1040 => x"C0C0C0BFF9C099C0",
 -1039 => x"C0C0C0BFF9C0B090",
 -1038 => x"C0C0C0BFF9C0B080",
 -1037 => x"C0C0C0BFF9C0B0F8",
 -1036 => x"C0C0C0BFF9C0B082",
 -1035 => x"C0C0C0BFF9C0B092",
 -1034 => x"C0C0C0BFF9C0B099",
 -1033 => x"C0C0C0BFF9C0B0B0",
 -1032 => x"C0C0C0BFF9C0B0A4",
 -1031 => x"C0C0C0BFF9C0B0F9",
 -1030 => x"C0C0C0BFF9C0B0C0",
 -1029 => x"C0C0C0BFF9C0A490",
 -1028 => x"C0C0C0BFF9C0A480",
 -1027 => x"C0C0C0BFF9C0A4F8",
 -1026 => x"C0C0C0BFF9C0A482",
 -1025 => x"C0C0C0BFF9C0A492",
 -1024 => x"C0C0C0BFF9C0A499",
 -1023 => x"C0C0C0BFF9C0A4B0",
 -1022 => x"C0C0C0BFF9C0A4A4",
 -1021 => x"C0C0C0BFF9C0A4F9",
 -1020 => x"C0C0C0BFF9C0A4C0",
 -1019 => x"C0C0C0BFF9C0F990",
 -1018 => x"C0C0C0BFF9C0F980",
 -1017 => x"C0C0C0BFF9C0F9F8",
 -1016 => x"C0C0C0BFF9C0F982",
 -1015 => x"C0C0C0BFF9C0F992",
 -1014 => x"C0C0C0BFF9C0F999",
 -1013 => x"C0C0C0BFF9C0F9B0",
 -1012 => x"C0C0C0BFF9C0F9A4",
 -1011 => x"C0C0C0BFF9C0F9F9",
 -1010 => x"C0C0C0BFF9C0F9C0",
 -1009 => x"C0C0C0BFF9C0C090",
 -1008 => x"C0C0C0BFF9C0C080",
 -1007 => x"C0C0C0BFF9C0C0F8",
 -1006 => x"C0C0C0BFF9C0C082",
 -1005 => x"C0C0C0BFF9C0C092",
 -1004 => x"C0C0C0BFF9C0C099",
 -1003 => x"C0C0C0BFF9C0C0B0",
 -1002 => x"C0C0C0BFF9C0C0A4",
 -1001 => x"C0C0C0BFF9C0C0F9",
 -1000 => x"C0C0C0BFF9C0C0C0",
  -999 => x"C0C0C0C0BF909090",
  -998 => x"C0C0C0C0BF909080",
  -997 => x"C0C0C0C0BF9090F8",
  -996 => x"C0C0C0C0BF909082",
  -995 => x"C0C0C0C0BF909092",
  -994 => x"C0C0C0C0BF909099",
  -993 => x"C0C0C0C0BF9090B0",
  -992 => x"C0C0C0C0BF9090A4",
  -991 => x"C0C0C0C0BF9090F9",
  -990 => x"C0C0C0C0BF9090C0",
  -989 => x"C0C0C0C0BF908090",
  -988 => x"C0C0C0C0BF908080",
  -987 => x"C0C0C0C0BF9080F8",
  -986 => x"C0C0C0C0BF908082",
  -985 => x"C0C0C0C0BF908092",
  -984 => x"C0C0C0C0BF908099",
  -983 => x"C0C0C0C0BF9080B0",
  -982 => x"C0C0C0C0BF9080A4",
  -981 => x"C0C0C0C0BF9080F9",
  -980 => x"C0C0C0C0BF9080C0",
  -979 => x"C0C0C0C0BF90F890",
  -978 => x"C0C0C0C0BF90F880",
  -977 => x"C0C0C0C0BF90F8F8",
  -976 => x"C0C0C0C0BF90F882",
  -975 => x"C0C0C0C0BF90F892",
  -974 => x"C0C0C0C0BF90F899",
  -973 => x"C0C0C0C0BF90F8B0",
  -972 => x"C0C0C0C0BF90F8A4",
  -971 => x"C0C0C0C0BF90F8F9",
  -970 => x"C0C0C0C0BF90F8C0",
  -969 => x"C0C0C0C0BF908290",
  -968 => x"C0C0C0C0BF908280",
  -967 => x"C0C0C0C0BF9082F8",
  -966 => x"C0C0C0C0BF908282",
  -965 => x"C0C0C0C0BF908292",
  -964 => x"C0C0C0C0BF908299",
  -963 => x"C0C0C0C0BF9082B0",
  -962 => x"C0C0C0C0BF9082A4",
  -961 => x"C0C0C0C0BF9082F9",
  -960 => x"C0C0C0C0BF9082C0",
  -959 => x"C0C0C0C0BF909290",
  -958 => x"C0C0C0C0BF909280",
  -957 => x"C0C0C0C0BF9092F8",
  -956 => x"C0C0C0C0BF909282",
  -955 => x"C0C0C0C0BF909292",
  -954 => x"C0C0C0C0BF909299",
  -953 => x"C0C0C0C0BF9092B0",
  -952 => x"C0C0C0C0BF9092A4",
  -951 => x"C0C0C0C0BF9092F9",
  -950 => x"C0C0C0C0BF9092C0",
  -949 => x"C0C0C0C0BF909990",
  -948 => x"C0C0C0C0BF909980",
  -947 => x"C0C0C0C0BF9099F8",
  -946 => x"C0C0C0C0BF909982",
  -945 => x"C0C0C0C0BF909992",
  -944 => x"C0C0C0C0BF909999",
  -943 => x"C0C0C0C0BF9099B0",
  -942 => x"C0C0C0C0BF9099A4",
  -941 => x"C0C0C0C0BF9099F9",
  -940 => x"C0C0C0C0BF9099C0",
  -939 => x"C0C0C0C0BF90B090",
  -938 => x"C0C0C0C0BF90B080",
  -937 => x"C0C0C0C0BF90B0F8",
  -936 => x"C0C0C0C0BF90B082",
  -935 => x"C0C0C0C0BF90B092",
  -934 => x"C0C0C0C0BF90B099",
  -933 => x"C0C0C0C0BF90B0B0",
  -932 => x"C0C0C0C0BF90B0A4",
  -931 => x"C0C0C0C0BF90B0F9",
  -930 => x"C0C0C0C0BF90B0C0",
  -929 => x"C0C0C0C0BF90A490",
  -928 => x"C0C0C0C0BF90A480",
  -927 => x"C0C0C0C0BF90A4F8",
  -926 => x"C0C0C0C0BF90A482",
  -925 => x"C0C0C0C0BF90A492",
  -924 => x"C0C0C0C0BF90A499",
  -923 => x"C0C0C0C0BF90A4B0",
  -922 => x"C0C0C0C0BF90A4A4",
  -921 => x"C0C0C0C0BF90A4F9",
  -920 => x"C0C0C0C0BF90A4C0",
  -919 => x"C0C0C0C0BF90F990",
  -918 => x"C0C0C0C0BF90F980",
  -917 => x"C0C0C0C0BF90F9F8",
  -916 => x"C0C0C0C0BF90F982",
  -915 => x"C0C0C0C0BF90F992",
  -914 => x"C0C0C0C0BF90F999",
  -913 => x"C0C0C0C0BF90F9B0",
  -912 => x"C0C0C0C0BF90F9A4",
  -911 => x"C0C0C0C0BF90F9F9",
  -910 => x"C0C0C0C0BF90F9C0",
  -909 => x"C0C0C0C0BF90C090",
  -908 => x"C0C0C0C0BF90C080",
  -907 => x"C0C0C0C0BF90C0F8",
  -906 => x"C0C0C0C0BF90C082",
  -905 => x"C0C0C0C0BF90C092",
  -904 => x"C0C0C0C0BF90C099",
  -903 => x"C0C0C0C0BF90C0B0",
  -902 => x"C0C0C0C0BF90C0A4",
  -901 => x"C0C0C0C0BF90C0F9",
  -900 => x"C0C0C0C0BF90C0C0",
  -899 => x"C0C0C0C0BF809090",
  -898 => x"C0C0C0C0BF809080",
  -897 => x"C0C0C0C0BF8090F8",
  -896 => x"C0C0C0C0BF809082",
  -895 => x"C0C0C0C0BF809092",
  -894 => x"C0C0C0C0BF809099",
  -893 => x"C0C0C0C0BF8090B0",
  -892 => x"C0C0C0C0BF8090A4",
  -891 => x"C0C0C0C0BF8090F9",
  -890 => x"C0C0C0C0BF8090C0",
  -889 => x"C0C0C0C0BF808090",
  -888 => x"C0C0C0C0BF808080",
  -887 => x"C0C0C0C0BF8080F8",
  -886 => x"C0C0C0C0BF808082",
  -885 => x"C0C0C0C0BF808092",
  -884 => x"C0C0C0C0BF808099",
  -883 => x"C0C0C0C0BF8080B0",
  -882 => x"C0C0C0C0BF8080A4",
  -881 => x"C0C0C0C0BF8080F9",
  -880 => x"C0C0C0C0BF8080C0",
  -879 => x"C0C0C0C0BF80F890",
  -878 => x"C0C0C0C0BF80F880",
  -877 => x"C0C0C0C0BF80F8F8",
  -876 => x"C0C0C0C0BF80F882",
  -875 => x"C0C0C0C0BF80F892",
  -874 => x"C0C0C0C0BF80F899",
  -873 => x"C0C0C0C0BF80F8B0",
  -872 => x"C0C0C0C0BF80F8A4",
  -871 => x"C0C0C0C0BF80F8F9",
  -870 => x"C0C0C0C0BF80F8C0",
  -869 => x"C0C0C0C0BF808290",
  -868 => x"C0C0C0C0BF808280",
  -867 => x"C0C0C0C0BF8082F8",
  -866 => x"C0C0C0C0BF808282",
  -865 => x"C0C0C0C0BF808292",
  -864 => x"C0C0C0C0BF808299",
  -863 => x"C0C0C0C0BF8082B0",
  -862 => x"C0C0C0C0BF8082A4",
  -861 => x"C0C0C0C0BF8082F9",
  -860 => x"C0C0C0C0BF8082C0",
  -859 => x"C0C0C0C0BF809290",
  -858 => x"C0C0C0C0BF809280",
  -857 => x"C0C0C0C0BF8092F8",
  -856 => x"C0C0C0C0BF809282",
  -855 => x"C0C0C0C0BF809292",
  -854 => x"C0C0C0C0BF809299",
  -853 => x"C0C0C0C0BF8092B0",
  -852 => x"C0C0C0C0BF8092A4",
  -851 => x"C0C0C0C0BF8092F9",
  -850 => x"C0C0C0C0BF8092C0",
  -849 => x"C0C0C0C0BF809990",
  -848 => x"C0C0C0C0BF809980",
  -847 => x"C0C0C0C0BF8099F8",
  -846 => x"C0C0C0C0BF809982",
  -845 => x"C0C0C0C0BF809992",
  -844 => x"C0C0C0C0BF809999",
  -843 => x"C0C0C0C0BF8099B0",
  -842 => x"C0C0C0C0BF8099A4",
  -841 => x"C0C0C0C0BF8099F9",
  -840 => x"C0C0C0C0BF8099C0",
  -839 => x"C0C0C0C0BF80B090",
  -838 => x"C0C0C0C0BF80B080",
  -837 => x"C0C0C0C0BF80B0F8",
  -836 => x"C0C0C0C0BF80B082",
  -835 => x"C0C0C0C0BF80B092",
  -834 => x"C0C0C0C0BF80B099",
  -833 => x"C0C0C0C0BF80B0B0",
  -832 => x"C0C0C0C0BF80B0A4",
  -831 => x"C0C0C0C0BF80B0F9",
  -830 => x"C0C0C0C0BF80B0C0",
  -829 => x"C0C0C0C0BF80A490",
  -828 => x"C0C0C0C0BF80A480",
  -827 => x"C0C0C0C0BF80A4F8",
  -826 => x"C0C0C0C0BF80A482",
  -825 => x"C0C0C0C0BF80A492",
  -824 => x"C0C0C0C0BF80A499",
  -823 => x"C0C0C0C0BF80A4B0",
  -822 => x"C0C0C0C0BF80A4A4",
  -821 => x"C0C0C0C0BF80A4F9",
  -820 => x"C0C0C0C0BF80A4C0",
  -819 => x"C0C0C0C0BF80F990",
  -818 => x"C0C0C0C0BF80F980",
  -817 => x"C0C0C0C0BF80F9F8",
  -816 => x"C0C0C0C0BF80F982",
  -815 => x"C0C0C0C0BF80F992",
  -814 => x"C0C0C0C0BF80F999",
  -813 => x"C0C0C0C0BF80F9B0",
  -812 => x"C0C0C0C0BF80F9A4",
  -811 => x"C0C0C0C0BF80F9F9",
  -810 => x"C0C0C0C0BF80F9C0",
  -809 => x"C0C0C0C0BF80C090",
  -808 => x"C0C0C0C0BF80C080",
  -807 => x"C0C0C0C0BF80C0F8",
  -806 => x"C0C0C0C0BF80C082",
  -805 => x"C0C0C0C0BF80C092",
  -804 => x"C0C0C0C0BF80C099",
  -803 => x"C0C0C0C0BF80C0B0",
  -802 => x"C0C0C0C0BF80C0A4",
  -801 => x"C0C0C0C0BF80C0F9",
  -800 => x"C0C0C0C0BF80C0C0",
  -799 => x"C0C0C0C0BFF89090",
  -798 => x"C0C0C0C0BFF89080",
  -797 => x"C0C0C0C0BFF890F8",
  -796 => x"C0C0C0C0BFF89082",
  -795 => x"C0C0C0C0BFF89092",
  -794 => x"C0C0C0C0BFF89099",
  -793 => x"C0C0C0C0BFF890B0",
  -792 => x"C0C0C0C0BFF890A4",
  -791 => x"C0C0C0C0BFF890F9",
  -790 => x"C0C0C0C0BFF890C0",
  -789 => x"C0C0C0C0BFF88090",
  -788 => x"C0C0C0C0BFF88080",
  -787 => x"C0C0C0C0BFF880F8",
  -786 => x"C0C0C0C0BFF88082",
  -785 => x"C0C0C0C0BFF88092",
  -784 => x"C0C0C0C0BFF88099",
  -783 => x"C0C0C0C0BFF880B0",
  -782 => x"C0C0C0C0BFF880A4",
  -781 => x"C0C0C0C0BFF880F9",
  -780 => x"C0C0C0C0BFF880C0",
  -779 => x"C0C0C0C0BFF8F890",
  -778 => x"C0C0C0C0BFF8F880",
  -777 => x"C0C0C0C0BFF8F8F8",
  -776 => x"C0C0C0C0BFF8F882",
  -775 => x"C0C0C0C0BFF8F892",
  -774 => x"C0C0C0C0BFF8F899",
  -773 => x"C0C0C0C0BFF8F8B0",
  -772 => x"C0C0C0C0BFF8F8A4",
  -771 => x"C0C0C0C0BFF8F8F9",
  -770 => x"C0C0C0C0BFF8F8C0",
  -769 => x"C0C0C0C0BFF88290",
  -768 => x"C0C0C0C0BFF88280",
  -767 => x"C0C0C0C0BFF882F8",
  -766 => x"C0C0C0C0BFF88282",
  -765 => x"C0C0C0C0BFF88292",
  -764 => x"C0C0C0C0BFF88299",
  -763 => x"C0C0C0C0BFF882B0",
  -762 => x"C0C0C0C0BFF882A4",
  -761 => x"C0C0C0C0BFF882F9",
  -760 => x"C0C0C0C0BFF882C0",
  -759 => x"C0C0C0C0BFF89290",
  -758 => x"C0C0C0C0BFF89280",
  -757 => x"C0C0C0C0BFF892F8",
  -756 => x"C0C0C0C0BFF89282",
  -755 => x"C0C0C0C0BFF89292",
  -754 => x"C0C0C0C0BFF89299",
  -753 => x"C0C0C0C0BFF892B0",
  -752 => x"C0C0C0C0BFF892A4",
  -751 => x"C0C0C0C0BFF892F9",
  -750 => x"C0C0C0C0BFF892C0",
  -749 => x"C0C0C0C0BFF89990",
  -748 => x"C0C0C0C0BFF89980",
  -747 => x"C0C0C0C0BFF899F8",
  -746 => x"C0C0C0C0BFF89982",
  -745 => x"C0C0C0C0BFF89992",
  -744 => x"C0C0C0C0BFF89999",
  -743 => x"C0C0C0C0BFF899B0",
  -742 => x"C0C0C0C0BFF899A4",
  -741 => x"C0C0C0C0BFF899F9",
  -740 => x"C0C0C0C0BFF899C0",
  -739 => x"C0C0C0C0BFF8B090",
  -738 => x"C0C0C0C0BFF8B080",
  -737 => x"C0C0C0C0BFF8B0F8",
  -736 => x"C0C0C0C0BFF8B082",
  -735 => x"C0C0C0C0BFF8B092",
  -734 => x"C0C0C0C0BFF8B099",
  -733 => x"C0C0C0C0BFF8B0B0",
  -732 => x"C0C0C0C0BFF8B0A4",
  -731 => x"C0C0C0C0BFF8B0F9",
  -730 => x"C0C0C0C0BFF8B0C0",
  -729 => x"C0C0C0C0BFF8A490",
  -728 => x"C0C0C0C0BFF8A480",
  -727 => x"C0C0C0C0BFF8A4F8",
  -726 => x"C0C0C0C0BFF8A482",
  -725 => x"C0C0C0C0BFF8A492",
  -724 => x"C0C0C0C0BFF8A499",
  -723 => x"C0C0C0C0BFF8A4B0",
  -722 => x"C0C0C0C0BFF8A4A4",
  -721 => x"C0C0C0C0BFF8A4F9",
  -720 => x"C0C0C0C0BFF8A4C0",
  -719 => x"C0C0C0C0BFF8F990",
  -718 => x"C0C0C0C0BFF8F980",
  -717 => x"C0C0C0C0BFF8F9F8",
  -716 => x"C0C0C0C0BFF8F982",
  -715 => x"C0C0C0C0BFF8F992",
  -714 => x"C0C0C0C0BFF8F999",
  -713 => x"C0C0C0C0BFF8F9B0",
  -712 => x"C0C0C0C0BFF8F9A4",
  -711 => x"C0C0C0C0BFF8F9F9",
  -710 => x"C0C0C0C0BFF8F9C0",
  -709 => x"C0C0C0C0BFF8C090",
  -708 => x"C0C0C0C0BFF8C080",
  -707 => x"C0C0C0C0BFF8C0F8",
  -706 => x"C0C0C0C0BFF8C082",
  -705 => x"C0C0C0C0BFF8C092",
  -704 => x"C0C0C0C0BFF8C099",
  -703 => x"C0C0C0C0BFF8C0B0",
  -702 => x"C0C0C0C0BFF8C0A4",
  -701 => x"C0C0C0C0BFF8C0F9",
  -700 => x"C0C0C0C0BFF8C0C0",
  -699 => x"C0C0C0C0BF829090",
  -698 => x"C0C0C0C0BF829080",
  -697 => x"C0C0C0C0BF8290F8",
  -696 => x"C0C0C0C0BF829082",
  -695 => x"C0C0C0C0BF829092",
  -694 => x"C0C0C0C0BF829099",
  -693 => x"C0C0C0C0BF8290B0",
  -692 => x"C0C0C0C0BF8290A4",
  -691 => x"C0C0C0C0BF8290F9",
  -690 => x"C0C0C0C0BF8290C0",
  -689 => x"C0C0C0C0BF828090",
  -688 => x"C0C0C0C0BF828080",
  -687 => x"C0C0C0C0BF8280F8",
  -686 => x"C0C0C0C0BF828082",
  -685 => x"C0C0C0C0BF828092",
  -684 => x"C0C0C0C0BF828099",
  -683 => x"C0C0C0C0BF8280B0",
  -682 => x"C0C0C0C0BF8280A4",
  -681 => x"C0C0C0C0BF8280F9",
  -680 => x"C0C0C0C0BF8280C0",
  -679 => x"C0C0C0C0BF82F890",
  -678 => x"C0C0C0C0BF82F880",
  -677 => x"C0C0C0C0BF82F8F8",
  -676 => x"C0C0C0C0BF82F882",
  -675 => x"C0C0C0C0BF82F892",
  -674 => x"C0C0C0C0BF82F899",
  -673 => x"C0C0C0C0BF82F8B0",
  -672 => x"C0C0C0C0BF82F8A4",
  -671 => x"C0C0C0C0BF82F8F9",
  -670 => x"C0C0C0C0BF82F8C0",
  -669 => x"C0C0C0C0BF828290",
  -668 => x"C0C0C0C0BF828280",
  -667 => x"C0C0C0C0BF8282F8",
  -666 => x"C0C0C0C0BF828282",
  -665 => x"C0C0C0C0BF828292",
  -664 => x"C0C0C0C0BF828299",
  -663 => x"C0C0C0C0BF8282B0",
  -662 => x"C0C0C0C0BF8282A4",
  -661 => x"C0C0C0C0BF8282F9",
  -660 => x"C0C0C0C0BF8282C0",
  -659 => x"C0C0C0C0BF829290",
  -658 => x"C0C0C0C0BF829280",
  -657 => x"C0C0C0C0BF8292F8",
  -656 => x"C0C0C0C0BF829282",
  -655 => x"C0C0C0C0BF829292",
  -654 => x"C0C0C0C0BF829299",
  -653 => x"C0C0C0C0BF8292B0",
  -652 => x"C0C0C0C0BF8292A4",
  -651 => x"C0C0C0C0BF8292F9",
  -650 => x"C0C0C0C0BF8292C0",
  -649 => x"C0C0C0C0BF829990",
  -648 => x"C0C0C0C0BF829980",
  -647 => x"C0C0C0C0BF8299F8",
  -646 => x"C0C0C0C0BF829982",
  -645 => x"C0C0C0C0BF829992",
  -644 => x"C0C0C0C0BF829999",
  -643 => x"C0C0C0C0BF8299B0",
  -642 => x"C0C0C0C0BF8299A4",
  -641 => x"C0C0C0C0BF8299F9",
  -640 => x"C0C0C0C0BF8299C0",
  -639 => x"C0C0C0C0BF82B090",
  -638 => x"C0C0C0C0BF82B080",
  -637 => x"C0C0C0C0BF82B0F8",
  -636 => x"C0C0C0C0BF82B082",
  -635 => x"C0C0C0C0BF82B092",
  -634 => x"C0C0C0C0BF82B099",
  -633 => x"C0C0C0C0BF82B0B0",
  -632 => x"C0C0C0C0BF82B0A4",
  -631 => x"C0C0C0C0BF82B0F9",
  -630 => x"C0C0C0C0BF82B0C0",
  -629 => x"C0C0C0C0BF82A490",
  -628 => x"C0C0C0C0BF82A480",
  -627 => x"C0C0C0C0BF82A4F8",
  -626 => x"C0C0C0C0BF82A482",
  -625 => x"C0C0C0C0BF82A492",
  -624 => x"C0C0C0C0BF82A499",
  -623 => x"C0C0C0C0BF82A4B0",
  -622 => x"C0C0C0C0BF82A4A4",
  -621 => x"C0C0C0C0BF82A4F9",
  -620 => x"C0C0C0C0BF82A4C0",
  -619 => x"C0C0C0C0BF82F990",
  -618 => x"C0C0C0C0BF82F980",
  -617 => x"C0C0C0C0BF82F9F8",
  -616 => x"C0C0C0C0BF82F982",
  -615 => x"C0C0C0C0BF82F992",
  -614 => x"C0C0C0C0BF82F999",
  -613 => x"C0C0C0C0BF82F9B0",
  -612 => x"C0C0C0C0BF82F9A4",
  -611 => x"C0C0C0C0BF82F9F9",
  -610 => x"C0C0C0C0BF82F9C0",
  -609 => x"C0C0C0C0BF82C090",
  -608 => x"C0C0C0C0BF82C080",
  -607 => x"C0C0C0C0BF82C0F8",
  -606 => x"C0C0C0C0BF82C082",
  -605 => x"C0C0C0C0BF82C092",
  -604 => x"C0C0C0C0BF82C099",
  -603 => x"C0C0C0C0BF82C0B0",
  -602 => x"C0C0C0C0BF82C0A4",
  -601 => x"C0C0C0C0BF82C0F9",
  -600 => x"C0C0C0C0BF82C0C0",
  -599 => x"C0C0C0C0BF929090",
  -598 => x"C0C0C0C0BF929080",
  -597 => x"C0C0C0C0BF9290F8",
  -596 => x"C0C0C0C0BF929082",
  -595 => x"C0C0C0C0BF929092",
  -594 => x"C0C0C0C0BF929099",
  -593 => x"C0C0C0C0BF9290B0",
  -592 => x"C0C0C0C0BF9290A4",
  -591 => x"C0C0C0C0BF9290F9",
  -590 => x"C0C0C0C0BF9290C0",
  -589 => x"C0C0C0C0BF928090",
  -588 => x"C0C0C0C0BF928080",
  -587 => x"C0C0C0C0BF9280F8",
  -586 => x"C0C0C0C0BF928082",
  -585 => x"C0C0C0C0BF928092",
  -584 => x"C0C0C0C0BF928099",
  -583 => x"C0C0C0C0BF9280B0",
  -582 => x"C0C0C0C0BF9280A4",
  -581 => x"C0C0C0C0BF9280F9",
  -580 => x"C0C0C0C0BF9280C0",
  -579 => x"C0C0C0C0BF92F890",
  -578 => x"C0C0C0C0BF92F880",
  -577 => x"C0C0C0C0BF92F8F8",
  -576 => x"C0C0C0C0BF92F882",
  -575 => x"C0C0C0C0BF92F892",
  -574 => x"C0C0C0C0BF92F899",
  -573 => x"C0C0C0C0BF92F8B0",
  -572 => x"C0C0C0C0BF92F8A4",
  -571 => x"C0C0C0C0BF92F8F9",
  -570 => x"C0C0C0C0BF92F8C0",
  -569 => x"C0C0C0C0BF928290",
  -568 => x"C0C0C0C0BF928280",
  -567 => x"C0C0C0C0BF9282F8",
  -566 => x"C0C0C0C0BF928282",
  -565 => x"C0C0C0C0BF928292",
  -564 => x"C0C0C0C0BF928299",
  -563 => x"C0C0C0C0BF9282B0",
  -562 => x"C0C0C0C0BF9282A4",
  -561 => x"C0C0C0C0BF9282F9",
  -560 => x"C0C0C0C0BF9282C0",
  -559 => x"C0C0C0C0BF929290",
  -558 => x"C0C0C0C0BF929280",
  -557 => x"C0C0C0C0BF9292F8",
  -556 => x"C0C0C0C0BF929282",
  -555 => x"C0C0C0C0BF929292",
  -554 => x"C0C0C0C0BF929299",
  -553 => x"C0C0C0C0BF9292B0",
  -552 => x"C0C0C0C0BF9292A4",
  -551 => x"C0C0C0C0BF9292F9",
  -550 => x"C0C0C0C0BF9292C0",
  -549 => x"C0C0C0C0BF929990",
  -548 => x"C0C0C0C0BF929980",
  -547 => x"C0C0C0C0BF9299F8",
  -546 => x"C0C0C0C0BF929982",
  -545 => x"C0C0C0C0BF929992",
  -544 => x"C0C0C0C0BF929999",
  -543 => x"C0C0C0C0BF9299B0",
  -542 => x"C0C0C0C0BF9299A4",
  -541 => x"C0C0C0C0BF9299F9",
  -540 => x"C0C0C0C0BF9299C0",
  -539 => x"C0C0C0C0BF92B090",
  -538 => x"C0C0C0C0BF92B080",
  -537 => x"C0C0C0C0BF92B0F8",
  -536 => x"C0C0C0C0BF92B082",
  -535 => x"C0C0C0C0BF92B092",
  -534 => x"C0C0C0C0BF92B099",
  -533 => x"C0C0C0C0BF92B0B0",
  -532 => x"C0C0C0C0BF92B0A4",
  -531 => x"C0C0C0C0BF92B0F9",
  -530 => x"C0C0C0C0BF92B0C0",
  -529 => x"C0C0C0C0BF92A490",
  -528 => x"C0C0C0C0BF92A480",
  -527 => x"C0C0C0C0BF92A4F8",
  -526 => x"C0C0C0C0BF92A482",
  -525 => x"C0C0C0C0BF92A492",
  -524 => x"C0C0C0C0BF92A499",
  -523 => x"C0C0C0C0BF92A4B0",
  -522 => x"C0C0C0C0BF92A4A4",
  -521 => x"C0C0C0C0BF92A4F9",
  -520 => x"C0C0C0C0BF92A4C0",
  -519 => x"C0C0C0C0BF92F990",
  -518 => x"C0C0C0C0BF92F980",
  -517 => x"C0C0C0C0BF92F9F8",
  -516 => x"C0C0C0C0BF92F982",
  -515 => x"C0C0C0C0BF92F992",
  -514 => x"C0C0C0C0BF92F999",
  -513 => x"C0C0C0C0BF92F9B0",
  -512 => x"C0C0C0C0BF92F9A4",
  -511 => x"C0C0C0C0BF92F9F9",
  -510 => x"C0C0C0C0BF92F9C0",
  -509 => x"C0C0C0C0BF92C090",
  -508 => x"C0C0C0C0BF92C080",
  -507 => x"C0C0C0C0BF92C0F8",
  -506 => x"C0C0C0C0BF92C082",
  -505 => x"C0C0C0C0BF92C092",
  -504 => x"C0C0C0C0BF92C099",
  -503 => x"C0C0C0C0BF92C0B0",
  -502 => x"C0C0C0C0BF92C0A4",
  -501 => x"C0C0C0C0BF92C0F9",
  -500 => x"C0C0C0C0BF92C0C0",
  -499 => x"C0C0C0C0BF999090",
  -498 => x"C0C0C0C0BF999080",
  -497 => x"C0C0C0C0BF9990F8",
  -496 => x"C0C0C0C0BF999082",
  -495 => x"C0C0C0C0BF999092",
  -494 => x"C0C0C0C0BF999099",
  -493 => x"C0C0C0C0BF9990B0",
  -492 => x"C0C0C0C0BF9990A4",
  -491 => x"C0C0C0C0BF9990F9",
  -490 => x"C0C0C0C0BF9990C0",
  -489 => x"C0C0C0C0BF998090",
  -488 => x"C0C0C0C0BF998080",
  -487 => x"C0C0C0C0BF9980F8",
  -486 => x"C0C0C0C0BF998082",
  -485 => x"C0C0C0C0BF998092",
  -484 => x"C0C0C0C0BF998099",
  -483 => x"C0C0C0C0BF9980B0",
  -482 => x"C0C0C0C0BF9980A4",
  -481 => x"C0C0C0C0BF9980F9",
  -480 => x"C0C0C0C0BF9980C0",
  -479 => x"C0C0C0C0BF99F890",
  -478 => x"C0C0C0C0BF99F880",
  -477 => x"C0C0C0C0BF99F8F8",
  -476 => x"C0C0C0C0BF99F882",
  -475 => x"C0C0C0C0BF99F892",
  -474 => x"C0C0C0C0BF99F899",
  -473 => x"C0C0C0C0BF99F8B0",
  -472 => x"C0C0C0C0BF99F8A4",
  -471 => x"C0C0C0C0BF99F8F9",
  -470 => x"C0C0C0C0BF99F8C0",
  -469 => x"C0C0C0C0BF998290",
  -468 => x"C0C0C0C0BF998280",
  -467 => x"C0C0C0C0BF9982F8",
  -466 => x"C0C0C0C0BF998282",
  -465 => x"C0C0C0C0BF998292",
  -464 => x"C0C0C0C0BF998299",
  -463 => x"C0C0C0C0BF9982B0",
  -462 => x"C0C0C0C0BF9982A4",
  -461 => x"C0C0C0C0BF9982F9",
  -460 => x"C0C0C0C0BF9982C0",
  -459 => x"C0C0C0C0BF999290",
  -458 => x"C0C0C0C0BF999280",
  -457 => x"C0C0C0C0BF9992F8",
  -456 => x"C0C0C0C0BF999282",
  -455 => x"C0C0C0C0BF999292",
  -454 => x"C0C0C0C0BF999299",
  -453 => x"C0C0C0C0BF9992B0",
  -452 => x"C0C0C0C0BF9992A4",
  -451 => x"C0C0C0C0BF9992F9",
  -450 => x"C0C0C0C0BF9992C0",
  -449 => x"C0C0C0C0BF999990",
  -448 => x"C0C0C0C0BF999980",
  -447 => x"C0C0C0C0BF9999F8",
  -446 => x"C0C0C0C0BF999982",
  -445 => x"C0C0C0C0BF999992",
  -444 => x"C0C0C0C0BF999999",
  -443 => x"C0C0C0C0BF9999B0",
  -442 => x"C0C0C0C0BF9999A4",
  -441 => x"C0C0C0C0BF9999F9",
  -440 => x"C0C0C0C0BF9999C0",
  -439 => x"C0C0C0C0BF99B090",
  -438 => x"C0C0C0C0BF99B080",
  -437 => x"C0C0C0C0BF99B0F8",
  -436 => x"C0C0C0C0BF99B082",
  -435 => x"C0C0C0C0BF99B092",
  -434 => x"C0C0C0C0BF99B099",
  -433 => x"C0C0C0C0BF99B0B0",
  -432 => x"C0C0C0C0BF99B0A4",
  -431 => x"C0C0C0C0BF99B0F9",
  -430 => x"C0C0C0C0BF99B0C0",
  -429 => x"C0C0C0C0BF99A490",
  -428 => x"C0C0C0C0BF99A480",
  -427 => x"C0C0C0C0BF99A4F8",
  -426 => x"C0C0C0C0BF99A482",
  -425 => x"C0C0C0C0BF99A492",
  -424 => x"C0C0C0C0BF99A499",
  -423 => x"C0C0C0C0BF99A4B0",
  -422 => x"C0C0C0C0BF99A4A4",
  -421 => x"C0C0C0C0BF99A4F9",
  -420 => x"C0C0C0C0BF99A4C0",
  -419 => x"C0C0C0C0BF99F990",
  -418 => x"C0C0C0C0BF99F980",
  -417 => x"C0C0C0C0BF99F9F8",
  -416 => x"C0C0C0C0BF99F982",
  -415 => x"C0C0C0C0BF99F992",
  -414 => x"C0C0C0C0BF99F999",
  -413 => x"C0C0C0C0BF99F9B0",
  -412 => x"C0C0C0C0BF99F9A4",
  -411 => x"C0C0C0C0BF99F9F9",
  -410 => x"C0C0C0C0BF99F9C0",
  -409 => x"C0C0C0C0BF99C090",
  -408 => x"C0C0C0C0BF99C080",
  -407 => x"C0C0C0C0BF99C0F8",
  -406 => x"C0C0C0C0BF99C082",
  -405 => x"C0C0C0C0BF99C092",
  -404 => x"C0C0C0C0BF99C099",
  -403 => x"C0C0C0C0BF99C0B0",
  -402 => x"C0C0C0C0BF99C0A4",
  -401 => x"C0C0C0C0BF99C0F9",
  -400 => x"C0C0C0C0BF99C0C0",
  -399 => x"C0C0C0C0BFB09090",
  -398 => x"C0C0C0C0BFB09080",
  -397 => x"C0C0C0C0BFB090F8",
  -396 => x"C0C0C0C0BFB09082",
  -395 => x"C0C0C0C0BFB09092",
  -394 => x"C0C0C0C0BFB09099",
  -393 => x"C0C0C0C0BFB090B0",
  -392 => x"C0C0C0C0BFB090A4",
  -391 => x"C0C0C0C0BFB090F9",
  -390 => x"C0C0C0C0BFB090C0",
  -389 => x"C0C0C0C0BFB08090",
  -388 => x"C0C0C0C0BFB08080",
  -387 => x"C0C0C0C0BFB080F8",
  -386 => x"C0C0C0C0BFB08082",
  -385 => x"C0C0C0C0BFB08092",
  -384 => x"C0C0C0C0BFB08099",
  -383 => x"C0C0C0C0BFB080B0",
  -382 => x"C0C0C0C0BFB080A4",
  -381 => x"C0C0C0C0BFB080F9",
  -380 => x"C0C0C0C0BFB080C0",
  -379 => x"C0C0C0C0BFB0F890",
  -378 => x"C0C0C0C0BFB0F880",
  -377 => x"C0C0C0C0BFB0F8F8",
  -376 => x"C0C0C0C0BFB0F882",
  -375 => x"C0C0C0C0BFB0F892",
  -374 => x"C0C0C0C0BFB0F899",
  -373 => x"C0C0C0C0BFB0F8B0",
  -372 => x"C0C0C0C0BFB0F8A4",
  -371 => x"C0C0C0C0BFB0F8F9",
  -370 => x"C0C0C0C0BFB0F8C0",
  -369 => x"C0C0C0C0BFB08290",
  -368 => x"C0C0C0C0BFB08280",
  -367 => x"C0C0C0C0BFB082F8",
  -366 => x"C0C0C0C0BFB08282",
  -365 => x"C0C0C0C0BFB08292",
  -364 => x"C0C0C0C0BFB08299",
  -363 => x"C0C0C0C0BFB082B0",
  -362 => x"C0C0C0C0BFB082A4",
  -361 => x"C0C0C0C0BFB082F9",
  -360 => x"C0C0C0C0BFB082C0",
  -359 => x"C0C0C0C0BFB09290",
  -358 => x"C0C0C0C0BFB09280",
  -357 => x"C0C0C0C0BFB092F8",
  -356 => x"C0C0C0C0BFB09282",
  -355 => x"C0C0C0C0BFB09292",
  -354 => x"C0C0C0C0BFB09299",
  -353 => x"C0C0C0C0BFB092B0",
  -352 => x"C0C0C0C0BFB092A4",
  -351 => x"C0C0C0C0BFB092F9",
  -350 => x"C0C0C0C0BFB092C0",
  -349 => x"C0C0C0C0BFB09990",
  -348 => x"C0C0C0C0BFB09980",
  -347 => x"C0C0C0C0BFB099F8",
  -346 => x"C0C0C0C0BFB09982",
  -345 => x"C0C0C0C0BFB09992",
  -344 => x"C0C0C0C0BFB09999",
  -343 => x"C0C0C0C0BFB099B0",
  -342 => x"C0C0C0C0BFB099A4",
  -341 => x"C0C0C0C0BFB099F9",
  -340 => x"C0C0C0C0BFB099C0",
  -339 => x"C0C0C0C0BFB0B090",
  -338 => x"C0C0C0C0BFB0B080",
  -337 => x"C0C0C0C0BFB0B0F8",
  -336 => x"C0C0C0C0BFB0B082",
  -335 => x"C0C0C0C0BFB0B092",
  -334 => x"C0C0C0C0BFB0B099",
  -333 => x"C0C0C0C0BFB0B0B0",
  -332 => x"C0C0C0C0BFB0B0A4",
  -331 => x"C0C0C0C0BFB0B0F9",
  -330 => x"C0C0C0C0BFB0B0C0",
  -329 => x"C0C0C0C0BFB0A490",
  -328 => x"C0C0C0C0BFB0A480",
  -327 => x"C0C0C0C0BFB0A4F8",
  -326 => x"C0C0C0C0BFB0A482",
  -325 => x"C0C0C0C0BFB0A492",
  -324 => x"C0C0C0C0BFB0A499",
  -323 => x"C0C0C0C0BFB0A4B0",
  -322 => x"C0C0C0C0BFB0A4A4",
  -321 => x"C0C0C0C0BFB0A4F9",
  -320 => x"C0C0C0C0BFB0A4C0",
  -319 => x"C0C0C0C0BFB0F990",
  -318 => x"C0C0C0C0BFB0F980",
  -317 => x"C0C0C0C0BFB0F9F8",
  -316 => x"C0C0C0C0BFB0F982",
  -315 => x"C0C0C0C0BFB0F992",
  -314 => x"C0C0C0C0BFB0F999",
  -313 => x"C0C0C0C0BFB0F9B0",
  -312 => x"C0C0C0C0BFB0F9A4",
  -311 => x"C0C0C0C0BFB0F9F9",
  -310 => x"C0C0C0C0BFB0F9C0",
  -309 => x"C0C0C0C0BFB0C090",
  -308 => x"C0C0C0C0BFB0C080",
  -307 => x"C0C0C0C0BFB0C0F8",
  -306 => x"C0C0C0C0BFB0C082",
  -305 => x"C0C0C0C0BFB0C092",
  -304 => x"C0C0C0C0BFB0C099",
  -303 => x"C0C0C0C0BFB0C0B0",
  -302 => x"C0C0C0C0BFB0C0A4",
  -301 => x"C0C0C0C0BFB0C0F9",
  -300 => x"C0C0C0C0BFB0C0C0",
  -299 => x"C0C0C0C0BFA49090",
  -298 => x"C0C0C0C0BFA49080",
  -297 => x"C0C0C0C0BFA490F8",
  -296 => x"C0C0C0C0BFA49082",
  -295 => x"C0C0C0C0BFA49092",
  -294 => x"C0C0C0C0BFA49099",
  -293 => x"C0C0C0C0BFA490B0",
  -292 => x"C0C0C0C0BFA490A4",
  -291 => x"C0C0C0C0BFA490F9",
  -290 => x"C0C0C0C0BFA490C0",
  -289 => x"C0C0C0C0BFA48090",
  -288 => x"C0C0C0C0BFA48080",
  -287 => x"C0C0C0C0BFA480F8",
  -286 => x"C0C0C0C0BFA48082",
  -285 => x"C0C0C0C0BFA48092",
  -284 => x"C0C0C0C0BFA48099",
  -283 => x"C0C0C0C0BFA480B0",
  -282 => x"C0C0C0C0BFA480A4",
  -281 => x"C0C0C0C0BFA480F9",
  -280 => x"C0C0C0C0BFA480C0",
  -279 => x"C0C0C0C0BFA4F890",
  -278 => x"C0C0C0C0BFA4F880",
  -277 => x"C0C0C0C0BFA4F8F8",
  -276 => x"C0C0C0C0BFA4F882",
  -275 => x"C0C0C0C0BFA4F892",
  -274 => x"C0C0C0C0BFA4F899",
  -273 => x"C0C0C0C0BFA4F8B0",
  -272 => x"C0C0C0C0BFA4F8A4",
  -271 => x"C0C0C0C0BFA4F8F9",
  -270 => x"C0C0C0C0BFA4F8C0",
  -269 => x"C0C0C0C0BFA48290",
  -268 => x"C0C0C0C0BFA48280",
  -267 => x"C0C0C0C0BFA482F8",
  -266 => x"C0C0C0C0BFA48282",
  -265 => x"C0C0C0C0BFA48292",
  -264 => x"C0C0C0C0BFA48299",
  -263 => x"C0C0C0C0BFA482B0",
  -262 => x"C0C0C0C0BFA482A4",
  -261 => x"C0C0C0C0BFA482F9",
  -260 => x"C0C0C0C0BFA482C0",
  -259 => x"C0C0C0C0BFA49290",
  -258 => x"C0C0C0C0BFA49280",
  -257 => x"C0C0C0C0BFA492F8",
  -256 => x"C0C0C0C0BFA49282",
  -255 => x"C0C0C0C0BFA49292",
  -254 => x"C0C0C0C0BFA49299",
  -253 => x"C0C0C0C0BFA492B0",
  -252 => x"C0C0C0C0BFA492A4",
  -251 => x"C0C0C0C0BFA492F9",
  -250 => x"C0C0C0C0BFA492C0",
  -249 => x"C0C0C0C0BFA49990",
  -248 => x"C0C0C0C0BFA49980",
  -247 => x"C0C0C0C0BFA499F8",
  -246 => x"C0C0C0C0BFA49982",
  -245 => x"C0C0C0C0BFA49992",
  -244 => x"C0C0C0C0BFA49999",
  -243 => x"C0C0C0C0BFA499B0",
  -242 => x"C0C0C0C0BFA499A4",
  -241 => x"C0C0C0C0BFA499F9",
  -240 => x"C0C0C0C0BFA499C0",
  -239 => x"C0C0C0C0BFA4B090",
  -238 => x"C0C0C0C0BFA4B080",
  -237 => x"C0C0C0C0BFA4B0F8",
  -236 => x"C0C0C0C0BFA4B082",
  -235 => x"C0C0C0C0BFA4B092",
  -234 => x"C0C0C0C0BFA4B099",
  -233 => x"C0C0C0C0BFA4B0B0",
  -232 => x"C0C0C0C0BFA4B0A4",
  -231 => x"C0C0C0C0BFA4B0F9",
  -230 => x"C0C0C0C0BFA4B0C0",
  -229 => x"C0C0C0C0BFA4A490",
  -228 => x"C0C0C0C0BFA4A480",
  -227 => x"C0C0C0C0BFA4A4F8",
  -226 => x"C0C0C0C0BFA4A482",
  -225 => x"C0C0C0C0BFA4A492",
  -224 => x"C0C0C0C0BFA4A499",
  -223 => x"C0C0C0C0BFA4A4B0",
  -222 => x"C0C0C0C0BFA4A4A4",
  -221 => x"C0C0C0C0BFA4A4F9",
  -220 => x"C0C0C0C0BFA4A4C0",
  -219 => x"C0C0C0C0BFA4F990",
  -218 => x"C0C0C0C0BFA4F980",
  -217 => x"C0C0C0C0BFA4F9F8",
  -216 => x"C0C0C0C0BFA4F982",
  -215 => x"C0C0C0C0BFA4F992",
  -214 => x"C0C0C0C0BFA4F999",
  -213 => x"C0C0C0C0BFA4F9B0",
  -212 => x"C0C0C0C0BFA4F9A4",
  -211 => x"C0C0C0C0BFA4F9F9",
  -210 => x"C0C0C0C0BFA4F9C0",
  -209 => x"C0C0C0C0BFA4C090",
  -208 => x"C0C0C0C0BFA4C080",
  -207 => x"C0C0C0C0BFA4C0F8",
  -206 => x"C0C0C0C0BFA4C082",
  -205 => x"C0C0C0C0BFA4C092",
  -204 => x"C0C0C0C0BFA4C099",
  -203 => x"C0C0C0C0BFA4C0B0",
  -202 => x"C0C0C0C0BFA4C0A4",
  -201 => x"C0C0C0C0BFA4C0F9",
  -200 => x"C0C0C0C0BFA4C0C0",
  -199 => x"C0C0C0C0BFF99090",
  -198 => x"C0C0C0C0BFF99080",
  -197 => x"C0C0C0C0BFF990F8",
  -196 => x"C0C0C0C0BFF99082",
  -195 => x"C0C0C0C0BFF99092",
  -194 => x"C0C0C0C0BFF99099",
  -193 => x"C0C0C0C0BFF990B0",
  -192 => x"C0C0C0C0BFF990A4",
  -191 => x"C0C0C0C0BFF990F9",
  -190 => x"C0C0C0C0BFF990C0",
  -189 => x"C0C0C0C0BFF98090",
  -188 => x"C0C0C0C0BFF98080",
  -187 => x"C0C0C0C0BFF980F8",
  -186 => x"C0C0C0C0BFF98082",
  -185 => x"C0C0C0C0BFF98092",
  -184 => x"C0C0C0C0BFF98099",
  -183 => x"C0C0C0C0BFF980B0",
  -182 => x"C0C0C0C0BFF980A4",
  -181 => x"C0C0C0C0BFF980F9",
  -180 => x"C0C0C0C0BFF980C0",
  -179 => x"C0C0C0C0BFF9F890",
  -178 => x"C0C0C0C0BFF9F880",
  -177 => x"C0C0C0C0BFF9F8F8",
  -176 => x"C0C0C0C0BFF9F882",
  -175 => x"C0C0C0C0BFF9F892",
  -174 => x"C0C0C0C0BFF9F899",
  -173 => x"C0C0C0C0BFF9F8B0",
  -172 => x"C0C0C0C0BFF9F8A4",
  -171 => x"C0C0C0C0BFF9F8F9",
  -170 => x"C0C0C0C0BFF9F8C0",
  -169 => x"C0C0C0C0BFF98290",
  -168 => x"C0C0C0C0BFF98280",
  -167 => x"C0C0C0C0BFF982F8",
  -166 => x"C0C0C0C0BFF98282",
  -165 => x"C0C0C0C0BFF98292",
  -164 => x"C0C0C0C0BFF98299",
  -163 => x"C0C0C0C0BFF982B0",
  -162 => x"C0C0C0C0BFF982A4",
  -161 => x"C0C0C0C0BFF982F9",
  -160 => x"C0C0C0C0BFF982C0",
  -159 => x"C0C0C0C0BFF99290",
  -158 => x"C0C0C0C0BFF99280",
  -157 => x"C0C0C0C0BFF992F8",
  -156 => x"C0C0C0C0BFF99282",
  -155 => x"C0C0C0C0BFF99292",
  -154 => x"C0C0C0C0BFF99299",
  -153 => x"C0C0C0C0BFF992B0",
  -152 => x"C0C0C0C0BFF992A4",
  -151 => x"C0C0C0C0BFF992F9",
  -150 => x"C0C0C0C0BFF992C0",
  -149 => x"C0C0C0C0BFF99990",
  -148 => x"C0C0C0C0BFF99980",
  -147 => x"C0C0C0C0BFF999F8",
  -146 => x"C0C0C0C0BFF99982",
  -145 => x"C0C0C0C0BFF99992",
  -144 => x"C0C0C0C0BFF99999",
  -143 => x"C0C0C0C0BFF999B0",
  -142 => x"C0C0C0C0BFF999A4",
  -141 => x"C0C0C0C0BFF999F9",
  -140 => x"C0C0C0C0BFF999C0",
  -139 => x"C0C0C0C0BFF9B090",
  -138 => x"C0C0C0C0BFF9B080",
  -137 => x"C0C0C0C0BFF9B0F8",
  -136 => x"C0C0C0C0BFF9B082",
  -135 => x"C0C0C0C0BFF9B092",
  -134 => x"C0C0C0C0BFF9B099",
  -133 => x"C0C0C0C0BFF9B0B0",
  -132 => x"C0C0C0C0BFF9B0A4",
  -131 => x"C0C0C0C0BFF9B0F9",
  -130 => x"C0C0C0C0BFF9B0C0",
  -129 => x"C0C0C0C0BFF9A490",
  -128 => x"C0C0C0C0BFF9A480",
  -127 => x"C0C0C0C0BFF9A4F8",
  -126 => x"C0C0C0C0BFF9A482",
  -125 => x"C0C0C0C0BFF9A492",
  -124 => x"C0C0C0C0BFF9A499",
  -123 => x"C0C0C0C0BFF9A4B0",
  -122 => x"C0C0C0C0BFF9A4A4",
  -121 => x"C0C0C0C0BFF9A4F9",
  -120 => x"C0C0C0C0BFF9A4C0",
  -119 => x"C0C0C0C0BFF9F990",
  -118 => x"C0C0C0C0BFF9F980",
  -117 => x"C0C0C0C0BFF9F9F8",
  -116 => x"C0C0C0C0BFF9F982",
  -115 => x"C0C0C0C0BFF9F992",
  -114 => x"C0C0C0C0BFF9F999",
  -113 => x"C0C0C0C0BFF9F9B0",
  -112 => x"C0C0C0C0BFF9F9A4",
  -111 => x"C0C0C0C0BFF9F9F9",
  -110 => x"C0C0C0C0BFF9F9C0",
  -109 => x"C0C0C0C0BFF9C090",
  -108 => x"C0C0C0C0BFF9C080",
  -107 => x"C0C0C0C0BFF9C0F8",
  -106 => x"C0C0C0C0BFF9C082",
  -105 => x"C0C0C0C0BFF9C092",
  -104 => x"C0C0C0C0BFF9C099",
  -103 => x"C0C0C0C0BFF9C0B0",
  -102 => x"C0C0C0C0BFF9C0A4",
  -101 => x"C0C0C0C0BFF9C0F9",
  -100 => x"C0C0C0C0BFF9C0C0",
   -99 => x"C0C0C0C0C0BF9090",
   -98 => x"C0C0C0C0C0BF9080",
   -97 => x"C0C0C0C0C0BF90F8",
   -96 => x"C0C0C0C0C0BF9082",
   -95 => x"C0C0C0C0C0BF9092",
   -94 => x"C0C0C0C0C0BF9099",
   -93 => x"C0C0C0C0C0BF90B0",
   -92 => x"C0C0C0C0C0BF90A4",
   -91 => x"C0C0C0C0C0BF90F9",
   -90 => x"C0C0C0C0C0BF90C0",
   -89 => x"C0C0C0C0C0BF8090",
   -88 => x"C0C0C0C0C0BF8080",
   -87 => x"C0C0C0C0C0BF80F8",
   -86 => x"C0C0C0C0C0BF8082",
   -85 => x"C0C0C0C0C0BF8092",
   -84 => x"C0C0C0C0C0BF8099",
   -83 => x"C0C0C0C0C0BF80B0",
   -82 => x"C0C0C0C0C0BF80A4",
   -81 => x"C0C0C0C0C0BF80F9",
   -80 => x"C0C0C0C0C0BF80C0",
   -79 => x"C0C0C0C0C0BFF890",
   -78 => x"C0C0C0C0C0BFF880",
   -77 => x"C0C0C0C0C0BFF8F8",
   -76 => x"C0C0C0C0C0BFF882",
   -75 => x"C0C0C0C0C0BFF892",
   -74 => x"C0C0C0C0C0BFF899",
   -73 => x"C0C0C0C0C0BFF8B0",
   -72 => x"C0C0C0C0C0BFF8A4",
   -71 => x"C0C0C0C0C0BFF8F9",
   -70 => x"C0C0C0C0C0BFF8C0",
   -69 => x"C0C0C0C0C0BF8290",
   -68 => x"C0C0C0C0C0BF8280",
   -67 => x"C0C0C0C0C0BF82F8",
   -66 => x"C0C0C0C0C0BF8282",
   -65 => x"C0C0C0C0C0BF8292",
   -64 => x"C0C0C0C0C0BF8299",
   -63 => x"C0C0C0C0C0BF82B0",
   -62 => x"C0C0C0C0C0BF82A4",
   -61 => x"C0C0C0C0C0BF82F9",
   -60 => x"C0C0C0C0C0BF82C0",
   -59 => x"C0C0C0C0C0BF9290",
   -58 => x"C0C0C0C0C0BF9280",
   -57 => x"C0C0C0C0C0BF92F8",
   -56 => x"C0C0C0C0C0BF9282",
   -55 => x"C0C0C0C0C0BF9292",
   -54 => x"C0C0C0C0C0BF9299",
   -53 => x"C0C0C0C0C0BF92B0",
   -52 => x"C0C0C0C0C0BF92A4",
   -51 => x"C0C0C0C0C0BF92F9",
   -50 => x"C0C0C0C0C0BF92C0",
   -49 => x"C0C0C0C0C0BF9990",
   -48 => x"C0C0C0C0C0BF9980",
   -47 => x"C0C0C0C0C0BF99F8",
   -46 => x"C0C0C0C0C0BF9982",
   -45 => x"C0C0C0C0C0BF9992",
   -44 => x"C0C0C0C0C0BF9999",
   -43 => x"C0C0C0C0C0BF99B0",
   -42 => x"C0C0C0C0C0BF99A4",
   -41 => x"C0C0C0C0C0BF99F9",
   -40 => x"C0C0C0C0C0BF99C0",
   -39 => x"C0C0C0C0C0BFB090",
   -38 => x"C0C0C0C0C0BFB080",
   -37 => x"C0C0C0C0C0BFB0F8",
   -36 => x"C0C0C0C0C0BFB082",
   -35 => x"C0C0C0C0C0BFB092",
   -34 => x"C0C0C0C0C0BFB099",
   -33 => x"C0C0C0C0C0BFB0B0",
   -32 => x"C0C0C0C0C0BFB0A4",
   -31 => x"C0C0C0C0C0BFB0F9",
   -30 => x"C0C0C0C0C0BFB0C0",
   -29 => x"C0C0C0C0C0BFA490",
   -28 => x"C0C0C0C0C0BFA480",
   -27 => x"C0C0C0C0C0BFA4F8",
   -26 => x"C0C0C0C0C0BFA482",
   -25 => x"C0C0C0C0C0BFA492",
   -24 => x"C0C0C0C0C0BFA499",
   -23 => x"C0C0C0C0C0BFA4B0",
   -22 => x"C0C0C0C0C0BFA4A4",
   -21 => x"C0C0C0C0C0BFA4F9",
   -20 => x"C0C0C0C0C0BFA4C0",
   -19 => x"C0C0C0C0C0BFF990",
   -18 => x"C0C0C0C0C0BFF980",
   -17 => x"C0C0C0C0C0BFF9F8",
   -16 => x"C0C0C0C0C0BFF982",
   -15 => x"C0C0C0C0C0BFF992",
   -14 => x"C0C0C0C0C0BFF999",
   -13 => x"C0C0C0C0C0BFF9B0",
   -12 => x"C0C0C0C0C0BFF9A4",
   -11 => x"C0C0C0C0C0BFF9F9",
   -10 => x"C0C0C0C0C0BFF9C0",
    -9 => x"C0C0C0C0C0C0BF90",
    -8 => x"C0C0C0C0C0C0BF80",
    -7 => x"C0C0C0C0C0C0BFF8",
    -6 => x"C0C0C0C0C0C0BF82",
    -5 => x"C0C0C0C0C0C0BF92",
    -4 => x"C0C0C0C0C0C0BF99",
    -3 => x"C0C0C0C0C0C0BFB0",
    -2 => x"C0C0C0C0C0C0BFA4",
    -1 => x"C0C0C0C0C0C0BFF9",
     0 => x"C0C0C0C0C0C0C0C0",
     1 => x"C0C0C0C0C0C0C0F9",
     2 => x"C0C0C0C0C0C0C0A4",
     3 => x"C0C0C0C0C0C0C0B0",
     4 => x"C0C0C0C0C0C0C099",
     5 => x"C0C0C0C0C0C0C092",
     6 => x"C0C0C0C0C0C0C082",
     7 => x"C0C0C0C0C0C0C0F8",
     8 => x"C0C0C0C0C0C0C080",
     9 => x"C0C0C0C0C0C0C090",
    10 => x"C0C0C0C0C0C0F9C0",
    11 => x"C0C0C0C0C0C0F9F9",
    12 => x"C0C0C0C0C0C0F9A4",
    13 => x"C0C0C0C0C0C0F9B0",
    14 => x"C0C0C0C0C0C0F999",
    15 => x"C0C0C0C0C0C0F992",
    16 => x"C0C0C0C0C0C0F982",
    17 => x"C0C0C0C0C0C0F9F8",
    18 => x"C0C0C0C0C0C0F980",
    19 => x"C0C0C0C0C0C0F990",
    20 => x"C0C0C0C0C0C0A4C0",
    21 => x"C0C0C0C0C0C0A4F9",
    22 => x"C0C0C0C0C0C0A4A4",
    23 => x"C0C0C0C0C0C0A4B0",
    24 => x"C0C0C0C0C0C0A499",
    25 => x"C0C0C0C0C0C0A492",
    26 => x"C0C0C0C0C0C0A482",
    27 => x"C0C0C0C0C0C0A4F8",
    28 => x"C0C0C0C0C0C0A480",
    29 => x"C0C0C0C0C0C0A490",
    30 => x"C0C0C0C0C0C0B0C0",
    31 => x"C0C0C0C0C0C0B0F9",
    32 => x"C0C0C0C0C0C0B0A4",
    33 => x"C0C0C0C0C0C0B0B0",
    34 => x"C0C0C0C0C0C0B099",
    35 => x"C0C0C0C0C0C0B092",
    36 => x"C0C0C0C0C0C0B082",
    37 => x"C0C0C0C0C0C0B0F8",
    38 => x"C0C0C0C0C0C0B080",
    39 => x"C0C0C0C0C0C0B090",
    40 => x"C0C0C0C0C0C099C0",
    41 => x"C0C0C0C0C0C099F9",
    42 => x"C0C0C0C0C0C099A4",
    43 => x"C0C0C0C0C0C099B0",
    44 => x"C0C0C0C0C0C09999",
    45 => x"C0C0C0C0C0C09992",
    46 => x"C0C0C0C0C0C09982",
    47 => x"C0C0C0C0C0C099F8",
    48 => x"C0C0C0C0C0C09980",
    49 => x"C0C0C0C0C0C09990",
    50 => x"C0C0C0C0C0C092C0",
    51 => x"C0C0C0C0C0C092F9",
    52 => x"C0C0C0C0C0C092A4",
    53 => x"C0C0C0C0C0C092B0",
    54 => x"C0C0C0C0C0C09299",
    55 => x"C0C0C0C0C0C09292",
    56 => x"C0C0C0C0C0C09282",
    57 => x"C0C0C0C0C0C092F8",
    58 => x"C0C0C0C0C0C09280",
    59 => x"C0C0C0C0C0C09290",
    60 => x"C0C0C0C0C0C082C0",
    61 => x"C0C0C0C0C0C082F9",
    62 => x"C0C0C0C0C0C082A4",
    63 => x"C0C0C0C0C0C082B0",
    64 => x"C0C0C0C0C0C08299",
    65 => x"C0C0C0C0C0C08292",
    66 => x"C0C0C0C0C0C08282",
    67 => x"C0C0C0C0C0C082F8",
    68 => x"C0C0C0C0C0C08280",
    69 => x"C0C0C0C0C0C08290",
    70 => x"C0C0C0C0C0C0F8C0",
    71 => x"C0C0C0C0C0C0F8F9",
    72 => x"C0C0C0C0C0C0F8A4",
    73 => x"C0C0C0C0C0C0F8B0",
    74 => x"C0C0C0C0C0C0F899",
    75 => x"C0C0C0C0C0C0F892",
    76 => x"C0C0C0C0C0C0F882",
    77 => x"C0C0C0C0C0C0F8F8",
    78 => x"C0C0C0C0C0C0F880",
    79 => x"C0C0C0C0C0C0F890",
    80 => x"C0C0C0C0C0C080C0",
    81 => x"C0C0C0C0C0C080F9",
    82 => x"C0C0C0C0C0C080A4",
    83 => x"C0C0C0C0C0C080B0",
    84 => x"C0C0C0C0C0C08099",
    85 => x"C0C0C0C0C0C08092",
    86 => x"C0C0C0C0C0C08082",
    87 => x"C0C0C0C0C0C080F8",
    88 => x"C0C0C0C0C0C08080",
    89 => x"C0C0C0C0C0C08090",
    90 => x"C0C0C0C0C0C090C0",
    91 => x"C0C0C0C0C0C090F9",
    92 => x"C0C0C0C0C0C090A4",
    93 => x"C0C0C0C0C0C090B0",
    94 => x"C0C0C0C0C0C09099",
    95 => x"C0C0C0C0C0C09092",
    96 => x"C0C0C0C0C0C09082",
    97 => x"C0C0C0C0C0C090F8",
    98 => x"C0C0C0C0C0C09080",
    99 => x"C0C0C0C0C0C09090",
   100 => x"C0C0C0C0C0F9C0C0",
   101 => x"C0C0C0C0C0F9C0F9",
   102 => x"C0C0C0C0C0F9C0A4",
   103 => x"C0C0C0C0C0F9C0B0",
   104 => x"C0C0C0C0C0F9C099",
   105 => x"C0C0C0C0C0F9C092",
   106 => x"C0C0C0C0C0F9C082",
   107 => x"C0C0C0C0C0F9C0F8",
   108 => x"C0C0C0C0C0F9C080",
   109 => x"C0C0C0C0C0F9C090",
   110 => x"C0C0C0C0C0F9F9C0",
   111 => x"C0C0C0C0C0F9F9F9",
   112 => x"C0C0C0C0C0F9F9A4",
   113 => x"C0C0C0C0C0F9F9B0",
   114 => x"C0C0C0C0C0F9F999",
   115 => x"C0C0C0C0C0F9F992",
   116 => x"C0C0C0C0C0F9F982",
   117 => x"C0C0C0C0C0F9F9F8",
   118 => x"C0C0C0C0C0F9F980",
   119 => x"C0C0C0C0C0F9F990",
   120 => x"C0C0C0C0C0F9A4C0",
   121 => x"C0C0C0C0C0F9A4F9",
   122 => x"C0C0C0C0C0F9A4A4",
   123 => x"C0C0C0C0C0F9A4B0",
   124 => x"C0C0C0C0C0F9A499",
   125 => x"C0C0C0C0C0F9A492",
   126 => x"C0C0C0C0C0F9A482",
   127 => x"C0C0C0C0C0F9A4F8",
   128 => x"C0C0C0C0C0F9A480",
   129 => x"C0C0C0C0C0F9A490",
   130 => x"C0C0C0C0C0F9B0C0",
   131 => x"C0C0C0C0C0F9B0F9",
   132 => x"C0C0C0C0C0F9B0A4",
   133 => x"C0C0C0C0C0F9B0B0",
   134 => x"C0C0C0C0C0F9B099",
   135 => x"C0C0C0C0C0F9B092",
   136 => x"C0C0C0C0C0F9B082",
   137 => x"C0C0C0C0C0F9B0F8",
   138 => x"C0C0C0C0C0F9B080",
   139 => x"C0C0C0C0C0F9B090",
   140 => x"C0C0C0C0C0F999C0",
   141 => x"C0C0C0C0C0F999F9",
   142 => x"C0C0C0C0C0F999A4",
   143 => x"C0C0C0C0C0F999B0",
   144 => x"C0C0C0C0C0F99999",
   145 => x"C0C0C0C0C0F99992",
   146 => x"C0C0C0C0C0F99982",
   147 => x"C0C0C0C0C0F999F8",
   148 => x"C0C0C0C0C0F99980",
   149 => x"C0C0C0C0C0F99990",
   150 => x"C0C0C0C0C0F992C0",
   151 => x"C0C0C0C0C0F992F9",
   152 => x"C0C0C0C0C0F992A4",
   153 => x"C0C0C0C0C0F992B0",
   154 => x"C0C0C0C0C0F99299",
   155 => x"C0C0C0C0C0F99292",
   156 => x"C0C0C0C0C0F99282",
   157 => x"C0C0C0C0C0F992F8",
   158 => x"C0C0C0C0C0F99280",
   159 => x"C0C0C0C0C0F99290",
   160 => x"C0C0C0C0C0F982C0",
   161 => x"C0C0C0C0C0F982F9",
   162 => x"C0C0C0C0C0F982A4",
   163 => x"C0C0C0C0C0F982B0",
   164 => x"C0C0C0C0C0F98299",
   165 => x"C0C0C0C0C0F98292",
   166 => x"C0C0C0C0C0F98282",
   167 => x"C0C0C0C0C0F982F8",
   168 => x"C0C0C0C0C0F98280",
   169 => x"C0C0C0C0C0F98290",
   170 => x"C0C0C0C0C0F9F8C0",
   171 => x"C0C0C0C0C0F9F8F9",
   172 => x"C0C0C0C0C0F9F8A4",
   173 => x"C0C0C0C0C0F9F8B0",
   174 => x"C0C0C0C0C0F9F899",
   175 => x"C0C0C0C0C0F9F892",
   176 => x"C0C0C0C0C0F9F882",
   177 => x"C0C0C0C0C0F9F8F8",
   178 => x"C0C0C0C0C0F9F880",
   179 => x"C0C0C0C0C0F9F890",
   180 => x"C0C0C0C0C0F980C0",
   181 => x"C0C0C0C0C0F980F9",
   182 => x"C0C0C0C0C0F980A4",
   183 => x"C0C0C0C0C0F980B0",
   184 => x"C0C0C0C0C0F98099",
   185 => x"C0C0C0C0C0F98092",
   186 => x"C0C0C0C0C0F98082",
   187 => x"C0C0C0C0C0F980F8",
   188 => x"C0C0C0C0C0F98080",
   189 => x"C0C0C0C0C0F98090",
   190 => x"C0C0C0C0C0F990C0",
   191 => x"C0C0C0C0C0F990F9",
   192 => x"C0C0C0C0C0F990A4",
   193 => x"C0C0C0C0C0F990B0",
   194 => x"C0C0C0C0C0F99099",
   195 => x"C0C0C0C0C0F99092",
   196 => x"C0C0C0C0C0F99082",
   197 => x"C0C0C0C0C0F990F8",
   198 => x"C0C0C0C0C0F99080",
   199 => x"C0C0C0C0C0F99090",
   200 => x"C0C0C0C0C0A4C0C0",
   201 => x"C0C0C0C0C0A4C0F9",
   202 => x"C0C0C0C0C0A4C0A4",
   203 => x"C0C0C0C0C0A4C0B0",
   204 => x"C0C0C0C0C0A4C099",
   205 => x"C0C0C0C0C0A4C092",
   206 => x"C0C0C0C0C0A4C082",
   207 => x"C0C0C0C0C0A4C0F8",
   208 => x"C0C0C0C0C0A4C080",
   209 => x"C0C0C0C0C0A4C090",
   210 => x"C0C0C0C0C0A4F9C0",
   211 => x"C0C0C0C0C0A4F9F9",
   212 => x"C0C0C0C0C0A4F9A4",
   213 => x"C0C0C0C0C0A4F9B0",
   214 => x"C0C0C0C0C0A4F999",
   215 => x"C0C0C0C0C0A4F992",
   216 => x"C0C0C0C0C0A4F982",
   217 => x"C0C0C0C0C0A4F9F8",
   218 => x"C0C0C0C0C0A4F980",
   219 => x"C0C0C0C0C0A4F990",
   220 => x"C0C0C0C0C0A4A4C0",
   221 => x"C0C0C0C0C0A4A4F9",
   222 => x"C0C0C0C0C0A4A4A4",
   223 => x"C0C0C0C0C0A4A4B0",
   224 => x"C0C0C0C0C0A4A499",
   225 => x"C0C0C0C0C0A4A492",
   226 => x"C0C0C0C0C0A4A482",
   227 => x"C0C0C0C0C0A4A4F8",
   228 => x"C0C0C0C0C0A4A480",
   229 => x"C0C0C0C0C0A4A490",
   230 => x"C0C0C0C0C0A4B0C0",
   231 => x"C0C0C0C0C0A4B0F9",
   232 => x"C0C0C0C0C0A4B0A4",
   233 => x"C0C0C0C0C0A4B0B0",
   234 => x"C0C0C0C0C0A4B099",
   235 => x"C0C0C0C0C0A4B092",
   236 => x"C0C0C0C0C0A4B082",
   237 => x"C0C0C0C0C0A4B0F8",
   238 => x"C0C0C0C0C0A4B080",
   239 => x"C0C0C0C0C0A4B090",
   240 => x"C0C0C0C0C0A499C0",
   241 => x"C0C0C0C0C0A499F9",
   242 => x"C0C0C0C0C0A499A4",
   243 => x"C0C0C0C0C0A499B0",
   244 => x"C0C0C0C0C0A49999",
   245 => x"C0C0C0C0C0A49992",
   246 => x"C0C0C0C0C0A49982",
   247 => x"C0C0C0C0C0A499F8",
   248 => x"C0C0C0C0C0A49980",
   249 => x"C0C0C0C0C0A49990",
   250 => x"C0C0C0C0C0A492C0",
   251 => x"C0C0C0C0C0A492F9",
   252 => x"C0C0C0C0C0A492A4",
   253 => x"C0C0C0C0C0A492B0",
   254 => x"C0C0C0C0C0A49299",
   255 => x"C0C0C0C0C0A49292",
   256 => x"C0C0C0C0C0A49282",
   257 => x"C0C0C0C0C0A492F8",
   258 => x"C0C0C0C0C0A49280",
   259 => x"C0C0C0C0C0A49290",
   260 => x"C0C0C0C0C0A482C0",
   261 => x"C0C0C0C0C0A482F9",
   262 => x"C0C0C0C0C0A482A4",
   263 => x"C0C0C0C0C0A482B0",
   264 => x"C0C0C0C0C0A48299",
   265 => x"C0C0C0C0C0A48292",
   266 => x"C0C0C0C0C0A48282",
   267 => x"C0C0C0C0C0A482F8",
   268 => x"C0C0C0C0C0A48280",
   269 => x"C0C0C0C0C0A48290",
   270 => x"C0C0C0C0C0A4F8C0",
   271 => x"C0C0C0C0C0A4F8F9",
   272 => x"C0C0C0C0C0A4F8A4",
   273 => x"C0C0C0C0C0A4F8B0",
   274 => x"C0C0C0C0C0A4F899",
   275 => x"C0C0C0C0C0A4F892",
   276 => x"C0C0C0C0C0A4F882",
   277 => x"C0C0C0C0C0A4F8F8",
   278 => x"C0C0C0C0C0A4F880",
   279 => x"C0C0C0C0C0A4F890",
   280 => x"C0C0C0C0C0A480C0",
   281 => x"C0C0C0C0C0A480F9",
   282 => x"C0C0C0C0C0A480A4",
   283 => x"C0C0C0C0C0A480B0",
   284 => x"C0C0C0C0C0A48099",
   285 => x"C0C0C0C0C0A48092",
   286 => x"C0C0C0C0C0A48082",
   287 => x"C0C0C0C0C0A480F8",
   288 => x"C0C0C0C0C0A48080",
   289 => x"C0C0C0C0C0A48090",
   290 => x"C0C0C0C0C0A490C0",
   291 => x"C0C0C0C0C0A490F9",
   292 => x"C0C0C0C0C0A490A4",
   293 => x"C0C0C0C0C0A490B0",
   294 => x"C0C0C0C0C0A49099",
   295 => x"C0C0C0C0C0A49092",
   296 => x"C0C0C0C0C0A49082",
   297 => x"C0C0C0C0C0A490F8",
   298 => x"C0C0C0C0C0A49080",
   299 => x"C0C0C0C0C0A49090",
   300 => x"C0C0C0C0C0B0C0C0",
   301 => x"C0C0C0C0C0B0C0F9",
   302 => x"C0C0C0C0C0B0C0A4",
   303 => x"C0C0C0C0C0B0C0B0",
   304 => x"C0C0C0C0C0B0C099",
   305 => x"C0C0C0C0C0B0C092",
   306 => x"C0C0C0C0C0B0C082",
   307 => x"C0C0C0C0C0B0C0F8",
   308 => x"C0C0C0C0C0B0C080",
   309 => x"C0C0C0C0C0B0C090",
   310 => x"C0C0C0C0C0B0F9C0",
   311 => x"C0C0C0C0C0B0F9F9",
   312 => x"C0C0C0C0C0B0F9A4",
   313 => x"C0C0C0C0C0B0F9B0",
   314 => x"C0C0C0C0C0B0F999",
   315 => x"C0C0C0C0C0B0F992",
   316 => x"C0C0C0C0C0B0F982",
   317 => x"C0C0C0C0C0B0F9F8",
   318 => x"C0C0C0C0C0B0F980",
   319 => x"C0C0C0C0C0B0F990",
   320 => x"C0C0C0C0C0B0A4C0",
   321 => x"C0C0C0C0C0B0A4F9",
   322 => x"C0C0C0C0C0B0A4A4",
   323 => x"C0C0C0C0C0B0A4B0",
   324 => x"C0C0C0C0C0B0A499",
   325 => x"C0C0C0C0C0B0A492",
   326 => x"C0C0C0C0C0B0A482",
   327 => x"C0C0C0C0C0B0A4F8",
   328 => x"C0C0C0C0C0B0A480",
   329 => x"C0C0C0C0C0B0A490",
   330 => x"C0C0C0C0C0B0B0C0",
   331 => x"C0C0C0C0C0B0B0F9",
   332 => x"C0C0C0C0C0B0B0A4",
   333 => x"C0C0C0C0C0B0B0B0",
   334 => x"C0C0C0C0C0B0B099",
   335 => x"C0C0C0C0C0B0B092",
   336 => x"C0C0C0C0C0B0B082",
   337 => x"C0C0C0C0C0B0B0F8",
   338 => x"C0C0C0C0C0B0B080",
   339 => x"C0C0C0C0C0B0B090",
   340 => x"C0C0C0C0C0B099C0",
   341 => x"C0C0C0C0C0B099F9",
   342 => x"C0C0C0C0C0B099A4",
   343 => x"C0C0C0C0C0B099B0",
   344 => x"C0C0C0C0C0B09999",
   345 => x"C0C0C0C0C0B09992",
   346 => x"C0C0C0C0C0B09982",
   347 => x"C0C0C0C0C0B099F8",
   348 => x"C0C0C0C0C0B09980",
   349 => x"C0C0C0C0C0B09990",
   350 => x"C0C0C0C0C0B092C0",
   351 => x"C0C0C0C0C0B092F9",
   352 => x"C0C0C0C0C0B092A4",
   353 => x"C0C0C0C0C0B092B0",
   354 => x"C0C0C0C0C0B09299",
   355 => x"C0C0C0C0C0B09292",
   356 => x"C0C0C0C0C0B09282",
   357 => x"C0C0C0C0C0B092F8",
   358 => x"C0C0C0C0C0B09280",
   359 => x"C0C0C0C0C0B09290",
   360 => x"C0C0C0C0C0B082C0",
   361 => x"C0C0C0C0C0B082F9",
   362 => x"C0C0C0C0C0B082A4",
   363 => x"C0C0C0C0C0B082B0",
   364 => x"C0C0C0C0C0B08299",
   365 => x"C0C0C0C0C0B08292",
   366 => x"C0C0C0C0C0B08282",
   367 => x"C0C0C0C0C0B082F8",
   368 => x"C0C0C0C0C0B08280",
   369 => x"C0C0C0C0C0B08290",
   370 => x"C0C0C0C0C0B0F8C0",
   371 => x"C0C0C0C0C0B0F8F9",
   372 => x"C0C0C0C0C0B0F8A4",
   373 => x"C0C0C0C0C0B0F8B0",
   374 => x"C0C0C0C0C0B0F899",
   375 => x"C0C0C0C0C0B0F892",
   376 => x"C0C0C0C0C0B0F882",
   377 => x"C0C0C0C0C0B0F8F8",
   378 => x"C0C0C0C0C0B0F880",
   379 => x"C0C0C0C0C0B0F890",
   380 => x"C0C0C0C0C0B080C0",
   381 => x"C0C0C0C0C0B080F9",
   382 => x"C0C0C0C0C0B080A4",
   383 => x"C0C0C0C0C0B080B0",
   384 => x"C0C0C0C0C0B08099",
   385 => x"C0C0C0C0C0B08092",
   386 => x"C0C0C0C0C0B08082",
   387 => x"C0C0C0C0C0B080F8",
   388 => x"C0C0C0C0C0B08080",
   389 => x"C0C0C0C0C0B08090",
   390 => x"C0C0C0C0C0B090C0",
   391 => x"C0C0C0C0C0B090F9",
   392 => x"C0C0C0C0C0B090A4",
   393 => x"C0C0C0C0C0B090B0",
   394 => x"C0C0C0C0C0B09099",
   395 => x"C0C0C0C0C0B09092",
   396 => x"C0C0C0C0C0B09082",
   397 => x"C0C0C0C0C0B090F8",
   398 => x"C0C0C0C0C0B09080",
   399 => x"C0C0C0C0C0B09090",
   400 => x"C0C0C0C0C099C0C0",
   401 => x"C0C0C0C0C099C0F9",
   402 => x"C0C0C0C0C099C0A4",
   403 => x"C0C0C0C0C099C0B0",
   404 => x"C0C0C0C0C099C099",
   405 => x"C0C0C0C0C099C092",
   406 => x"C0C0C0C0C099C082",
   407 => x"C0C0C0C0C099C0F8",
   408 => x"C0C0C0C0C099C080",
   409 => x"C0C0C0C0C099C090",
   410 => x"C0C0C0C0C099F9C0",
   411 => x"C0C0C0C0C099F9F9",
   412 => x"C0C0C0C0C099F9A4",
   413 => x"C0C0C0C0C099F9B0",
   414 => x"C0C0C0C0C099F999",
   415 => x"C0C0C0C0C099F992",
   416 => x"C0C0C0C0C099F982",
   417 => x"C0C0C0C0C099F9F8",
   418 => x"C0C0C0C0C099F980",
   419 => x"C0C0C0C0C099F990",
   420 => x"C0C0C0C0C099A4C0",
   421 => x"C0C0C0C0C099A4F9",
   422 => x"C0C0C0C0C099A4A4",
   423 => x"C0C0C0C0C099A4B0",
   424 => x"C0C0C0C0C099A499",
   425 => x"C0C0C0C0C099A492",
   426 => x"C0C0C0C0C099A482",
   427 => x"C0C0C0C0C099A4F8",
   428 => x"C0C0C0C0C099A480",
   429 => x"C0C0C0C0C099A490",
   430 => x"C0C0C0C0C099B0C0",
   431 => x"C0C0C0C0C099B0F9",
   432 => x"C0C0C0C0C099B0A4",
   433 => x"C0C0C0C0C099B0B0",
   434 => x"C0C0C0C0C099B099",
   435 => x"C0C0C0C0C099B092",
   436 => x"C0C0C0C0C099B082",
   437 => x"C0C0C0C0C099B0F8",
   438 => x"C0C0C0C0C099B080",
   439 => x"C0C0C0C0C099B090",
   440 => x"C0C0C0C0C09999C0",
   441 => x"C0C0C0C0C09999F9",
   442 => x"C0C0C0C0C09999A4",
   443 => x"C0C0C0C0C09999B0",
   444 => x"C0C0C0C0C0999999",
   445 => x"C0C0C0C0C0999992",
   446 => x"C0C0C0C0C0999982",
   447 => x"C0C0C0C0C09999F8",
   448 => x"C0C0C0C0C0999980",
   449 => x"C0C0C0C0C0999990",
   450 => x"C0C0C0C0C09992C0",
   451 => x"C0C0C0C0C09992F9",
   452 => x"C0C0C0C0C09992A4",
   453 => x"C0C0C0C0C09992B0",
   454 => x"C0C0C0C0C0999299",
   455 => x"C0C0C0C0C0999292",
   456 => x"C0C0C0C0C0999282",
   457 => x"C0C0C0C0C09992F8",
   458 => x"C0C0C0C0C0999280",
   459 => x"C0C0C0C0C0999290",
   460 => x"C0C0C0C0C09982C0",
   461 => x"C0C0C0C0C09982F9",
   462 => x"C0C0C0C0C09982A4",
   463 => x"C0C0C0C0C09982B0",
   464 => x"C0C0C0C0C0998299",
   465 => x"C0C0C0C0C0998292",
   466 => x"C0C0C0C0C0998282",
   467 => x"C0C0C0C0C09982F8",
   468 => x"C0C0C0C0C0998280",
   469 => x"C0C0C0C0C0998290",
   470 => x"C0C0C0C0C099F8C0",
   471 => x"C0C0C0C0C099F8F9",
   472 => x"C0C0C0C0C099F8A4",
   473 => x"C0C0C0C0C099F8B0",
   474 => x"C0C0C0C0C099F899",
   475 => x"C0C0C0C0C099F892",
   476 => x"C0C0C0C0C099F882",
   477 => x"C0C0C0C0C099F8F8",
   478 => x"C0C0C0C0C099F880",
   479 => x"C0C0C0C0C099F890",
   480 => x"C0C0C0C0C09980C0",
   481 => x"C0C0C0C0C09980F9",
   482 => x"C0C0C0C0C09980A4",
   483 => x"C0C0C0C0C09980B0",
   484 => x"C0C0C0C0C0998099",
   485 => x"C0C0C0C0C0998092",
   486 => x"C0C0C0C0C0998082",
   487 => x"C0C0C0C0C09980F8",
   488 => x"C0C0C0C0C0998080",
   489 => x"C0C0C0C0C0998090",
   490 => x"C0C0C0C0C09990C0",
   491 => x"C0C0C0C0C09990F9",
   492 => x"C0C0C0C0C09990A4",
   493 => x"C0C0C0C0C09990B0",
   494 => x"C0C0C0C0C0999099",
   495 => x"C0C0C0C0C0999092",
   496 => x"C0C0C0C0C0999082",
   497 => x"C0C0C0C0C09990F8",
   498 => x"C0C0C0C0C0999080",
   499 => x"C0C0C0C0C0999090",
   500 => x"C0C0C0C0C092C0C0",
   501 => x"C0C0C0C0C092C0F9",
   502 => x"C0C0C0C0C092C0A4",
   503 => x"C0C0C0C0C092C0B0",
   504 => x"C0C0C0C0C092C099",
   505 => x"C0C0C0C0C092C092",
   506 => x"C0C0C0C0C092C082",
   507 => x"C0C0C0C0C092C0F8",
   508 => x"C0C0C0C0C092C080",
   509 => x"C0C0C0C0C092C090",
   510 => x"C0C0C0C0C092F9C0",
   511 => x"C0C0C0C0C092F9F9",
   512 => x"C0C0C0C0C092F9A4",
   513 => x"C0C0C0C0C092F9B0",
   514 => x"C0C0C0C0C092F999",
   515 => x"C0C0C0C0C092F992",
   516 => x"C0C0C0C0C092F982",
   517 => x"C0C0C0C0C092F9F8",
   518 => x"C0C0C0C0C092F980",
   519 => x"C0C0C0C0C092F990",
   520 => x"C0C0C0C0C092A4C0",
   521 => x"C0C0C0C0C092A4F9",
   522 => x"C0C0C0C0C092A4A4",
   523 => x"C0C0C0C0C092A4B0",
   524 => x"C0C0C0C0C092A499",
   525 => x"C0C0C0C0C092A492",
   526 => x"C0C0C0C0C092A482",
   527 => x"C0C0C0C0C092A4F8",
   528 => x"C0C0C0C0C092A480",
   529 => x"C0C0C0C0C092A490",
   530 => x"C0C0C0C0C092B0C0",
   531 => x"C0C0C0C0C092B0F9",
   532 => x"C0C0C0C0C092B0A4",
   533 => x"C0C0C0C0C092B0B0",
   534 => x"C0C0C0C0C092B099",
   535 => x"C0C0C0C0C092B092",
   536 => x"C0C0C0C0C092B082",
   537 => x"C0C0C0C0C092B0F8",
   538 => x"C0C0C0C0C092B080",
   539 => x"C0C0C0C0C092B090",
   540 => x"C0C0C0C0C09299C0",
   541 => x"C0C0C0C0C09299F9",
   542 => x"C0C0C0C0C09299A4",
   543 => x"C0C0C0C0C09299B0",
   544 => x"C0C0C0C0C0929999",
   545 => x"C0C0C0C0C0929992",
   546 => x"C0C0C0C0C0929982",
   547 => x"C0C0C0C0C09299F8",
   548 => x"C0C0C0C0C0929980",
   549 => x"C0C0C0C0C0929990",
   550 => x"C0C0C0C0C09292C0",
   551 => x"C0C0C0C0C09292F9",
   552 => x"C0C0C0C0C09292A4",
   553 => x"C0C0C0C0C09292B0",
   554 => x"C0C0C0C0C0929299",
   555 => x"C0C0C0C0C0929292",
   556 => x"C0C0C0C0C0929282",
   557 => x"C0C0C0C0C09292F8",
   558 => x"C0C0C0C0C0929280",
   559 => x"C0C0C0C0C0929290",
   560 => x"C0C0C0C0C09282C0",
   561 => x"C0C0C0C0C09282F9",
   562 => x"C0C0C0C0C09282A4",
   563 => x"C0C0C0C0C09282B0",
   564 => x"C0C0C0C0C0928299",
   565 => x"C0C0C0C0C0928292",
   566 => x"C0C0C0C0C0928282",
   567 => x"C0C0C0C0C09282F8",
   568 => x"C0C0C0C0C0928280",
   569 => x"C0C0C0C0C0928290",
   570 => x"C0C0C0C0C092F8C0",
   571 => x"C0C0C0C0C092F8F9",
   572 => x"C0C0C0C0C092F8A4",
   573 => x"C0C0C0C0C092F8B0",
   574 => x"C0C0C0C0C092F899",
   575 => x"C0C0C0C0C092F892",
   576 => x"C0C0C0C0C092F882",
   577 => x"C0C0C0C0C092F8F8",
   578 => x"C0C0C0C0C092F880",
   579 => x"C0C0C0C0C092F890",
   580 => x"C0C0C0C0C09280C0",
   581 => x"C0C0C0C0C09280F9",
   582 => x"C0C0C0C0C09280A4",
   583 => x"C0C0C0C0C09280B0",
   584 => x"C0C0C0C0C0928099",
   585 => x"C0C0C0C0C0928092",
   586 => x"C0C0C0C0C0928082",
   587 => x"C0C0C0C0C09280F8",
   588 => x"C0C0C0C0C0928080",
   589 => x"C0C0C0C0C0928090",
   590 => x"C0C0C0C0C09290C0",
   591 => x"C0C0C0C0C09290F9",
   592 => x"C0C0C0C0C09290A4",
   593 => x"C0C0C0C0C09290B0",
   594 => x"C0C0C0C0C0929099",
   595 => x"C0C0C0C0C0929092",
   596 => x"C0C0C0C0C0929082",
   597 => x"C0C0C0C0C09290F8",
   598 => x"C0C0C0C0C0929080",
   599 => x"C0C0C0C0C0929090",
   600 => x"C0C0C0C0C082C0C0",
   601 => x"C0C0C0C0C082C0F9",
   602 => x"C0C0C0C0C082C0A4",
   603 => x"C0C0C0C0C082C0B0",
   604 => x"C0C0C0C0C082C099",
   605 => x"C0C0C0C0C082C092",
   606 => x"C0C0C0C0C082C082",
   607 => x"C0C0C0C0C082C0F8",
   608 => x"C0C0C0C0C082C080",
   609 => x"C0C0C0C0C082C090",
   610 => x"C0C0C0C0C082F9C0",
   611 => x"C0C0C0C0C082F9F9",
   612 => x"C0C0C0C0C082F9A4",
   613 => x"C0C0C0C0C082F9B0",
   614 => x"C0C0C0C0C082F999",
   615 => x"C0C0C0C0C082F992",
   616 => x"C0C0C0C0C082F982",
   617 => x"C0C0C0C0C082F9F8",
   618 => x"C0C0C0C0C082F980",
   619 => x"C0C0C0C0C082F990",
   620 => x"C0C0C0C0C082A4C0",
   621 => x"C0C0C0C0C082A4F9",
   622 => x"C0C0C0C0C082A4A4",
   623 => x"C0C0C0C0C082A4B0",
   624 => x"C0C0C0C0C082A499",
   625 => x"C0C0C0C0C082A492",
   626 => x"C0C0C0C0C082A482",
   627 => x"C0C0C0C0C082A4F8",
   628 => x"C0C0C0C0C082A480",
   629 => x"C0C0C0C0C082A490",
   630 => x"C0C0C0C0C082B0C0",
   631 => x"C0C0C0C0C082B0F9",
   632 => x"C0C0C0C0C082B0A4",
   633 => x"C0C0C0C0C082B0B0",
   634 => x"C0C0C0C0C082B099",
   635 => x"C0C0C0C0C082B092",
   636 => x"C0C0C0C0C082B082",
   637 => x"C0C0C0C0C082B0F8",
   638 => x"C0C0C0C0C082B080",
   639 => x"C0C0C0C0C082B090",
   640 => x"C0C0C0C0C08299C0",
   641 => x"C0C0C0C0C08299F9",
   642 => x"C0C0C0C0C08299A4",
   643 => x"C0C0C0C0C08299B0",
   644 => x"C0C0C0C0C0829999",
   645 => x"C0C0C0C0C0829992",
   646 => x"C0C0C0C0C0829982",
   647 => x"C0C0C0C0C08299F8",
   648 => x"C0C0C0C0C0829980",
   649 => x"C0C0C0C0C0829990",
   650 => x"C0C0C0C0C08292C0",
   651 => x"C0C0C0C0C08292F9",
   652 => x"C0C0C0C0C08292A4",
   653 => x"C0C0C0C0C08292B0",
   654 => x"C0C0C0C0C0829299",
   655 => x"C0C0C0C0C0829292",
   656 => x"C0C0C0C0C0829282",
   657 => x"C0C0C0C0C08292F8",
   658 => x"C0C0C0C0C0829280",
   659 => x"C0C0C0C0C0829290",
   660 => x"C0C0C0C0C08282C0",
   661 => x"C0C0C0C0C08282F9",
   662 => x"C0C0C0C0C08282A4",
   663 => x"C0C0C0C0C08282B0",
   664 => x"C0C0C0C0C0828299",
   665 => x"C0C0C0C0C0828292",
   666 => x"C0C0C0C0C0828282",
   667 => x"C0C0C0C0C08282F8",
   668 => x"C0C0C0C0C0828280",
   669 => x"C0C0C0C0C0828290",
   670 => x"C0C0C0C0C082F8C0",
   671 => x"C0C0C0C0C082F8F9",
   672 => x"C0C0C0C0C082F8A4",
   673 => x"C0C0C0C0C082F8B0",
   674 => x"C0C0C0C0C082F899",
   675 => x"C0C0C0C0C082F892",
   676 => x"C0C0C0C0C082F882",
   677 => x"C0C0C0C0C082F8F8",
   678 => x"C0C0C0C0C082F880",
   679 => x"C0C0C0C0C082F890",
   680 => x"C0C0C0C0C08280C0",
   681 => x"C0C0C0C0C08280F9",
   682 => x"C0C0C0C0C08280A4",
   683 => x"C0C0C0C0C08280B0",
   684 => x"C0C0C0C0C0828099",
   685 => x"C0C0C0C0C0828092",
   686 => x"C0C0C0C0C0828082",
   687 => x"C0C0C0C0C08280F8",
   688 => x"C0C0C0C0C0828080",
   689 => x"C0C0C0C0C0828090",
   690 => x"C0C0C0C0C08290C0",
   691 => x"C0C0C0C0C08290F9",
   692 => x"C0C0C0C0C08290A4",
   693 => x"C0C0C0C0C08290B0",
   694 => x"C0C0C0C0C0829099",
   695 => x"C0C0C0C0C0829092",
   696 => x"C0C0C0C0C0829082",
   697 => x"C0C0C0C0C08290F8",
   698 => x"C0C0C0C0C0829080",
   699 => x"C0C0C0C0C0829090",
   700 => x"C0C0C0C0C0F8C0C0",
   701 => x"C0C0C0C0C0F8C0F9",
   702 => x"C0C0C0C0C0F8C0A4",
   703 => x"C0C0C0C0C0F8C0B0",
   704 => x"C0C0C0C0C0F8C099",
   705 => x"C0C0C0C0C0F8C092",
   706 => x"C0C0C0C0C0F8C082",
   707 => x"C0C0C0C0C0F8C0F8",
   708 => x"C0C0C0C0C0F8C080",
   709 => x"C0C0C0C0C0F8C090",
   710 => x"C0C0C0C0C0F8F9C0",
   711 => x"C0C0C0C0C0F8F9F9",
   712 => x"C0C0C0C0C0F8F9A4",
   713 => x"C0C0C0C0C0F8F9B0",
   714 => x"C0C0C0C0C0F8F999",
   715 => x"C0C0C0C0C0F8F992",
   716 => x"C0C0C0C0C0F8F982",
   717 => x"C0C0C0C0C0F8F9F8",
   718 => x"C0C0C0C0C0F8F980",
   719 => x"C0C0C0C0C0F8F990",
   720 => x"C0C0C0C0C0F8A4C0",
   721 => x"C0C0C0C0C0F8A4F9",
   722 => x"C0C0C0C0C0F8A4A4",
   723 => x"C0C0C0C0C0F8A4B0",
   724 => x"C0C0C0C0C0F8A499",
   725 => x"C0C0C0C0C0F8A492",
   726 => x"C0C0C0C0C0F8A482",
   727 => x"C0C0C0C0C0F8A4F8",
   728 => x"C0C0C0C0C0F8A480",
   729 => x"C0C0C0C0C0F8A490",
   730 => x"C0C0C0C0C0F8B0C0",
   731 => x"C0C0C0C0C0F8B0F9",
   732 => x"C0C0C0C0C0F8B0A4",
   733 => x"C0C0C0C0C0F8B0B0",
   734 => x"C0C0C0C0C0F8B099",
   735 => x"C0C0C0C0C0F8B092",
   736 => x"C0C0C0C0C0F8B082",
   737 => x"C0C0C0C0C0F8B0F8",
   738 => x"C0C0C0C0C0F8B080",
   739 => x"C0C0C0C0C0F8B090",
   740 => x"C0C0C0C0C0F899C0",
   741 => x"C0C0C0C0C0F899F9",
   742 => x"C0C0C0C0C0F899A4",
   743 => x"C0C0C0C0C0F899B0",
   744 => x"C0C0C0C0C0F89999",
   745 => x"C0C0C0C0C0F89992",
   746 => x"C0C0C0C0C0F89982",
   747 => x"C0C0C0C0C0F899F8",
   748 => x"C0C0C0C0C0F89980",
   749 => x"C0C0C0C0C0F89990",
   750 => x"C0C0C0C0C0F892C0",
   751 => x"C0C0C0C0C0F892F9",
   752 => x"C0C0C0C0C0F892A4",
   753 => x"C0C0C0C0C0F892B0",
   754 => x"C0C0C0C0C0F89299",
   755 => x"C0C0C0C0C0F89292",
   756 => x"C0C0C0C0C0F89282",
   757 => x"C0C0C0C0C0F892F8",
   758 => x"C0C0C0C0C0F89280",
   759 => x"C0C0C0C0C0F89290",
   760 => x"C0C0C0C0C0F882C0",
   761 => x"C0C0C0C0C0F882F9",
   762 => x"C0C0C0C0C0F882A4",
   763 => x"C0C0C0C0C0F882B0",
   764 => x"C0C0C0C0C0F88299",
   765 => x"C0C0C0C0C0F88292",
   766 => x"C0C0C0C0C0F88282",
   767 => x"C0C0C0C0C0F882F8",
   768 => x"C0C0C0C0C0F88280",
   769 => x"C0C0C0C0C0F88290",
   770 => x"C0C0C0C0C0F8F8C0",
   771 => x"C0C0C0C0C0F8F8F9",
   772 => x"C0C0C0C0C0F8F8A4",
   773 => x"C0C0C0C0C0F8F8B0",
   774 => x"C0C0C0C0C0F8F899",
   775 => x"C0C0C0C0C0F8F892",
   776 => x"C0C0C0C0C0F8F882",
   777 => x"C0C0C0C0C0F8F8F8",
   778 => x"C0C0C0C0C0F8F880",
   779 => x"C0C0C0C0C0F8F890",
   780 => x"C0C0C0C0C0F880C0",
   781 => x"C0C0C0C0C0F880F9",
   782 => x"C0C0C0C0C0F880A4",
   783 => x"C0C0C0C0C0F880B0",
   784 => x"C0C0C0C0C0F88099",
   785 => x"C0C0C0C0C0F88092",
   786 => x"C0C0C0C0C0F88082",
   787 => x"C0C0C0C0C0F880F8",
   788 => x"C0C0C0C0C0F88080",
   789 => x"C0C0C0C0C0F88090",
   790 => x"C0C0C0C0C0F890C0",
   791 => x"C0C0C0C0C0F890F9",
   792 => x"C0C0C0C0C0F890A4",
   793 => x"C0C0C0C0C0F890B0",
   794 => x"C0C0C0C0C0F89099",
   795 => x"C0C0C0C0C0F89092",
   796 => x"C0C0C0C0C0F89082",
   797 => x"C0C0C0C0C0F890F8",
   798 => x"C0C0C0C0C0F89080",
   799 => x"C0C0C0C0C0F89090",
   800 => x"C0C0C0C0C080C0C0",
   801 => x"C0C0C0C0C080C0F9",
   802 => x"C0C0C0C0C080C0A4",
   803 => x"C0C0C0C0C080C0B0",
   804 => x"C0C0C0C0C080C099",
   805 => x"C0C0C0C0C080C092",
   806 => x"C0C0C0C0C080C082",
   807 => x"C0C0C0C0C080C0F8",
   808 => x"C0C0C0C0C080C080",
   809 => x"C0C0C0C0C080C090",
   810 => x"C0C0C0C0C080F9C0",
   811 => x"C0C0C0C0C080F9F9",
   812 => x"C0C0C0C0C080F9A4",
   813 => x"C0C0C0C0C080F9B0",
   814 => x"C0C0C0C0C080F999",
   815 => x"C0C0C0C0C080F992",
   816 => x"C0C0C0C0C080F982",
   817 => x"C0C0C0C0C080F9F8",
   818 => x"C0C0C0C0C080F980",
   819 => x"C0C0C0C0C080F990",
   820 => x"C0C0C0C0C080A4C0",
   821 => x"C0C0C0C0C080A4F9",
   822 => x"C0C0C0C0C080A4A4",
   823 => x"C0C0C0C0C080A4B0",
   824 => x"C0C0C0C0C080A499",
   825 => x"C0C0C0C0C080A492",
   826 => x"C0C0C0C0C080A482",
   827 => x"C0C0C0C0C080A4F8",
   828 => x"C0C0C0C0C080A480",
   829 => x"C0C0C0C0C080A490",
   830 => x"C0C0C0C0C080B0C0",
   831 => x"C0C0C0C0C080B0F9",
   832 => x"C0C0C0C0C080B0A4",
   833 => x"C0C0C0C0C080B0B0",
   834 => x"C0C0C0C0C080B099",
   835 => x"C0C0C0C0C080B092",
   836 => x"C0C0C0C0C080B082",
   837 => x"C0C0C0C0C080B0F8",
   838 => x"C0C0C0C0C080B080",
   839 => x"C0C0C0C0C080B090",
   840 => x"C0C0C0C0C08099C0",
   841 => x"C0C0C0C0C08099F9",
   842 => x"C0C0C0C0C08099A4",
   843 => x"C0C0C0C0C08099B0",
   844 => x"C0C0C0C0C0809999",
   845 => x"C0C0C0C0C0809992",
   846 => x"C0C0C0C0C0809982",
   847 => x"C0C0C0C0C08099F8",
   848 => x"C0C0C0C0C0809980",
   849 => x"C0C0C0C0C0809990",
   850 => x"C0C0C0C0C08092C0",
   851 => x"C0C0C0C0C08092F9",
   852 => x"C0C0C0C0C08092A4",
   853 => x"C0C0C0C0C08092B0",
   854 => x"C0C0C0C0C0809299",
   855 => x"C0C0C0C0C0809292",
   856 => x"C0C0C0C0C0809282",
   857 => x"C0C0C0C0C08092F8",
   858 => x"C0C0C0C0C0809280",
   859 => x"C0C0C0C0C0809290",
   860 => x"C0C0C0C0C08082C0",
   861 => x"C0C0C0C0C08082F9",
   862 => x"C0C0C0C0C08082A4",
   863 => x"C0C0C0C0C08082B0",
   864 => x"C0C0C0C0C0808299",
   865 => x"C0C0C0C0C0808292",
   866 => x"C0C0C0C0C0808282",
   867 => x"C0C0C0C0C08082F8",
   868 => x"C0C0C0C0C0808280",
   869 => x"C0C0C0C0C0808290",
   870 => x"C0C0C0C0C080F8C0",
   871 => x"C0C0C0C0C080F8F9",
   872 => x"C0C0C0C0C080F8A4",
   873 => x"C0C0C0C0C080F8B0",
   874 => x"C0C0C0C0C080F899",
   875 => x"C0C0C0C0C080F892",
   876 => x"C0C0C0C0C080F882",
   877 => x"C0C0C0C0C080F8F8",
   878 => x"C0C0C0C0C080F880",
   879 => x"C0C0C0C0C080F890",
   880 => x"C0C0C0C0C08080C0",
   881 => x"C0C0C0C0C08080F9",
   882 => x"C0C0C0C0C08080A4",
   883 => x"C0C0C0C0C08080B0",
   884 => x"C0C0C0C0C0808099",
   885 => x"C0C0C0C0C0808092",
   886 => x"C0C0C0C0C0808082",
   887 => x"C0C0C0C0C08080F8",
   888 => x"C0C0C0C0C0808080",
   889 => x"C0C0C0C0C0808090",
   890 => x"C0C0C0C0C08090C0",
   891 => x"C0C0C0C0C08090F9",
   892 => x"C0C0C0C0C08090A4",
   893 => x"C0C0C0C0C08090B0",
   894 => x"C0C0C0C0C0809099",
   895 => x"C0C0C0C0C0809092",
   896 => x"C0C0C0C0C0809082",
   897 => x"C0C0C0C0C08090F8",
   898 => x"C0C0C0C0C0809080",
   899 => x"C0C0C0C0C0809090",
   900 => x"C0C0C0C0C090C0C0",
   901 => x"C0C0C0C0C090C0F9",
   902 => x"C0C0C0C0C090C0A4",
   903 => x"C0C0C0C0C090C0B0",
   904 => x"C0C0C0C0C090C099",
   905 => x"C0C0C0C0C090C092",
   906 => x"C0C0C0C0C090C082",
   907 => x"C0C0C0C0C090C0F8",
   908 => x"C0C0C0C0C090C080",
   909 => x"C0C0C0C0C090C090",
   910 => x"C0C0C0C0C090F9C0",
   911 => x"C0C0C0C0C090F9F9",
   912 => x"C0C0C0C0C090F9A4",
   913 => x"C0C0C0C0C090F9B0",
   914 => x"C0C0C0C0C090F999",
   915 => x"C0C0C0C0C090F992",
   916 => x"C0C0C0C0C090F982",
   917 => x"C0C0C0C0C090F9F8",
   918 => x"C0C0C0C0C090F980",
   919 => x"C0C0C0C0C090F990",
   920 => x"C0C0C0C0C090A4C0",
   921 => x"C0C0C0C0C090A4F9",
   922 => x"C0C0C0C0C090A4A4",
   923 => x"C0C0C0C0C090A4B0",
   924 => x"C0C0C0C0C090A499",
   925 => x"C0C0C0C0C090A492",
   926 => x"C0C0C0C0C090A482",
   927 => x"C0C0C0C0C090A4F8",
   928 => x"C0C0C0C0C090A480",
   929 => x"C0C0C0C0C090A490",
   930 => x"C0C0C0C0C090B0C0",
   931 => x"C0C0C0C0C090B0F9",
   932 => x"C0C0C0C0C090B0A4",
   933 => x"C0C0C0C0C090B0B0",
   934 => x"C0C0C0C0C090B099",
   935 => x"C0C0C0C0C090B092",
   936 => x"C0C0C0C0C090B082",
   937 => x"C0C0C0C0C090B0F8",
   938 => x"C0C0C0C0C090B080",
   939 => x"C0C0C0C0C090B090",
   940 => x"C0C0C0C0C09099C0",
   941 => x"C0C0C0C0C09099F9",
   942 => x"C0C0C0C0C09099A4",
   943 => x"C0C0C0C0C09099B0",
   944 => x"C0C0C0C0C0909999",
   945 => x"C0C0C0C0C0909992",
   946 => x"C0C0C0C0C0909982",
   947 => x"C0C0C0C0C09099F8",
   948 => x"C0C0C0C0C0909980",
   949 => x"C0C0C0C0C0909990",
   950 => x"C0C0C0C0C09092C0",
   951 => x"C0C0C0C0C09092F9",
   952 => x"C0C0C0C0C09092A4",
   953 => x"C0C0C0C0C09092B0",
   954 => x"C0C0C0C0C0909299",
   955 => x"C0C0C0C0C0909292",
   956 => x"C0C0C0C0C0909282",
   957 => x"C0C0C0C0C09092F8",
   958 => x"C0C0C0C0C0909280",
   959 => x"C0C0C0C0C0909290",
   960 => x"C0C0C0C0C09082C0",
   961 => x"C0C0C0C0C09082F9",
   962 => x"C0C0C0C0C09082A4",
   963 => x"C0C0C0C0C09082B0",
   964 => x"C0C0C0C0C0908299",
   965 => x"C0C0C0C0C0908292",
   966 => x"C0C0C0C0C0908282",
   967 => x"C0C0C0C0C09082F8",
   968 => x"C0C0C0C0C0908280",
   969 => x"C0C0C0C0C0908290",
   970 => x"C0C0C0C0C090F8C0",
   971 => x"C0C0C0C0C090F8F9",
   972 => x"C0C0C0C0C090F8A4",
   973 => x"C0C0C0C0C090F8B0",
   974 => x"C0C0C0C0C090F899",
   975 => x"C0C0C0C0C090F892",
   976 => x"C0C0C0C0C090F882",
   977 => x"C0C0C0C0C090F8F8",
   978 => x"C0C0C0C0C090F880",
   979 => x"C0C0C0C0C090F890",
   980 => x"C0C0C0C0C09080C0",
   981 => x"C0C0C0C0C09080F9",
   982 => x"C0C0C0C0C09080A4",
   983 => x"C0C0C0C0C09080B0",
   984 => x"C0C0C0C0C0908099",
   985 => x"C0C0C0C0C0908092",
   986 => x"C0C0C0C0C0908082",
   987 => x"C0C0C0C0C09080F8",
   988 => x"C0C0C0C0C0908080",
   989 => x"C0C0C0C0C0908090",
   990 => x"C0C0C0C0C09090C0",
   991 => x"C0C0C0C0C09090F9",
   992 => x"C0C0C0C0C09090A4",
   993 => x"C0C0C0C0C09090B0",
   994 => x"C0C0C0C0C0909099",
   995 => x"C0C0C0C0C0909092",
   996 => x"C0C0C0C0C0909082",
   997 => x"C0C0C0C0C09090F8",
   998 => x"C0C0C0C0C0909080",
   999 => x"C0C0C0C0C0909090",
  1000 => x"C0C0C0C0F9C0C0C0",
  1001 => x"C0C0C0C0F9C0C0F9",
  1002 => x"C0C0C0C0F9C0C0A4",
  1003 => x"C0C0C0C0F9C0C0B0",
  1004 => x"C0C0C0C0F9C0C099",
  1005 => x"C0C0C0C0F9C0C092",
  1006 => x"C0C0C0C0F9C0C082",
  1007 => x"C0C0C0C0F9C0C0F8",
  1008 => x"C0C0C0C0F9C0C080",
  1009 => x"C0C0C0C0F9C0C090",
  1010 => x"C0C0C0C0F9C0F9C0",
  1011 => x"C0C0C0C0F9C0F9F9",
  1012 => x"C0C0C0C0F9C0F9A4",
  1013 => x"C0C0C0C0F9C0F9B0",
  1014 => x"C0C0C0C0F9C0F999",
  1015 => x"C0C0C0C0F9C0F992",
  1016 => x"C0C0C0C0F9C0F982",
  1017 => x"C0C0C0C0F9C0F9F8",
  1018 => x"C0C0C0C0F9C0F980",
  1019 => x"C0C0C0C0F9C0F990",
  1020 => x"C0C0C0C0F9C0A4C0",
  1021 => x"C0C0C0C0F9C0A4F9",
  1022 => x"C0C0C0C0F9C0A4A4",
  1023 => x"C0C0C0C0F9C0A4B0",
  1024 => x"C0C0C0C0F9C0A499",
  1025 => x"C0C0C0C0F9C0A492",
  1026 => x"C0C0C0C0F9C0A482",
  1027 => x"C0C0C0C0F9C0A4F8",
  1028 => x"C0C0C0C0F9C0A480",
  1029 => x"C0C0C0C0F9C0A490",
  1030 => x"C0C0C0C0F9C0B0C0",
  1031 => x"C0C0C0C0F9C0B0F9",
  1032 => x"C0C0C0C0F9C0B0A4",
  1033 => x"C0C0C0C0F9C0B0B0",
  1034 => x"C0C0C0C0F9C0B099",
  1035 => x"C0C0C0C0F9C0B092",
  1036 => x"C0C0C0C0F9C0B082",
  1037 => x"C0C0C0C0F9C0B0F8",
  1038 => x"C0C0C0C0F9C0B080",
  1039 => x"C0C0C0C0F9C0B090",
  1040 => x"C0C0C0C0F9C099C0",
  1041 => x"C0C0C0C0F9C099F9",
  1042 => x"C0C0C0C0F9C099A4",
  1043 => x"C0C0C0C0F9C099B0",
  1044 => x"C0C0C0C0F9C09999",
  1045 => x"C0C0C0C0F9C09992",
  1046 => x"C0C0C0C0F9C09982",
  1047 => x"C0C0C0C0F9C099F8",
  1048 => x"C0C0C0C0F9C09980",
  1049 => x"C0C0C0C0F9C09990",
  1050 => x"C0C0C0C0F9C092C0",
  1051 => x"C0C0C0C0F9C092F9",
  1052 => x"C0C0C0C0F9C092A4",
  1053 => x"C0C0C0C0F9C092B0",
  1054 => x"C0C0C0C0F9C09299",
  1055 => x"C0C0C0C0F9C09292",
  1056 => x"C0C0C0C0F9C09282",
  1057 => x"C0C0C0C0F9C092F8",
  1058 => x"C0C0C0C0F9C09280",
  1059 => x"C0C0C0C0F9C09290",
  1060 => x"C0C0C0C0F9C082C0",
  1061 => x"C0C0C0C0F9C082F9",
  1062 => x"C0C0C0C0F9C082A4",
  1063 => x"C0C0C0C0F9C082B0",
  1064 => x"C0C0C0C0F9C08299",
  1065 => x"C0C0C0C0F9C08292",
  1066 => x"C0C0C0C0F9C08282",
  1067 => x"C0C0C0C0F9C082F8",
  1068 => x"C0C0C0C0F9C08280",
  1069 => x"C0C0C0C0F9C08290",
  1070 => x"C0C0C0C0F9C0F8C0",
  1071 => x"C0C0C0C0F9C0F8F9",
  1072 => x"C0C0C0C0F9C0F8A4",
  1073 => x"C0C0C0C0F9C0F8B0",
  1074 => x"C0C0C0C0F9C0F899",
  1075 => x"C0C0C0C0F9C0F892",
  1076 => x"C0C0C0C0F9C0F882",
  1077 => x"C0C0C0C0F9C0F8F8",
  1078 => x"C0C0C0C0F9C0F880",
  1079 => x"C0C0C0C0F9C0F890",
  1080 => x"C0C0C0C0F9C080C0",
  1081 => x"C0C0C0C0F9C080F9",
  1082 => x"C0C0C0C0F9C080A4",
  1083 => x"C0C0C0C0F9C080B0",
  1084 => x"C0C0C0C0F9C08099",
  1085 => x"C0C0C0C0F9C08092",
  1086 => x"C0C0C0C0F9C08082",
  1087 => x"C0C0C0C0F9C080F8",
  1088 => x"C0C0C0C0F9C08080",
  1089 => x"C0C0C0C0F9C08090",
  1090 => x"C0C0C0C0F9C090C0",
  1091 => x"C0C0C0C0F9C090F9",
  1092 => x"C0C0C0C0F9C090A4",
  1093 => x"C0C0C0C0F9C090B0",
  1094 => x"C0C0C0C0F9C09099",
  1095 => x"C0C0C0C0F9C09092",
  1096 => x"C0C0C0C0F9C09082",
  1097 => x"C0C0C0C0F9C090F8",
  1098 => x"C0C0C0C0F9C09080",
  1099 => x"C0C0C0C0F9C09090",
  1100 => x"C0C0C0C0F9F9C0C0",
  1101 => x"C0C0C0C0F9F9C0F9",
  1102 => x"C0C0C0C0F9F9C0A4",
  1103 => x"C0C0C0C0F9F9C0B0",
  1104 => x"C0C0C0C0F9F9C099",
  1105 => x"C0C0C0C0F9F9C092",
  1106 => x"C0C0C0C0F9F9C082",
  1107 => x"C0C0C0C0F9F9C0F8",
  1108 => x"C0C0C0C0F9F9C080",
  1109 => x"C0C0C0C0F9F9C090",
  1110 => x"C0C0C0C0F9F9F9C0",
  1111 => x"C0C0C0C0F9F9F9F9",
  1112 => x"C0C0C0C0F9F9F9A4",
  1113 => x"C0C0C0C0F9F9F9B0",
  1114 => x"C0C0C0C0F9F9F999",
  1115 => x"C0C0C0C0F9F9F992",
  1116 => x"C0C0C0C0F9F9F982",
  1117 => x"C0C0C0C0F9F9F9F8",
  1118 => x"C0C0C0C0F9F9F980",
  1119 => x"C0C0C0C0F9F9F990",
  1120 => x"C0C0C0C0F9F9A4C0",
  1121 => x"C0C0C0C0F9F9A4F9",
  1122 => x"C0C0C0C0F9F9A4A4",
  1123 => x"C0C0C0C0F9F9A4B0",
  1124 => x"C0C0C0C0F9F9A499",
  1125 => x"C0C0C0C0F9F9A492",
  1126 => x"C0C0C0C0F9F9A482",
  1127 => x"C0C0C0C0F9F9A4F8",
  1128 => x"C0C0C0C0F9F9A480",
  1129 => x"C0C0C0C0F9F9A490",
  1130 => x"C0C0C0C0F9F9B0C0",
  1131 => x"C0C0C0C0F9F9B0F9",
  1132 => x"C0C0C0C0F9F9B0A4",
  1133 => x"C0C0C0C0F9F9B0B0",
  1134 => x"C0C0C0C0F9F9B099",
  1135 => x"C0C0C0C0F9F9B092",
  1136 => x"C0C0C0C0F9F9B082",
  1137 => x"C0C0C0C0F9F9B0F8",
  1138 => x"C0C0C0C0F9F9B080",
  1139 => x"C0C0C0C0F9F9B090",
  1140 => x"C0C0C0C0F9F999C0",
  1141 => x"C0C0C0C0F9F999F9",
  1142 => x"C0C0C0C0F9F999A4",
  1143 => x"C0C0C0C0F9F999B0",
  1144 => x"C0C0C0C0F9F99999",
  1145 => x"C0C0C0C0F9F99992",
  1146 => x"C0C0C0C0F9F99982",
  1147 => x"C0C0C0C0F9F999F8",
  1148 => x"C0C0C0C0F9F99980",
  1149 => x"C0C0C0C0F9F99990",
  1150 => x"C0C0C0C0F9F992C0",
  1151 => x"C0C0C0C0F9F992F9",
  1152 => x"C0C0C0C0F9F992A4",
  1153 => x"C0C0C0C0F9F992B0",
  1154 => x"C0C0C0C0F9F99299",
  1155 => x"C0C0C0C0F9F99292",
  1156 => x"C0C0C0C0F9F99282",
  1157 => x"C0C0C0C0F9F992F8",
  1158 => x"C0C0C0C0F9F99280",
  1159 => x"C0C0C0C0F9F99290",
  1160 => x"C0C0C0C0F9F982C0",
  1161 => x"C0C0C0C0F9F982F9",
  1162 => x"C0C0C0C0F9F982A4",
  1163 => x"C0C0C0C0F9F982B0",
  1164 => x"C0C0C0C0F9F98299",
  1165 => x"C0C0C0C0F9F98292",
  1166 => x"C0C0C0C0F9F98282",
  1167 => x"C0C0C0C0F9F982F8",
  1168 => x"C0C0C0C0F9F98280",
  1169 => x"C0C0C0C0F9F98290",
  1170 => x"C0C0C0C0F9F9F8C0",
  1171 => x"C0C0C0C0F9F9F8F9",
  1172 => x"C0C0C0C0F9F9F8A4",
  1173 => x"C0C0C0C0F9F9F8B0",
  1174 => x"C0C0C0C0F9F9F899",
  1175 => x"C0C0C0C0F9F9F892",
  1176 => x"C0C0C0C0F9F9F882",
  1177 => x"C0C0C0C0F9F9F8F8",
  1178 => x"C0C0C0C0F9F9F880",
  1179 => x"C0C0C0C0F9F9F890",
  1180 => x"C0C0C0C0F9F980C0",
  1181 => x"C0C0C0C0F9F980F9",
  1182 => x"C0C0C0C0F9F980A4",
  1183 => x"C0C0C0C0F9F980B0",
  1184 => x"C0C0C0C0F9F98099",
  1185 => x"C0C0C0C0F9F98092",
  1186 => x"C0C0C0C0F9F98082",
  1187 => x"C0C0C0C0F9F980F8",
  1188 => x"C0C0C0C0F9F98080",
  1189 => x"C0C0C0C0F9F98090",
  1190 => x"C0C0C0C0F9F990C0",
  1191 => x"C0C0C0C0F9F990F9",
  1192 => x"C0C0C0C0F9F990A4",
  1193 => x"C0C0C0C0F9F990B0",
  1194 => x"C0C0C0C0F9F99099",
  1195 => x"C0C0C0C0F9F99092",
  1196 => x"C0C0C0C0F9F99082",
  1197 => x"C0C0C0C0F9F990F8",
  1198 => x"C0C0C0C0F9F99080",
  1199 => x"C0C0C0C0F9F99090",
  1200 => x"C0C0C0C0F9A4C0C0",
  1201 => x"C0C0C0C0F9A4C0F9",
  1202 => x"C0C0C0C0F9A4C0A4",
  1203 => x"C0C0C0C0F9A4C0B0",
  1204 => x"C0C0C0C0F9A4C099",
  1205 => x"C0C0C0C0F9A4C092",
  1206 => x"C0C0C0C0F9A4C082",
  1207 => x"C0C0C0C0F9A4C0F8",
  1208 => x"C0C0C0C0F9A4C080",
  1209 => x"C0C0C0C0F9A4C090",
  1210 => x"C0C0C0C0F9A4F9C0",
  1211 => x"C0C0C0C0F9A4F9F9",
  1212 => x"C0C0C0C0F9A4F9A4",
  1213 => x"C0C0C0C0F9A4F9B0",
  1214 => x"C0C0C0C0F9A4F999",
  1215 => x"C0C0C0C0F9A4F992",
  1216 => x"C0C0C0C0F9A4F982",
  1217 => x"C0C0C0C0F9A4F9F8",
  1218 => x"C0C0C0C0F9A4F980",
  1219 => x"C0C0C0C0F9A4F990",
  1220 => x"C0C0C0C0F9A4A4C0",
  1221 => x"C0C0C0C0F9A4A4F9",
  1222 => x"C0C0C0C0F9A4A4A4",
  1223 => x"C0C0C0C0F9A4A4B0",
  1224 => x"C0C0C0C0F9A4A499",
  1225 => x"C0C0C0C0F9A4A492",
  1226 => x"C0C0C0C0F9A4A482",
  1227 => x"C0C0C0C0F9A4A4F8",
  1228 => x"C0C0C0C0F9A4A480",
  1229 => x"C0C0C0C0F9A4A490",
  1230 => x"C0C0C0C0F9A4B0C0",
  1231 => x"C0C0C0C0F9A4B0F9",
  1232 => x"C0C0C0C0F9A4B0A4",
  1233 => x"C0C0C0C0F9A4B0B0",
  1234 => x"C0C0C0C0F9A4B099",
  1235 => x"C0C0C0C0F9A4B092",
  1236 => x"C0C0C0C0F9A4B082",
  1237 => x"C0C0C0C0F9A4B0F8",
  1238 => x"C0C0C0C0F9A4B080",
  1239 => x"C0C0C0C0F9A4B090",
  1240 => x"C0C0C0C0F9A499C0",
  1241 => x"C0C0C0C0F9A499F9",
  1242 => x"C0C0C0C0F9A499A4",
  1243 => x"C0C0C0C0F9A499B0",
  1244 => x"C0C0C0C0F9A49999",
  1245 => x"C0C0C0C0F9A49992",
  1246 => x"C0C0C0C0F9A49982",
  1247 => x"C0C0C0C0F9A499F8",
  1248 => x"C0C0C0C0F9A49980",
  1249 => x"C0C0C0C0F9A49990",
  1250 => x"C0C0C0C0F9A492C0",
  1251 => x"C0C0C0C0F9A492F9",
  1252 => x"C0C0C0C0F9A492A4",
  1253 => x"C0C0C0C0F9A492B0",
  1254 => x"C0C0C0C0F9A49299",
  1255 => x"C0C0C0C0F9A49292",
  1256 => x"C0C0C0C0F9A49282",
  1257 => x"C0C0C0C0F9A492F8",
  1258 => x"C0C0C0C0F9A49280",
  1259 => x"C0C0C0C0F9A49290",
  1260 => x"C0C0C0C0F9A482C0",
  1261 => x"C0C0C0C0F9A482F9",
  1262 => x"C0C0C0C0F9A482A4",
  1263 => x"C0C0C0C0F9A482B0",
  1264 => x"C0C0C0C0F9A48299",
  1265 => x"C0C0C0C0F9A48292",
  1266 => x"C0C0C0C0F9A48282",
  1267 => x"C0C0C0C0F9A482F8",
  1268 => x"C0C0C0C0F9A48280",
  1269 => x"C0C0C0C0F9A48290",
  1270 => x"C0C0C0C0F9A4F8C0",
  1271 => x"C0C0C0C0F9A4F8F9",
  1272 => x"C0C0C0C0F9A4F8A4",
  1273 => x"C0C0C0C0F9A4F8B0",
  1274 => x"C0C0C0C0F9A4F899",
  1275 => x"C0C0C0C0F9A4F892",
  1276 => x"C0C0C0C0F9A4F882",
  1277 => x"C0C0C0C0F9A4F8F8",
  1278 => x"C0C0C0C0F9A4F880",
  1279 => x"C0C0C0C0F9A4F890",
  1280 => x"C0C0C0C0F9A480C0",
  1281 => x"C0C0C0C0F9A480F9",
  1282 => x"C0C0C0C0F9A480A4",
  1283 => x"C0C0C0C0F9A480B0",
  1284 => x"C0C0C0C0F9A48099",
  1285 => x"C0C0C0C0F9A48092",
  1286 => x"C0C0C0C0F9A48082",
  1287 => x"C0C0C0C0F9A480F8",
  1288 => x"C0C0C0C0F9A48080",
  1289 => x"C0C0C0C0F9A48090",
  1290 => x"C0C0C0C0F9A490C0",
  1291 => x"C0C0C0C0F9A490F9",
  1292 => x"C0C0C0C0F9A490A4",
  1293 => x"C0C0C0C0F9A490B0",
  1294 => x"C0C0C0C0F9A49099",
  1295 => x"C0C0C0C0F9A49092",
  1296 => x"C0C0C0C0F9A49082",
  1297 => x"C0C0C0C0F9A490F8",
  1298 => x"C0C0C0C0F9A49080",
  1299 => x"C0C0C0C0F9A49090",
  1300 => x"C0C0C0C0F9B0C0C0",
  1301 => x"C0C0C0C0F9B0C0F9",
  1302 => x"C0C0C0C0F9B0C0A4",
  1303 => x"C0C0C0C0F9B0C0B0",
  1304 => x"C0C0C0C0F9B0C099",
  1305 => x"C0C0C0C0F9B0C092",
  1306 => x"C0C0C0C0F9B0C082",
  1307 => x"C0C0C0C0F9B0C0F8",
  1308 => x"C0C0C0C0F9B0C080",
  1309 => x"C0C0C0C0F9B0C090",
  1310 => x"C0C0C0C0F9B0F9C0",
  1311 => x"C0C0C0C0F9B0F9F9",
  1312 => x"C0C0C0C0F9B0F9A4",
  1313 => x"C0C0C0C0F9B0F9B0",
  1314 => x"C0C0C0C0F9B0F999",
  1315 => x"C0C0C0C0F9B0F992",
  1316 => x"C0C0C0C0F9B0F982",
  1317 => x"C0C0C0C0F9B0F9F8",
  1318 => x"C0C0C0C0F9B0F980",
  1319 => x"C0C0C0C0F9B0F990",
  1320 => x"C0C0C0C0F9B0A4C0",
  1321 => x"C0C0C0C0F9B0A4F9",
  1322 => x"C0C0C0C0F9B0A4A4",
  1323 => x"C0C0C0C0F9B0A4B0",
  1324 => x"C0C0C0C0F9B0A499",
  1325 => x"C0C0C0C0F9B0A492",
  1326 => x"C0C0C0C0F9B0A482",
  1327 => x"C0C0C0C0F9B0A4F8",
  1328 => x"C0C0C0C0F9B0A480",
  1329 => x"C0C0C0C0F9B0A490",
  1330 => x"C0C0C0C0F9B0B0C0",
  1331 => x"C0C0C0C0F9B0B0F9",
  1332 => x"C0C0C0C0F9B0B0A4",
  1333 => x"C0C0C0C0F9B0B0B0",
  1334 => x"C0C0C0C0F9B0B099",
  1335 => x"C0C0C0C0F9B0B092",
  1336 => x"C0C0C0C0F9B0B082",
  1337 => x"C0C0C0C0F9B0B0F8",
  1338 => x"C0C0C0C0F9B0B080",
  1339 => x"C0C0C0C0F9B0B090",
  1340 => x"C0C0C0C0F9B099C0",
  1341 => x"C0C0C0C0F9B099F9",
  1342 => x"C0C0C0C0F9B099A4",
  1343 => x"C0C0C0C0F9B099B0",
  1344 => x"C0C0C0C0F9B09999",
  1345 => x"C0C0C0C0F9B09992",
  1346 => x"C0C0C0C0F9B09982",
  1347 => x"C0C0C0C0F9B099F8",
  1348 => x"C0C0C0C0F9B09980",
  1349 => x"C0C0C0C0F9B09990",
  1350 => x"C0C0C0C0F9B092C0",
  1351 => x"C0C0C0C0F9B092F9",
  1352 => x"C0C0C0C0F9B092A4",
  1353 => x"C0C0C0C0F9B092B0",
  1354 => x"C0C0C0C0F9B09299",
  1355 => x"C0C0C0C0F9B09292",
  1356 => x"C0C0C0C0F9B09282",
  1357 => x"C0C0C0C0F9B092F8",
  1358 => x"C0C0C0C0F9B09280",
  1359 => x"C0C0C0C0F9B09290",
  1360 => x"C0C0C0C0F9B082C0",
  1361 => x"C0C0C0C0F9B082F9",
  1362 => x"C0C0C0C0F9B082A4",
  1363 => x"C0C0C0C0F9B082B0",
  1364 => x"C0C0C0C0F9B08299",
  1365 => x"C0C0C0C0F9B08292",
  1366 => x"C0C0C0C0F9B08282",
  1367 => x"C0C0C0C0F9B082F8",
  1368 => x"C0C0C0C0F9B08280",
  1369 => x"C0C0C0C0F9B08290",
  1370 => x"C0C0C0C0F9B0F8C0",
  1371 => x"C0C0C0C0F9B0F8F9",
  1372 => x"C0C0C0C0F9B0F8A4",
  1373 => x"C0C0C0C0F9B0F8B0",
  1374 => x"C0C0C0C0F9B0F899",
  1375 => x"C0C0C0C0F9B0F892",
  1376 => x"C0C0C0C0F9B0F882",
  1377 => x"C0C0C0C0F9B0F8F8",
  1378 => x"C0C0C0C0F9B0F880",
  1379 => x"C0C0C0C0F9B0F890",
  1380 => x"C0C0C0C0F9B080C0",
  1381 => x"C0C0C0C0F9B080F9",
  1382 => x"C0C0C0C0F9B080A4",
  1383 => x"C0C0C0C0F9B080B0",
  1384 => x"C0C0C0C0F9B08099",
  1385 => x"C0C0C0C0F9B08092",
  1386 => x"C0C0C0C0F9B08082",
  1387 => x"C0C0C0C0F9B080F8",
  1388 => x"C0C0C0C0F9B08080",
  1389 => x"C0C0C0C0F9B08090",
  1390 => x"C0C0C0C0F9B090C0",
  1391 => x"C0C0C0C0F9B090F9",
  1392 => x"C0C0C0C0F9B090A4",
  1393 => x"C0C0C0C0F9B090B0",
  1394 => x"C0C0C0C0F9B09099",
  1395 => x"C0C0C0C0F9B09092",
  1396 => x"C0C0C0C0F9B09082",
  1397 => x"C0C0C0C0F9B090F8",
  1398 => x"C0C0C0C0F9B09080",
  1399 => x"C0C0C0C0F9B09090",
  1400 => x"C0C0C0C0F999C0C0",
  1401 => x"C0C0C0C0F999C0F9",
  1402 => x"C0C0C0C0F999C0A4",
  1403 => x"C0C0C0C0F999C0B0",
  1404 => x"C0C0C0C0F999C099",
  1405 => x"C0C0C0C0F999C092",
  1406 => x"C0C0C0C0F999C082",
  1407 => x"C0C0C0C0F999C0F8",
  1408 => x"C0C0C0C0F999C080",
  1409 => x"C0C0C0C0F999C090",
  1410 => x"C0C0C0C0F999F9C0",
  1411 => x"C0C0C0C0F999F9F9",
  1412 => x"C0C0C0C0F999F9A4",
  1413 => x"C0C0C0C0F999F9B0",
  1414 => x"C0C0C0C0F999F999",
  1415 => x"C0C0C0C0F999F992",
  1416 => x"C0C0C0C0F999F982",
  1417 => x"C0C0C0C0F999F9F8",
  1418 => x"C0C0C0C0F999F980",
  1419 => x"C0C0C0C0F999F990",
  1420 => x"C0C0C0C0F999A4C0",
  1421 => x"C0C0C0C0F999A4F9",
  1422 => x"C0C0C0C0F999A4A4",
  1423 => x"C0C0C0C0F999A4B0",
  1424 => x"C0C0C0C0F999A499",
  1425 => x"C0C0C0C0F999A492",
  1426 => x"C0C0C0C0F999A482",
  1427 => x"C0C0C0C0F999A4F8",
  1428 => x"C0C0C0C0F999A480",
  1429 => x"C0C0C0C0F999A490",
  1430 => x"C0C0C0C0F999B0C0",
  1431 => x"C0C0C0C0F999B0F9",
  1432 => x"C0C0C0C0F999B0A4",
  1433 => x"C0C0C0C0F999B0B0",
  1434 => x"C0C0C0C0F999B099",
  1435 => x"C0C0C0C0F999B092",
  1436 => x"C0C0C0C0F999B082",
  1437 => x"C0C0C0C0F999B0F8",
  1438 => x"C0C0C0C0F999B080",
  1439 => x"C0C0C0C0F999B090",
  1440 => x"C0C0C0C0F99999C0",
  1441 => x"C0C0C0C0F99999F9",
  1442 => x"C0C0C0C0F99999A4",
  1443 => x"C0C0C0C0F99999B0",
  1444 => x"C0C0C0C0F9999999",
  1445 => x"C0C0C0C0F9999992",
  1446 => x"C0C0C0C0F9999982",
  1447 => x"C0C0C0C0F99999F8",
  1448 => x"C0C0C0C0F9999980",
  1449 => x"C0C0C0C0F9999990",
  1450 => x"C0C0C0C0F99992C0",
  1451 => x"C0C0C0C0F99992F9",
  1452 => x"C0C0C0C0F99992A4",
  1453 => x"C0C0C0C0F99992B0",
  1454 => x"C0C0C0C0F9999299",
  1455 => x"C0C0C0C0F9999292",
  1456 => x"C0C0C0C0F9999282",
  1457 => x"C0C0C0C0F99992F8",
  1458 => x"C0C0C0C0F9999280",
  1459 => x"C0C0C0C0F9999290",
  1460 => x"C0C0C0C0F99982C0",
  1461 => x"C0C0C0C0F99982F9",
  1462 => x"C0C0C0C0F99982A4",
  1463 => x"C0C0C0C0F99982B0",
  1464 => x"C0C0C0C0F9998299",
  1465 => x"C0C0C0C0F9998292",
  1466 => x"C0C0C0C0F9998282",
  1467 => x"C0C0C0C0F99982F8",
  1468 => x"C0C0C0C0F9998280",
  1469 => x"C0C0C0C0F9998290",
  1470 => x"C0C0C0C0F999F8C0",
  1471 => x"C0C0C0C0F999F8F9",
  1472 => x"C0C0C0C0F999F8A4",
  1473 => x"C0C0C0C0F999F8B0",
  1474 => x"C0C0C0C0F999F899",
  1475 => x"C0C0C0C0F999F892",
  1476 => x"C0C0C0C0F999F882",
  1477 => x"C0C0C0C0F999F8F8",
  1478 => x"C0C0C0C0F999F880",
  1479 => x"C0C0C0C0F999F890",
  1480 => x"C0C0C0C0F99980C0",
  1481 => x"C0C0C0C0F99980F9",
  1482 => x"C0C0C0C0F99980A4",
  1483 => x"C0C0C0C0F99980B0",
  1484 => x"C0C0C0C0F9998099",
  1485 => x"C0C0C0C0F9998092",
  1486 => x"C0C0C0C0F9998082",
  1487 => x"C0C0C0C0F99980F8",
  1488 => x"C0C0C0C0F9998080",
  1489 => x"C0C0C0C0F9998090",
  1490 => x"C0C0C0C0F99990C0",
  1491 => x"C0C0C0C0F99990F9",
  1492 => x"C0C0C0C0F99990A4",
  1493 => x"C0C0C0C0F99990B0",
  1494 => x"C0C0C0C0F9999099",
  1495 => x"C0C0C0C0F9999092",
  1496 => x"C0C0C0C0F9999082",
  1497 => x"C0C0C0C0F99990F8",
  1498 => x"C0C0C0C0F9999080",
  1499 => x"C0C0C0C0F9999090",
  1500 => x"C0C0C0C0F992C0C0",
  1501 => x"C0C0C0C0F992C0F9",
  1502 => x"C0C0C0C0F992C0A4",
  1503 => x"C0C0C0C0F992C0B0",
  1504 => x"C0C0C0C0F992C099",
  1505 => x"C0C0C0C0F992C092",
  1506 => x"C0C0C0C0F992C082",
  1507 => x"C0C0C0C0F992C0F8",
  1508 => x"C0C0C0C0F992C080",
  1509 => x"C0C0C0C0F992C090",
  1510 => x"C0C0C0C0F992F9C0",
  1511 => x"C0C0C0C0F992F9F9",
  1512 => x"C0C0C0C0F992F9A4",
  1513 => x"C0C0C0C0F992F9B0",
  1514 => x"C0C0C0C0F992F999",
  1515 => x"C0C0C0C0F992F992",
  1516 => x"C0C0C0C0F992F982",
  1517 => x"C0C0C0C0F992F9F8",
  1518 => x"C0C0C0C0F992F980",
  1519 => x"C0C0C0C0F992F990",
  1520 => x"C0C0C0C0F992A4C0",
  1521 => x"C0C0C0C0F992A4F9",
  1522 => x"C0C0C0C0F992A4A4",
  1523 => x"C0C0C0C0F992A4B0",
  1524 => x"C0C0C0C0F992A499",
  1525 => x"C0C0C0C0F992A492",
  1526 => x"C0C0C0C0F992A482",
  1527 => x"C0C0C0C0F992A4F8",
  1528 => x"C0C0C0C0F992A480",
  1529 => x"C0C0C0C0F992A490",
  1530 => x"C0C0C0C0F992B0C0",
  1531 => x"C0C0C0C0F992B0F9",
  1532 => x"C0C0C0C0F992B0A4",
  1533 => x"C0C0C0C0F992B0B0",
  1534 => x"C0C0C0C0F992B099",
  1535 => x"C0C0C0C0F992B092",
  1536 => x"C0C0C0C0F992B082",
  1537 => x"C0C0C0C0F992B0F8",
  1538 => x"C0C0C0C0F992B080",
  1539 => x"C0C0C0C0F992B090",
  1540 => x"C0C0C0C0F99299C0",
  1541 => x"C0C0C0C0F99299F9",
  1542 => x"C0C0C0C0F99299A4",
  1543 => x"C0C0C0C0F99299B0",
  1544 => x"C0C0C0C0F9929999",
  1545 => x"C0C0C0C0F9929992",
  1546 => x"C0C0C0C0F9929982",
  1547 => x"C0C0C0C0F99299F8",
  1548 => x"C0C0C0C0F9929980",
  1549 => x"C0C0C0C0F9929990",
  1550 => x"C0C0C0C0F99292C0",
  1551 => x"C0C0C0C0F99292F9",
  1552 => x"C0C0C0C0F99292A4",
  1553 => x"C0C0C0C0F99292B0",
  1554 => x"C0C0C0C0F9929299",
  1555 => x"C0C0C0C0F9929292",
  1556 => x"C0C0C0C0F9929282",
  1557 => x"C0C0C0C0F99292F8",
  1558 => x"C0C0C0C0F9929280",
  1559 => x"C0C0C0C0F9929290",
  1560 => x"C0C0C0C0F99282C0",
  1561 => x"C0C0C0C0F99282F9",
  1562 => x"C0C0C0C0F99282A4",
  1563 => x"C0C0C0C0F99282B0",
  1564 => x"C0C0C0C0F9928299",
  1565 => x"C0C0C0C0F9928292",
  1566 => x"C0C0C0C0F9928282",
  1567 => x"C0C0C0C0F99282F8",
  1568 => x"C0C0C0C0F9928280",
  1569 => x"C0C0C0C0F9928290",
  1570 => x"C0C0C0C0F992F8C0",
  1571 => x"C0C0C0C0F992F8F9",
  1572 => x"C0C0C0C0F992F8A4",
  1573 => x"C0C0C0C0F992F8B0",
  1574 => x"C0C0C0C0F992F899",
  1575 => x"C0C0C0C0F992F892",
  1576 => x"C0C0C0C0F992F882",
  1577 => x"C0C0C0C0F992F8F8",
  1578 => x"C0C0C0C0F992F880",
  1579 => x"C0C0C0C0F992F890",
  1580 => x"C0C0C0C0F99280C0",
  1581 => x"C0C0C0C0F99280F9",
  1582 => x"C0C0C0C0F99280A4",
  1583 => x"C0C0C0C0F99280B0",
  1584 => x"C0C0C0C0F9928099",
  1585 => x"C0C0C0C0F9928092",
  1586 => x"C0C0C0C0F9928082",
  1587 => x"C0C0C0C0F99280F8",
  1588 => x"C0C0C0C0F9928080",
  1589 => x"C0C0C0C0F9928090",
  1590 => x"C0C0C0C0F99290C0",
  1591 => x"C0C0C0C0F99290F9",
  1592 => x"C0C0C0C0F99290A4",
  1593 => x"C0C0C0C0F99290B0",
  1594 => x"C0C0C0C0F9929099",
  1595 => x"C0C0C0C0F9929092",
  1596 => x"C0C0C0C0F9929082",
  1597 => x"C0C0C0C0F99290F8",
  1598 => x"C0C0C0C0F9929080",
  1599 => x"C0C0C0C0F9929090",
  1600 => x"C0C0C0C0F982C0C0",
  1601 => x"C0C0C0C0F982C0F9",
  1602 => x"C0C0C0C0F982C0A4",
  1603 => x"C0C0C0C0F982C0B0",
  1604 => x"C0C0C0C0F982C099",
  1605 => x"C0C0C0C0F982C092",
  1606 => x"C0C0C0C0F982C082",
  1607 => x"C0C0C0C0F982C0F8",
  1608 => x"C0C0C0C0F982C080",
  1609 => x"C0C0C0C0F982C090",
  1610 => x"C0C0C0C0F982F9C0",
  1611 => x"C0C0C0C0F982F9F9",
  1612 => x"C0C0C0C0F982F9A4",
  1613 => x"C0C0C0C0F982F9B0",
  1614 => x"C0C0C0C0F982F999",
  1615 => x"C0C0C0C0F982F992",
  1616 => x"C0C0C0C0F982F982",
  1617 => x"C0C0C0C0F982F9F8",
  1618 => x"C0C0C0C0F982F980",
  1619 => x"C0C0C0C0F982F990",
  1620 => x"C0C0C0C0F982A4C0",
  1621 => x"C0C0C0C0F982A4F9",
  1622 => x"C0C0C0C0F982A4A4",
  1623 => x"C0C0C0C0F982A4B0",
  1624 => x"C0C0C0C0F982A499",
  1625 => x"C0C0C0C0F982A492",
  1626 => x"C0C0C0C0F982A482",
  1627 => x"C0C0C0C0F982A4F8",
  1628 => x"C0C0C0C0F982A480",
  1629 => x"C0C0C0C0F982A490",
  1630 => x"C0C0C0C0F982B0C0",
  1631 => x"C0C0C0C0F982B0F9",
  1632 => x"C0C0C0C0F982B0A4",
  1633 => x"C0C0C0C0F982B0B0",
  1634 => x"C0C0C0C0F982B099",
  1635 => x"C0C0C0C0F982B092",
  1636 => x"C0C0C0C0F982B082",
  1637 => x"C0C0C0C0F982B0F8",
  1638 => x"C0C0C0C0F982B080",
  1639 => x"C0C0C0C0F982B090",
  1640 => x"C0C0C0C0F98299C0",
  1641 => x"C0C0C0C0F98299F9",
  1642 => x"C0C0C0C0F98299A4",
  1643 => x"C0C0C0C0F98299B0",
  1644 => x"C0C0C0C0F9829999",
  1645 => x"C0C0C0C0F9829992",
  1646 => x"C0C0C0C0F9829982",
  1647 => x"C0C0C0C0F98299F8",
  1648 => x"C0C0C0C0F9829980",
  1649 => x"C0C0C0C0F9829990",
  1650 => x"C0C0C0C0F98292C0",
  1651 => x"C0C0C0C0F98292F9",
  1652 => x"C0C0C0C0F98292A4",
  1653 => x"C0C0C0C0F98292B0",
  1654 => x"C0C0C0C0F9829299",
  1655 => x"C0C0C0C0F9829292",
  1656 => x"C0C0C0C0F9829282",
  1657 => x"C0C0C0C0F98292F8",
  1658 => x"C0C0C0C0F9829280",
  1659 => x"C0C0C0C0F9829290",
  1660 => x"C0C0C0C0F98282C0",
  1661 => x"C0C0C0C0F98282F9",
  1662 => x"C0C0C0C0F98282A4",
  1663 => x"C0C0C0C0F98282B0",
  1664 => x"C0C0C0C0F9828299",
  1665 => x"C0C0C0C0F9828292",
  1666 => x"C0C0C0C0F9828282",
  1667 => x"C0C0C0C0F98282F8",
  1668 => x"C0C0C0C0F9828280",
  1669 => x"C0C0C0C0F9828290",
  1670 => x"C0C0C0C0F982F8C0",
  1671 => x"C0C0C0C0F982F8F9",
  1672 => x"C0C0C0C0F982F8A4",
  1673 => x"C0C0C0C0F982F8B0",
  1674 => x"C0C0C0C0F982F899",
  1675 => x"C0C0C0C0F982F892",
  1676 => x"C0C0C0C0F982F882",
  1677 => x"C0C0C0C0F982F8F8",
  1678 => x"C0C0C0C0F982F880",
  1679 => x"C0C0C0C0F982F890",
  1680 => x"C0C0C0C0F98280C0",
  1681 => x"C0C0C0C0F98280F9",
  1682 => x"C0C0C0C0F98280A4",
  1683 => x"C0C0C0C0F98280B0",
  1684 => x"C0C0C0C0F9828099",
  1685 => x"C0C0C0C0F9828092",
  1686 => x"C0C0C0C0F9828082",
  1687 => x"C0C0C0C0F98280F8",
  1688 => x"C0C0C0C0F9828080",
  1689 => x"C0C0C0C0F9828090",
  1690 => x"C0C0C0C0F98290C0",
  1691 => x"C0C0C0C0F98290F9",
  1692 => x"C0C0C0C0F98290A4",
  1693 => x"C0C0C0C0F98290B0",
  1694 => x"C0C0C0C0F9829099",
  1695 => x"C0C0C0C0F9829092",
  1696 => x"C0C0C0C0F9829082",
  1697 => x"C0C0C0C0F98290F8",
  1698 => x"C0C0C0C0F9829080",
  1699 => x"C0C0C0C0F9829090",
  1700 => x"C0C0C0C0F9F8C0C0",
  1701 => x"C0C0C0C0F9F8C0F9",
  1702 => x"C0C0C0C0F9F8C0A4",
  1703 => x"C0C0C0C0F9F8C0B0",
  1704 => x"C0C0C0C0F9F8C099",
  1705 => x"C0C0C0C0F9F8C092",
  1706 => x"C0C0C0C0F9F8C082",
  1707 => x"C0C0C0C0F9F8C0F8",
  1708 => x"C0C0C0C0F9F8C080",
  1709 => x"C0C0C0C0F9F8C090",
  1710 => x"C0C0C0C0F9F8F9C0",
  1711 => x"C0C0C0C0F9F8F9F9",
  1712 => x"C0C0C0C0F9F8F9A4",
  1713 => x"C0C0C0C0F9F8F9B0",
  1714 => x"C0C0C0C0F9F8F999",
  1715 => x"C0C0C0C0F9F8F992",
  1716 => x"C0C0C0C0F9F8F982",
  1717 => x"C0C0C0C0F9F8F9F8",
  1718 => x"C0C0C0C0F9F8F980",
  1719 => x"C0C0C0C0F9F8F990",
  1720 => x"C0C0C0C0F9F8A4C0",
  1721 => x"C0C0C0C0F9F8A4F9",
  1722 => x"C0C0C0C0F9F8A4A4",
  1723 => x"C0C0C0C0F9F8A4B0",
  1724 => x"C0C0C0C0F9F8A499",
  1725 => x"C0C0C0C0F9F8A492",
  1726 => x"C0C0C0C0F9F8A482",
  1727 => x"C0C0C0C0F9F8A4F8",
  1728 => x"C0C0C0C0F9F8A480",
  1729 => x"C0C0C0C0F9F8A490",
  1730 => x"C0C0C0C0F9F8B0C0",
  1731 => x"C0C0C0C0F9F8B0F9",
  1732 => x"C0C0C0C0F9F8B0A4",
  1733 => x"C0C0C0C0F9F8B0B0",
  1734 => x"C0C0C0C0F9F8B099",
  1735 => x"C0C0C0C0F9F8B092",
  1736 => x"C0C0C0C0F9F8B082",
  1737 => x"C0C0C0C0F9F8B0F8",
  1738 => x"C0C0C0C0F9F8B080",
  1739 => x"C0C0C0C0F9F8B090",
  1740 => x"C0C0C0C0F9F899C0",
  1741 => x"C0C0C0C0F9F899F9",
  1742 => x"C0C0C0C0F9F899A4",
  1743 => x"C0C0C0C0F9F899B0",
  1744 => x"C0C0C0C0F9F89999",
  1745 => x"C0C0C0C0F9F89992",
  1746 => x"C0C0C0C0F9F89982",
  1747 => x"C0C0C0C0F9F899F8",
  1748 => x"C0C0C0C0F9F89980",
  1749 => x"C0C0C0C0F9F89990",
  1750 => x"C0C0C0C0F9F892C0",
  1751 => x"C0C0C0C0F9F892F9",
  1752 => x"C0C0C0C0F9F892A4",
  1753 => x"C0C0C0C0F9F892B0",
  1754 => x"C0C0C0C0F9F89299",
  1755 => x"C0C0C0C0F9F89292",
  1756 => x"C0C0C0C0F9F89282",
  1757 => x"C0C0C0C0F9F892F8",
  1758 => x"C0C0C0C0F9F89280",
  1759 => x"C0C0C0C0F9F89290",
  1760 => x"C0C0C0C0F9F882C0",
  1761 => x"C0C0C0C0F9F882F9",
  1762 => x"C0C0C0C0F9F882A4",
  1763 => x"C0C0C0C0F9F882B0",
  1764 => x"C0C0C0C0F9F88299",
  1765 => x"C0C0C0C0F9F88292",
  1766 => x"C0C0C0C0F9F88282",
  1767 => x"C0C0C0C0F9F882F8",
  1768 => x"C0C0C0C0F9F88280",
  1769 => x"C0C0C0C0F9F88290",
  1770 => x"C0C0C0C0F9F8F8C0",
  1771 => x"C0C0C0C0F9F8F8F9",
  1772 => x"C0C0C0C0F9F8F8A4",
  1773 => x"C0C0C0C0F9F8F8B0",
  1774 => x"C0C0C0C0F9F8F899",
  1775 => x"C0C0C0C0F9F8F892",
  1776 => x"C0C0C0C0F9F8F882",
  1777 => x"C0C0C0C0F9F8F8F8",
  1778 => x"C0C0C0C0F9F8F880",
  1779 => x"C0C0C0C0F9F8F890",
  1780 => x"C0C0C0C0F9F880C0",
  1781 => x"C0C0C0C0F9F880F9",
  1782 => x"C0C0C0C0F9F880A4",
  1783 => x"C0C0C0C0F9F880B0",
  1784 => x"C0C0C0C0F9F88099",
  1785 => x"C0C0C0C0F9F88092",
  1786 => x"C0C0C0C0F9F88082",
  1787 => x"C0C0C0C0F9F880F8",
  1788 => x"C0C0C0C0F9F88080",
  1789 => x"C0C0C0C0F9F88090",
  1790 => x"C0C0C0C0F9F890C0",
  1791 => x"C0C0C0C0F9F890F9",
  1792 => x"C0C0C0C0F9F890A4",
  1793 => x"C0C0C0C0F9F890B0",
  1794 => x"C0C0C0C0F9F89099",
  1795 => x"C0C0C0C0F9F89092",
  1796 => x"C0C0C0C0F9F89082",
  1797 => x"C0C0C0C0F9F890F8",
  1798 => x"C0C0C0C0F9F89080",
  1799 => x"C0C0C0C0F9F89090",
  1800 => x"C0C0C0C0F980C0C0",
  1801 => x"C0C0C0C0F980C0F9",
  1802 => x"C0C0C0C0F980C0A4",
  1803 => x"C0C0C0C0F980C0B0",
  1804 => x"C0C0C0C0F980C099",
  1805 => x"C0C0C0C0F980C092",
  1806 => x"C0C0C0C0F980C082",
  1807 => x"C0C0C0C0F980C0F8",
  1808 => x"C0C0C0C0F980C080",
  1809 => x"C0C0C0C0F980C090",
  1810 => x"C0C0C0C0F980F9C0",
  1811 => x"C0C0C0C0F980F9F9",
  1812 => x"C0C0C0C0F980F9A4",
  1813 => x"C0C0C0C0F980F9B0",
  1814 => x"C0C0C0C0F980F999",
  1815 => x"C0C0C0C0F980F992",
  1816 => x"C0C0C0C0F980F982",
  1817 => x"C0C0C0C0F980F9F8",
  1818 => x"C0C0C0C0F980F980",
  1819 => x"C0C0C0C0F980F990",
  1820 => x"C0C0C0C0F980A4C0",
  1821 => x"C0C0C0C0F980A4F9",
  1822 => x"C0C0C0C0F980A4A4",
  1823 => x"C0C0C0C0F980A4B0",
  1824 => x"C0C0C0C0F980A499",
  1825 => x"C0C0C0C0F980A492",
  1826 => x"C0C0C0C0F980A482",
  1827 => x"C0C0C0C0F980A4F8",
  1828 => x"C0C0C0C0F980A480",
  1829 => x"C0C0C0C0F980A490",
  1830 => x"C0C0C0C0F980B0C0",
  1831 => x"C0C0C0C0F980B0F9",
  1832 => x"C0C0C0C0F980B0A4",
  1833 => x"C0C0C0C0F980B0B0",
  1834 => x"C0C0C0C0F980B099",
  1835 => x"C0C0C0C0F980B092",
  1836 => x"C0C0C0C0F980B082",
  1837 => x"C0C0C0C0F980B0F8",
  1838 => x"C0C0C0C0F980B080",
  1839 => x"C0C0C0C0F980B090",
  1840 => x"C0C0C0C0F98099C0",
  1841 => x"C0C0C0C0F98099F9",
  1842 => x"C0C0C0C0F98099A4",
  1843 => x"C0C0C0C0F98099B0",
  1844 => x"C0C0C0C0F9809999",
  1845 => x"C0C0C0C0F9809992",
  1846 => x"C0C0C0C0F9809982",
  1847 => x"C0C0C0C0F98099F8",
  1848 => x"C0C0C0C0F9809980",
  1849 => x"C0C0C0C0F9809990",
  1850 => x"C0C0C0C0F98092C0",
  1851 => x"C0C0C0C0F98092F9",
  1852 => x"C0C0C0C0F98092A4",
  1853 => x"C0C0C0C0F98092B0",
  1854 => x"C0C0C0C0F9809299",
  1855 => x"C0C0C0C0F9809292",
  1856 => x"C0C0C0C0F9809282",
  1857 => x"C0C0C0C0F98092F8",
  1858 => x"C0C0C0C0F9809280",
  1859 => x"C0C0C0C0F9809290",
  1860 => x"C0C0C0C0F98082C0",
  1861 => x"C0C0C0C0F98082F9",
  1862 => x"C0C0C0C0F98082A4",
  1863 => x"C0C0C0C0F98082B0",
  1864 => x"C0C0C0C0F9808299",
  1865 => x"C0C0C0C0F9808292",
  1866 => x"C0C0C0C0F9808282",
  1867 => x"C0C0C0C0F98082F8",
  1868 => x"C0C0C0C0F9808280",
  1869 => x"C0C0C0C0F9808290",
  1870 => x"C0C0C0C0F980F8C0",
  1871 => x"C0C0C0C0F980F8F9",
  1872 => x"C0C0C0C0F980F8A4",
  1873 => x"C0C0C0C0F980F8B0",
  1874 => x"C0C0C0C0F980F899",
  1875 => x"C0C0C0C0F980F892",
  1876 => x"C0C0C0C0F980F882",
  1877 => x"C0C0C0C0F980F8F8",
  1878 => x"C0C0C0C0F980F880",
  1879 => x"C0C0C0C0F980F890",
  1880 => x"C0C0C0C0F98080C0",
  1881 => x"C0C0C0C0F98080F9",
  1882 => x"C0C0C0C0F98080A4",
  1883 => x"C0C0C0C0F98080B0",
  1884 => x"C0C0C0C0F9808099",
  1885 => x"C0C0C0C0F9808092",
  1886 => x"C0C0C0C0F9808082",
  1887 => x"C0C0C0C0F98080F8",
  1888 => x"C0C0C0C0F9808080",
  1889 => x"C0C0C0C0F9808090",
  1890 => x"C0C0C0C0F98090C0",
  1891 => x"C0C0C0C0F98090F9",
  1892 => x"C0C0C0C0F98090A4",
  1893 => x"C0C0C0C0F98090B0",
  1894 => x"C0C0C0C0F9809099",
  1895 => x"C0C0C0C0F9809092",
  1896 => x"C0C0C0C0F9809082",
  1897 => x"C0C0C0C0F98090F8",
  1898 => x"C0C0C0C0F9809080",
  1899 => x"C0C0C0C0F9809090",
  1900 => x"C0C0C0C0F990C0C0",
  1901 => x"C0C0C0C0F990C0F9",
  1902 => x"C0C0C0C0F990C0A4",
  1903 => x"C0C0C0C0F990C0B0",
  1904 => x"C0C0C0C0F990C099",
  1905 => x"C0C0C0C0F990C092",
  1906 => x"C0C0C0C0F990C082",
  1907 => x"C0C0C0C0F990C0F8",
  1908 => x"C0C0C0C0F990C080",
  1909 => x"C0C0C0C0F990C090",
  1910 => x"C0C0C0C0F990F9C0",
  1911 => x"C0C0C0C0F990F9F9",
  1912 => x"C0C0C0C0F990F9A4",
  1913 => x"C0C0C0C0F990F9B0",
  1914 => x"C0C0C0C0F990F999",
  1915 => x"C0C0C0C0F990F992",
  1916 => x"C0C0C0C0F990F982",
  1917 => x"C0C0C0C0F990F9F8",
  1918 => x"C0C0C0C0F990F980",
  1919 => x"C0C0C0C0F990F990",
  1920 => x"C0C0C0C0F990A4C0",
  1921 => x"C0C0C0C0F990A4F9",
  1922 => x"C0C0C0C0F990A4A4",
  1923 => x"C0C0C0C0F990A4B0",
  1924 => x"C0C0C0C0F990A499",
  1925 => x"C0C0C0C0F990A492",
  1926 => x"C0C0C0C0F990A482",
  1927 => x"C0C0C0C0F990A4F8",
  1928 => x"C0C0C0C0F990A480",
  1929 => x"C0C0C0C0F990A490",
  1930 => x"C0C0C0C0F990B0C0",
  1931 => x"C0C0C0C0F990B0F9",
  1932 => x"C0C0C0C0F990B0A4",
  1933 => x"C0C0C0C0F990B0B0",
  1934 => x"C0C0C0C0F990B099",
  1935 => x"C0C0C0C0F990B092",
  1936 => x"C0C0C0C0F990B082",
  1937 => x"C0C0C0C0F990B0F8",
  1938 => x"C0C0C0C0F990B080",
  1939 => x"C0C0C0C0F990B090",
  1940 => x"C0C0C0C0F99099C0",
  1941 => x"C0C0C0C0F99099F9",
  1942 => x"C0C0C0C0F99099A4",
  1943 => x"C0C0C0C0F99099B0",
  1944 => x"C0C0C0C0F9909999",
  1945 => x"C0C0C0C0F9909992",
  1946 => x"C0C0C0C0F9909982",
  1947 => x"C0C0C0C0F99099F8",
  1948 => x"C0C0C0C0F9909980",
  1949 => x"C0C0C0C0F9909990",
  1950 => x"C0C0C0C0F99092C0",
  1951 => x"C0C0C0C0F99092F9",
  1952 => x"C0C0C0C0F99092A4",
  1953 => x"C0C0C0C0F99092B0",
  1954 => x"C0C0C0C0F9909299",
  1955 => x"C0C0C0C0F9909292",
  1956 => x"C0C0C0C0F9909282",
  1957 => x"C0C0C0C0F99092F8",
  1958 => x"C0C0C0C0F9909280",
  1959 => x"C0C0C0C0F9909290",
  1960 => x"C0C0C0C0F99082C0",
  1961 => x"C0C0C0C0F99082F9",
  1962 => x"C0C0C0C0F99082A4",
  1963 => x"C0C0C0C0F99082B0",
  1964 => x"C0C0C0C0F9908299",
  1965 => x"C0C0C0C0F9908292",
  1966 => x"C0C0C0C0F9908282",
  1967 => x"C0C0C0C0F99082F8",
  1968 => x"C0C0C0C0F9908280",
  1969 => x"C0C0C0C0F9908290",
  1970 => x"C0C0C0C0F990F8C0",
  1971 => x"C0C0C0C0F990F8F9",
  1972 => x"C0C0C0C0F990F8A4",
  1973 => x"C0C0C0C0F990F8B0",
  1974 => x"C0C0C0C0F990F899",
  1975 => x"C0C0C0C0F990F892",
  1976 => x"C0C0C0C0F990F882",
  1977 => x"C0C0C0C0F990F8F8",
  1978 => x"C0C0C0C0F990F880",
  1979 => x"C0C0C0C0F990F890",
  1980 => x"C0C0C0C0F99080C0",
  1981 => x"C0C0C0C0F99080F9",
  1982 => x"C0C0C0C0F99080A4",
  1983 => x"C0C0C0C0F99080B0",
  1984 => x"C0C0C0C0F9908099",
  1985 => x"C0C0C0C0F9908092",
  1986 => x"C0C0C0C0F9908082",
  1987 => x"C0C0C0C0F99080F8",
  1988 => x"C0C0C0C0F9908080",
  1989 => x"C0C0C0C0F9908090",
  1990 => x"C0C0C0C0F99090C0",
  1991 => x"C0C0C0C0F99090F9",
  1992 => x"C0C0C0C0F99090A4",
  1993 => x"C0C0C0C0F99090B0",
  1994 => x"C0C0C0C0F9909099",
  1995 => x"C0C0C0C0F9909092",
  1996 => x"C0C0C0C0F9909082",
  1997 => x"C0C0C0C0F99090F8",
  1998 => x"C0C0C0C0F9909080",
  1999 => x"C0C0C0C0F9909090",
  2000 => x"C0C0C0C0A4C0C0C0",
  2001 => x"C0C0C0C0A4C0C0F9",
  2002 => x"C0C0C0C0A4C0C0A4",
  2003 => x"C0C0C0C0A4C0C0B0",
  2004 => x"C0C0C0C0A4C0C099",
  2005 => x"C0C0C0C0A4C0C092",
  2006 => x"C0C0C0C0A4C0C082",
  2007 => x"C0C0C0C0A4C0C0F8",
  2008 => x"C0C0C0C0A4C0C080",
  2009 => x"C0C0C0C0A4C0C090",
  2010 => x"C0C0C0C0A4C0F9C0",
  2011 => x"C0C0C0C0A4C0F9F9",
  2012 => x"C0C0C0C0A4C0F9A4",
  2013 => x"C0C0C0C0A4C0F9B0",
  2014 => x"C0C0C0C0A4C0F999",
  2015 => x"C0C0C0C0A4C0F992",
  2016 => x"C0C0C0C0A4C0F982",
  2017 => x"C0C0C0C0A4C0F9F8",
  2018 => x"C0C0C0C0A4C0F980",
  2019 => x"C0C0C0C0A4C0F990",
  2020 => x"C0C0C0C0A4C0A4C0",
  2021 => x"C0C0C0C0A4C0A4F9",
  2022 => x"C0C0C0C0A4C0A4A4",
  2023 => x"C0C0C0C0A4C0A4B0",
  2024 => x"C0C0C0C0A4C0A499",
  2025 => x"C0C0C0C0A4C0A492",
  2026 => x"C0C0C0C0A4C0A482",
  2027 => x"C0C0C0C0A4C0A4F8",
  2028 => x"C0C0C0C0A4C0A480",
  2029 => x"C0C0C0C0A4C0A490",
  2030 => x"C0C0C0C0A4C0B0C0",
  2031 => x"C0C0C0C0A4C0B0F9",
  2032 => x"C0C0C0C0A4C0B0A4",
  2033 => x"C0C0C0C0A4C0B0B0",
  2034 => x"C0C0C0C0A4C0B099",
  2035 => x"C0C0C0C0A4C0B092",
  2036 => x"C0C0C0C0A4C0B082",
  2037 => x"C0C0C0C0A4C0B0F8",
  2038 => x"C0C0C0C0A4C0B080",
  2039 => x"C0C0C0C0A4C0B090",
  2040 => x"C0C0C0C0A4C099C0",
  2041 => x"C0C0C0C0A4C099F9",
  2042 => x"C0C0C0C0A4C099A4",
  2043 => x"C0C0C0C0A4C099B0",
  2044 => x"C0C0C0C0A4C09999",
  2045 => x"C0C0C0C0A4C09992",
  2046 => x"C0C0C0C0A4C09982",
  2047 => x"C0C0C0C0A4C099F8",
  2048 => x"C0C0C0C0A4C09980",
  2049 => x"C0C0C0C0A4C09990",
  2050 => x"C0C0C0C0A4C092C0",
  2051 => x"C0C0C0C0A4C092F9",
  2052 => x"C0C0C0C0A4C092A4",
  2053 => x"C0C0C0C0A4C092B0",
  2054 => x"C0C0C0C0A4C09299",
  2055 => x"C0C0C0C0A4C09292",
  2056 => x"C0C0C0C0A4C09282",
  2057 => x"C0C0C0C0A4C092F8",
  2058 => x"C0C0C0C0A4C09280",
  2059 => x"C0C0C0C0A4C09290",
  2060 => x"C0C0C0C0A4C082C0",
  2061 => x"C0C0C0C0A4C082F9",
  2062 => x"C0C0C0C0A4C082A4",
  2063 => x"C0C0C0C0A4C082B0",
  2064 => x"C0C0C0C0A4C08299",
  2065 => x"C0C0C0C0A4C08292",
  2066 => x"C0C0C0C0A4C08282",
  2067 => x"C0C0C0C0A4C082F8",
  2068 => x"C0C0C0C0A4C08280",
  2069 => x"C0C0C0C0A4C08290",
  2070 => x"C0C0C0C0A4C0F8C0",
  2071 => x"C0C0C0C0A4C0F8F9",
  2072 => x"C0C0C0C0A4C0F8A4",
  2073 => x"C0C0C0C0A4C0F8B0",
  2074 => x"C0C0C0C0A4C0F899",
  2075 => x"C0C0C0C0A4C0F892",
  2076 => x"C0C0C0C0A4C0F882",
  2077 => x"C0C0C0C0A4C0F8F8",
  2078 => x"C0C0C0C0A4C0F880",
  2079 => x"C0C0C0C0A4C0F890",
  2080 => x"C0C0C0C0A4C080C0",
  2081 => x"C0C0C0C0A4C080F9",
  2082 => x"C0C0C0C0A4C080A4",
  2083 => x"C0C0C0C0A4C080B0",
  2084 => x"C0C0C0C0A4C08099",
  2085 => x"C0C0C0C0A4C08092",
  2086 => x"C0C0C0C0A4C08082",
  2087 => x"C0C0C0C0A4C080F8",
  2088 => x"C0C0C0C0A4C08080",
  2089 => x"C0C0C0C0A4C08090",
  2090 => x"C0C0C0C0A4C090C0",
  2091 => x"C0C0C0C0A4C090F9",
  2092 => x"C0C0C0C0A4C090A4",
  2093 => x"C0C0C0C0A4C090B0",
  2094 => x"C0C0C0C0A4C09099",
  2095 => x"C0C0C0C0A4C09092",
  2096 => x"C0C0C0C0A4C09082",
  2097 => x"C0C0C0C0A4C090F8",
  2098 => x"C0C0C0C0A4C09080",
  2099 => x"C0C0C0C0A4C09090",
  2100 => x"C0C0C0C0A4F9C0C0",
  2101 => x"C0C0C0C0A4F9C0F9",
  2102 => x"C0C0C0C0A4F9C0A4",
  2103 => x"C0C0C0C0A4F9C0B0",
  2104 => x"C0C0C0C0A4F9C099",
  2105 => x"C0C0C0C0A4F9C092",
  2106 => x"C0C0C0C0A4F9C082",
  2107 => x"C0C0C0C0A4F9C0F8",
  2108 => x"C0C0C0C0A4F9C080",
  2109 => x"C0C0C0C0A4F9C090",
  2110 => x"C0C0C0C0A4F9F9C0",
  2111 => x"C0C0C0C0A4F9F9F9",
  2112 => x"C0C0C0C0A4F9F9A4",
  2113 => x"C0C0C0C0A4F9F9B0",
  2114 => x"C0C0C0C0A4F9F999",
  2115 => x"C0C0C0C0A4F9F992",
  2116 => x"C0C0C0C0A4F9F982",
  2117 => x"C0C0C0C0A4F9F9F8",
  2118 => x"C0C0C0C0A4F9F980",
  2119 => x"C0C0C0C0A4F9F990",
  2120 => x"C0C0C0C0A4F9A4C0",
  2121 => x"C0C0C0C0A4F9A4F9",
  2122 => x"C0C0C0C0A4F9A4A4",
  2123 => x"C0C0C0C0A4F9A4B0",
  2124 => x"C0C0C0C0A4F9A499",
  2125 => x"C0C0C0C0A4F9A492",
  2126 => x"C0C0C0C0A4F9A482",
  2127 => x"C0C0C0C0A4F9A4F8",
  2128 => x"C0C0C0C0A4F9A480",
  2129 => x"C0C0C0C0A4F9A490",
  2130 => x"C0C0C0C0A4F9B0C0",
  2131 => x"C0C0C0C0A4F9B0F9",
  2132 => x"C0C0C0C0A4F9B0A4",
  2133 => x"C0C0C0C0A4F9B0B0",
  2134 => x"C0C0C0C0A4F9B099",
  2135 => x"C0C0C0C0A4F9B092",
  2136 => x"C0C0C0C0A4F9B082",
  2137 => x"C0C0C0C0A4F9B0F8",
  2138 => x"C0C0C0C0A4F9B080",
  2139 => x"C0C0C0C0A4F9B090",
  2140 => x"C0C0C0C0A4F999C0",
  2141 => x"C0C0C0C0A4F999F9",
  2142 => x"C0C0C0C0A4F999A4",
  2143 => x"C0C0C0C0A4F999B0",
  2144 => x"C0C0C0C0A4F99999",
  2145 => x"C0C0C0C0A4F99992",
  2146 => x"C0C0C0C0A4F99982",
  2147 => x"C0C0C0C0A4F999F8",
  2148 => x"C0C0C0C0A4F99980",
  2149 => x"C0C0C0C0A4F99990",
  2150 => x"C0C0C0C0A4F992C0",
  2151 => x"C0C0C0C0A4F992F9",
  2152 => x"C0C0C0C0A4F992A4",
  2153 => x"C0C0C0C0A4F992B0",
  2154 => x"C0C0C0C0A4F99299",
  2155 => x"C0C0C0C0A4F99292",
  2156 => x"C0C0C0C0A4F99282",
  2157 => x"C0C0C0C0A4F992F8",
  2158 => x"C0C0C0C0A4F99280",
  2159 => x"C0C0C0C0A4F99290",
  2160 => x"C0C0C0C0A4F982C0",
  2161 => x"C0C0C0C0A4F982F9",
  2162 => x"C0C0C0C0A4F982A4",
  2163 => x"C0C0C0C0A4F982B0",
  2164 => x"C0C0C0C0A4F98299",
  2165 => x"C0C0C0C0A4F98292",
  2166 => x"C0C0C0C0A4F98282",
  2167 => x"C0C0C0C0A4F982F8",
  2168 => x"C0C0C0C0A4F98280",
  2169 => x"C0C0C0C0A4F98290",
  2170 => x"C0C0C0C0A4F9F8C0",
  2171 => x"C0C0C0C0A4F9F8F9",
  2172 => x"C0C0C0C0A4F9F8A4",
  2173 => x"C0C0C0C0A4F9F8B0",
  2174 => x"C0C0C0C0A4F9F899",
  2175 => x"C0C0C0C0A4F9F892",
  2176 => x"C0C0C0C0A4F9F882",
  2177 => x"C0C0C0C0A4F9F8F8",
  2178 => x"C0C0C0C0A4F9F880",
  2179 => x"C0C0C0C0A4F9F890",
  2180 => x"C0C0C0C0A4F980C0",
  2181 => x"C0C0C0C0A4F980F9",
  2182 => x"C0C0C0C0A4F980A4",
  2183 => x"C0C0C0C0A4F980B0",
  2184 => x"C0C0C0C0A4F98099",
  2185 => x"C0C0C0C0A4F98092",
  2186 => x"C0C0C0C0A4F98082",
  2187 => x"C0C0C0C0A4F980F8",
  2188 => x"C0C0C0C0A4F98080",
  2189 => x"C0C0C0C0A4F98090",
  2190 => x"C0C0C0C0A4F990C0",
  2191 => x"C0C0C0C0A4F990F9",
  2192 => x"C0C0C0C0A4F990A4",
  2193 => x"C0C0C0C0A4F990B0",
  2194 => x"C0C0C0C0A4F99099",
  2195 => x"C0C0C0C0A4F99092",
  2196 => x"C0C0C0C0A4F99082",
  2197 => x"C0C0C0C0A4F990F8",
  2198 => x"C0C0C0C0A4F99080",
  2199 => x"C0C0C0C0A4F99090",
  2200 => x"C0C0C0C0A4A4C0C0",
  2201 => x"C0C0C0C0A4A4C0F9",
  2202 => x"C0C0C0C0A4A4C0A4",
  2203 => x"C0C0C0C0A4A4C0B0",
  2204 => x"C0C0C0C0A4A4C099",
  2205 => x"C0C0C0C0A4A4C092",
  2206 => x"C0C0C0C0A4A4C082",
  2207 => x"C0C0C0C0A4A4C0F8",
  2208 => x"C0C0C0C0A4A4C080",
  2209 => x"C0C0C0C0A4A4C090",
  2210 => x"C0C0C0C0A4A4F9C0",
  2211 => x"C0C0C0C0A4A4F9F9",
  2212 => x"C0C0C0C0A4A4F9A4",
  2213 => x"C0C0C0C0A4A4F9B0",
  2214 => x"C0C0C0C0A4A4F999",
  2215 => x"C0C0C0C0A4A4F992",
  2216 => x"C0C0C0C0A4A4F982",
  2217 => x"C0C0C0C0A4A4F9F8",
  2218 => x"C0C0C0C0A4A4F980",
  2219 => x"C0C0C0C0A4A4F990",
  2220 => x"C0C0C0C0A4A4A4C0",
  2221 => x"C0C0C0C0A4A4A4F9",
  2222 => x"C0C0C0C0A4A4A4A4",
  2223 => x"C0C0C0C0A4A4A4B0",
  2224 => x"C0C0C0C0A4A4A499",
  2225 => x"C0C0C0C0A4A4A492",
  2226 => x"C0C0C0C0A4A4A482",
  2227 => x"C0C0C0C0A4A4A4F8",
  2228 => x"C0C0C0C0A4A4A480",
  2229 => x"C0C0C0C0A4A4A490",
  2230 => x"C0C0C0C0A4A4B0C0",
  2231 => x"C0C0C0C0A4A4B0F9",
  2232 => x"C0C0C0C0A4A4B0A4",
  2233 => x"C0C0C0C0A4A4B0B0",
  2234 => x"C0C0C0C0A4A4B099",
  2235 => x"C0C0C0C0A4A4B092",
  2236 => x"C0C0C0C0A4A4B082",
  2237 => x"C0C0C0C0A4A4B0F8",
  2238 => x"C0C0C0C0A4A4B080",
  2239 => x"C0C0C0C0A4A4B090",
  2240 => x"C0C0C0C0A4A499C0",
  2241 => x"C0C0C0C0A4A499F9",
  2242 => x"C0C0C0C0A4A499A4",
  2243 => x"C0C0C0C0A4A499B0",
  2244 => x"C0C0C0C0A4A49999",
  2245 => x"C0C0C0C0A4A49992",
  2246 => x"C0C0C0C0A4A49982",
  2247 => x"C0C0C0C0A4A499F8",
  2248 => x"C0C0C0C0A4A49980",
  2249 => x"C0C0C0C0A4A49990",
  2250 => x"C0C0C0C0A4A492C0",
  2251 => x"C0C0C0C0A4A492F9",
  2252 => x"C0C0C0C0A4A492A4",
  2253 => x"C0C0C0C0A4A492B0",
  2254 => x"C0C0C0C0A4A49299",
  2255 => x"C0C0C0C0A4A49292",
  2256 => x"C0C0C0C0A4A49282",
  2257 => x"C0C0C0C0A4A492F8",
  2258 => x"C0C0C0C0A4A49280",
  2259 => x"C0C0C0C0A4A49290",
  2260 => x"C0C0C0C0A4A482C0",
  2261 => x"C0C0C0C0A4A482F9",
  2262 => x"C0C0C0C0A4A482A4",
  2263 => x"C0C0C0C0A4A482B0",
  2264 => x"C0C0C0C0A4A48299",
  2265 => x"C0C0C0C0A4A48292",
  2266 => x"C0C0C0C0A4A48282",
  2267 => x"C0C0C0C0A4A482F8",
  2268 => x"C0C0C0C0A4A48280",
  2269 => x"C0C0C0C0A4A48290",
  2270 => x"C0C0C0C0A4A4F8C0",
  2271 => x"C0C0C0C0A4A4F8F9",
  2272 => x"C0C0C0C0A4A4F8A4",
  2273 => x"C0C0C0C0A4A4F8B0",
  2274 => x"C0C0C0C0A4A4F899",
  2275 => x"C0C0C0C0A4A4F892",
  2276 => x"C0C0C0C0A4A4F882",
  2277 => x"C0C0C0C0A4A4F8F8",
  2278 => x"C0C0C0C0A4A4F880",
  2279 => x"C0C0C0C0A4A4F890",
  2280 => x"C0C0C0C0A4A480C0",
  2281 => x"C0C0C0C0A4A480F9",
  2282 => x"C0C0C0C0A4A480A4",
  2283 => x"C0C0C0C0A4A480B0",
  2284 => x"C0C0C0C0A4A48099",
  2285 => x"C0C0C0C0A4A48092",
  2286 => x"C0C0C0C0A4A48082",
  2287 => x"C0C0C0C0A4A480F8",
  2288 => x"C0C0C0C0A4A48080",
  2289 => x"C0C0C0C0A4A48090",
  2290 => x"C0C0C0C0A4A490C0",
  2291 => x"C0C0C0C0A4A490F9",
  2292 => x"C0C0C0C0A4A490A4",
  2293 => x"C0C0C0C0A4A490B0",
  2294 => x"C0C0C0C0A4A49099",
  2295 => x"C0C0C0C0A4A49092",
  2296 => x"C0C0C0C0A4A49082",
  2297 => x"C0C0C0C0A4A490F8",
  2298 => x"C0C0C0C0A4A49080",
  2299 => x"C0C0C0C0A4A49090",
  2300 => x"C0C0C0C0A4B0C0C0",
  2301 => x"C0C0C0C0A4B0C0F9",
  2302 => x"C0C0C0C0A4B0C0A4",
  2303 => x"C0C0C0C0A4B0C0B0",
  2304 => x"C0C0C0C0A4B0C099",
  2305 => x"C0C0C0C0A4B0C092",
  2306 => x"C0C0C0C0A4B0C082",
  2307 => x"C0C0C0C0A4B0C0F8",
  2308 => x"C0C0C0C0A4B0C080",
  2309 => x"C0C0C0C0A4B0C090",
  2310 => x"C0C0C0C0A4B0F9C0",
  2311 => x"C0C0C0C0A4B0F9F9",
  2312 => x"C0C0C0C0A4B0F9A4",
  2313 => x"C0C0C0C0A4B0F9B0",
  2314 => x"C0C0C0C0A4B0F999",
  2315 => x"C0C0C0C0A4B0F992",
  2316 => x"C0C0C0C0A4B0F982",
  2317 => x"C0C0C0C0A4B0F9F8",
  2318 => x"C0C0C0C0A4B0F980",
  2319 => x"C0C0C0C0A4B0F990",
  2320 => x"C0C0C0C0A4B0A4C0",
  2321 => x"C0C0C0C0A4B0A4F9",
  2322 => x"C0C0C0C0A4B0A4A4",
  2323 => x"C0C0C0C0A4B0A4B0",
  2324 => x"C0C0C0C0A4B0A499",
  2325 => x"C0C0C0C0A4B0A492",
  2326 => x"C0C0C0C0A4B0A482",
  2327 => x"C0C0C0C0A4B0A4F8",
  2328 => x"C0C0C0C0A4B0A480",
  2329 => x"C0C0C0C0A4B0A490",
  2330 => x"C0C0C0C0A4B0B0C0",
  2331 => x"C0C0C0C0A4B0B0F9",
  2332 => x"C0C0C0C0A4B0B0A4",
  2333 => x"C0C0C0C0A4B0B0B0",
  2334 => x"C0C0C0C0A4B0B099",
  2335 => x"C0C0C0C0A4B0B092",
  2336 => x"C0C0C0C0A4B0B082",
  2337 => x"C0C0C0C0A4B0B0F8",
  2338 => x"C0C0C0C0A4B0B080",
  2339 => x"C0C0C0C0A4B0B090",
  2340 => x"C0C0C0C0A4B099C0",
  2341 => x"C0C0C0C0A4B099F9",
  2342 => x"C0C0C0C0A4B099A4",
  2343 => x"C0C0C0C0A4B099B0",
  2344 => x"C0C0C0C0A4B09999",
  2345 => x"C0C0C0C0A4B09992",
  2346 => x"C0C0C0C0A4B09982",
  2347 => x"C0C0C0C0A4B099F8",
  2348 => x"C0C0C0C0A4B09980",
  2349 => x"C0C0C0C0A4B09990",
  2350 => x"C0C0C0C0A4B092C0",
  2351 => x"C0C0C0C0A4B092F9",
  2352 => x"C0C0C0C0A4B092A4",
  2353 => x"C0C0C0C0A4B092B0",
  2354 => x"C0C0C0C0A4B09299",
  2355 => x"C0C0C0C0A4B09292",
  2356 => x"C0C0C0C0A4B09282",
  2357 => x"C0C0C0C0A4B092F8",
  2358 => x"C0C0C0C0A4B09280",
  2359 => x"C0C0C0C0A4B09290",
  2360 => x"C0C0C0C0A4B082C0",
  2361 => x"C0C0C0C0A4B082F9",
  2362 => x"C0C0C0C0A4B082A4",
  2363 => x"C0C0C0C0A4B082B0",
  2364 => x"C0C0C0C0A4B08299",
  2365 => x"C0C0C0C0A4B08292",
  2366 => x"C0C0C0C0A4B08282",
  2367 => x"C0C0C0C0A4B082F8",
  2368 => x"C0C0C0C0A4B08280",
  2369 => x"C0C0C0C0A4B08290",
  2370 => x"C0C0C0C0A4B0F8C0",
  2371 => x"C0C0C0C0A4B0F8F9",
  2372 => x"C0C0C0C0A4B0F8A4",
  2373 => x"C0C0C0C0A4B0F8B0",
  2374 => x"C0C0C0C0A4B0F899",
  2375 => x"C0C0C0C0A4B0F892",
  2376 => x"C0C0C0C0A4B0F882",
  2377 => x"C0C0C0C0A4B0F8F8",
  2378 => x"C0C0C0C0A4B0F880",
  2379 => x"C0C0C0C0A4B0F890",
  2380 => x"C0C0C0C0A4B080C0",
  2381 => x"C0C0C0C0A4B080F9",
  2382 => x"C0C0C0C0A4B080A4",
  2383 => x"C0C0C0C0A4B080B0",
  2384 => x"C0C0C0C0A4B08099",
  2385 => x"C0C0C0C0A4B08092",
  2386 => x"C0C0C0C0A4B08082",
  2387 => x"C0C0C0C0A4B080F8",
  2388 => x"C0C0C0C0A4B08080",
  2389 => x"C0C0C0C0A4B08090",
  2390 => x"C0C0C0C0A4B090C0",
  2391 => x"C0C0C0C0A4B090F9",
  2392 => x"C0C0C0C0A4B090A4",
  2393 => x"C0C0C0C0A4B090B0",
  2394 => x"C0C0C0C0A4B09099",
  2395 => x"C0C0C0C0A4B09092",
  2396 => x"C0C0C0C0A4B09082",
  2397 => x"C0C0C0C0A4B090F8",
  2398 => x"C0C0C0C0A4B09080",
  2399 => x"C0C0C0C0A4B09090",
  2400 => x"C0C0C0C0A499C0C0",
  2401 => x"C0C0C0C0A499C0F9",
  2402 => x"C0C0C0C0A499C0A4",
  2403 => x"C0C0C0C0A499C0B0",
  2404 => x"C0C0C0C0A499C099",
  2405 => x"C0C0C0C0A499C092",
  2406 => x"C0C0C0C0A499C082",
  2407 => x"C0C0C0C0A499C0F8",
  2408 => x"C0C0C0C0A499C080",
  2409 => x"C0C0C0C0A499C090",
  2410 => x"C0C0C0C0A499F9C0",
  2411 => x"C0C0C0C0A499F9F9",
  2412 => x"C0C0C0C0A499F9A4",
  2413 => x"C0C0C0C0A499F9B0",
  2414 => x"C0C0C0C0A499F999",
  2415 => x"C0C0C0C0A499F992",
  2416 => x"C0C0C0C0A499F982",
  2417 => x"C0C0C0C0A499F9F8",
  2418 => x"C0C0C0C0A499F980",
  2419 => x"C0C0C0C0A499F990",
  2420 => x"C0C0C0C0A499A4C0",
  2421 => x"C0C0C0C0A499A4F9",
  2422 => x"C0C0C0C0A499A4A4",
  2423 => x"C0C0C0C0A499A4B0",
  2424 => x"C0C0C0C0A499A499",
  2425 => x"C0C0C0C0A499A492",
  2426 => x"C0C0C0C0A499A482",
  2427 => x"C0C0C0C0A499A4F8",
  2428 => x"C0C0C0C0A499A480",
  2429 => x"C0C0C0C0A499A490",
  2430 => x"C0C0C0C0A499B0C0",
  2431 => x"C0C0C0C0A499B0F9",
  2432 => x"C0C0C0C0A499B0A4",
  2433 => x"C0C0C0C0A499B0B0",
  2434 => x"C0C0C0C0A499B099",
  2435 => x"C0C0C0C0A499B092",
  2436 => x"C0C0C0C0A499B082",
  2437 => x"C0C0C0C0A499B0F8",
  2438 => x"C0C0C0C0A499B080",
  2439 => x"C0C0C0C0A499B090",
  2440 => x"C0C0C0C0A49999C0",
  2441 => x"C0C0C0C0A49999F9",
  2442 => x"C0C0C0C0A49999A4",
  2443 => x"C0C0C0C0A49999B0",
  2444 => x"C0C0C0C0A4999999",
  2445 => x"C0C0C0C0A4999992",
  2446 => x"C0C0C0C0A4999982",
  2447 => x"C0C0C0C0A49999F8",
  2448 => x"C0C0C0C0A4999980",
  2449 => x"C0C0C0C0A4999990",
  2450 => x"C0C0C0C0A49992C0",
  2451 => x"C0C0C0C0A49992F9",
  2452 => x"C0C0C0C0A49992A4",
  2453 => x"C0C0C0C0A49992B0",
  2454 => x"C0C0C0C0A4999299",
  2455 => x"C0C0C0C0A4999292",
  2456 => x"C0C0C0C0A4999282",
  2457 => x"C0C0C0C0A49992F8",
  2458 => x"C0C0C0C0A4999280",
  2459 => x"C0C0C0C0A4999290",
  2460 => x"C0C0C0C0A49982C0",
  2461 => x"C0C0C0C0A49982F9",
  2462 => x"C0C0C0C0A49982A4",
  2463 => x"C0C0C0C0A49982B0",
  2464 => x"C0C0C0C0A4998299",
  2465 => x"C0C0C0C0A4998292",
  2466 => x"C0C0C0C0A4998282",
  2467 => x"C0C0C0C0A49982F8",
  2468 => x"C0C0C0C0A4998280",
  2469 => x"C0C0C0C0A4998290",
  2470 => x"C0C0C0C0A499F8C0",
  2471 => x"C0C0C0C0A499F8F9",
  2472 => x"C0C0C0C0A499F8A4",
  2473 => x"C0C0C0C0A499F8B0",
  2474 => x"C0C0C0C0A499F899",
  2475 => x"C0C0C0C0A499F892",
  2476 => x"C0C0C0C0A499F882",
  2477 => x"C0C0C0C0A499F8F8",
  2478 => x"C0C0C0C0A499F880",
  2479 => x"C0C0C0C0A499F890",
  2480 => x"C0C0C0C0A49980C0",
  2481 => x"C0C0C0C0A49980F9",
  2482 => x"C0C0C0C0A49980A4",
  2483 => x"C0C0C0C0A49980B0",
  2484 => x"C0C0C0C0A4998099",
  2485 => x"C0C0C0C0A4998092",
  2486 => x"C0C0C0C0A4998082",
  2487 => x"C0C0C0C0A49980F8",
  2488 => x"C0C0C0C0A4998080",
  2489 => x"C0C0C0C0A4998090",
  2490 => x"C0C0C0C0A49990C0",
  2491 => x"C0C0C0C0A49990F9",
  2492 => x"C0C0C0C0A49990A4",
  2493 => x"C0C0C0C0A49990B0",
  2494 => x"C0C0C0C0A4999099",
  2495 => x"C0C0C0C0A4999092",
  2496 => x"C0C0C0C0A4999082",
  2497 => x"C0C0C0C0A49990F8",
  2498 => x"C0C0C0C0A4999080",
  2499 => x"C0C0C0C0A4999090",
  2500 => x"C0C0C0C0A492C0C0",
  2501 => x"C0C0C0C0A492C0F9",
  2502 => x"C0C0C0C0A492C0A4",
  2503 => x"C0C0C0C0A492C0B0",
  2504 => x"C0C0C0C0A492C099",
  2505 => x"C0C0C0C0A492C092",
  2506 => x"C0C0C0C0A492C082",
  2507 => x"C0C0C0C0A492C0F8",
  2508 => x"C0C0C0C0A492C080",
  2509 => x"C0C0C0C0A492C090",
  2510 => x"C0C0C0C0A492F9C0",
  2511 => x"C0C0C0C0A492F9F9",
  2512 => x"C0C0C0C0A492F9A4",
  2513 => x"C0C0C0C0A492F9B0",
  2514 => x"C0C0C0C0A492F999",
  2515 => x"C0C0C0C0A492F992",
  2516 => x"C0C0C0C0A492F982",
  2517 => x"C0C0C0C0A492F9F8",
  2518 => x"C0C0C0C0A492F980",
  2519 => x"C0C0C0C0A492F990",
  2520 => x"C0C0C0C0A492A4C0",
  2521 => x"C0C0C0C0A492A4F9",
  2522 => x"C0C0C0C0A492A4A4",
  2523 => x"C0C0C0C0A492A4B0",
  2524 => x"C0C0C0C0A492A499",
  2525 => x"C0C0C0C0A492A492",
  2526 => x"C0C0C0C0A492A482",
  2527 => x"C0C0C0C0A492A4F8",
  2528 => x"C0C0C0C0A492A480",
  2529 => x"C0C0C0C0A492A490",
  2530 => x"C0C0C0C0A492B0C0",
  2531 => x"C0C0C0C0A492B0F9",
  2532 => x"C0C0C0C0A492B0A4",
  2533 => x"C0C0C0C0A492B0B0",
  2534 => x"C0C0C0C0A492B099",
  2535 => x"C0C0C0C0A492B092",
  2536 => x"C0C0C0C0A492B082",
  2537 => x"C0C0C0C0A492B0F8",
  2538 => x"C0C0C0C0A492B080",
  2539 => x"C0C0C0C0A492B090",
  2540 => x"C0C0C0C0A49299C0",
  2541 => x"C0C0C0C0A49299F9",
  2542 => x"C0C0C0C0A49299A4",
  2543 => x"C0C0C0C0A49299B0",
  2544 => x"C0C0C0C0A4929999",
  2545 => x"C0C0C0C0A4929992",
  2546 => x"C0C0C0C0A4929982",
  2547 => x"C0C0C0C0A49299F8",
  2548 => x"C0C0C0C0A4929980",
  2549 => x"C0C0C0C0A4929990",
  2550 => x"C0C0C0C0A49292C0",
  2551 => x"C0C0C0C0A49292F9",
  2552 => x"C0C0C0C0A49292A4",
  2553 => x"C0C0C0C0A49292B0",
  2554 => x"C0C0C0C0A4929299",
  2555 => x"C0C0C0C0A4929292",
  2556 => x"C0C0C0C0A4929282",
  2557 => x"C0C0C0C0A49292F8",
  2558 => x"C0C0C0C0A4929280",
  2559 => x"C0C0C0C0A4929290",
  2560 => x"C0C0C0C0A49282C0",
  2561 => x"C0C0C0C0A49282F9",
  2562 => x"C0C0C0C0A49282A4",
  2563 => x"C0C0C0C0A49282B0",
  2564 => x"C0C0C0C0A4928299",
  2565 => x"C0C0C0C0A4928292",
  2566 => x"C0C0C0C0A4928282",
  2567 => x"C0C0C0C0A49282F8",
  2568 => x"C0C0C0C0A4928280",
  2569 => x"C0C0C0C0A4928290",
  2570 => x"C0C0C0C0A492F8C0",
  2571 => x"C0C0C0C0A492F8F9",
  2572 => x"C0C0C0C0A492F8A4",
  2573 => x"C0C0C0C0A492F8B0",
  2574 => x"C0C0C0C0A492F899",
  2575 => x"C0C0C0C0A492F892",
  2576 => x"C0C0C0C0A492F882",
  2577 => x"C0C0C0C0A492F8F8",
  2578 => x"C0C0C0C0A492F880",
  2579 => x"C0C0C0C0A492F890",
  2580 => x"C0C0C0C0A49280C0",
  2581 => x"C0C0C0C0A49280F9",
  2582 => x"C0C0C0C0A49280A4",
  2583 => x"C0C0C0C0A49280B0",
  2584 => x"C0C0C0C0A4928099",
  2585 => x"C0C0C0C0A4928092",
  2586 => x"C0C0C0C0A4928082",
  2587 => x"C0C0C0C0A49280F8",
  2588 => x"C0C0C0C0A4928080",
  2589 => x"C0C0C0C0A4928090",
  2590 => x"C0C0C0C0A49290C0",
  2591 => x"C0C0C0C0A49290F9",
  2592 => x"C0C0C0C0A49290A4",
  2593 => x"C0C0C0C0A49290B0",
  2594 => x"C0C0C0C0A4929099",
  2595 => x"C0C0C0C0A4929092",
  2596 => x"C0C0C0C0A4929082",
  2597 => x"C0C0C0C0A49290F8",
  2598 => x"C0C0C0C0A4929080",
  2599 => x"C0C0C0C0A4929090",
  2600 => x"C0C0C0C0A482C0C0",
  2601 => x"C0C0C0C0A482C0F9",
  2602 => x"C0C0C0C0A482C0A4",
  2603 => x"C0C0C0C0A482C0B0",
  2604 => x"C0C0C0C0A482C099",
  2605 => x"C0C0C0C0A482C092",
  2606 => x"C0C0C0C0A482C082",
  2607 => x"C0C0C0C0A482C0F8",
  2608 => x"C0C0C0C0A482C080",
  2609 => x"C0C0C0C0A482C090",
  2610 => x"C0C0C0C0A482F9C0",
  2611 => x"C0C0C0C0A482F9F9",
  2612 => x"C0C0C0C0A482F9A4",
  2613 => x"C0C0C0C0A482F9B0",
  2614 => x"C0C0C0C0A482F999",
  2615 => x"C0C0C0C0A482F992",
  2616 => x"C0C0C0C0A482F982",
  2617 => x"C0C0C0C0A482F9F8",
  2618 => x"C0C0C0C0A482F980",
  2619 => x"C0C0C0C0A482F990",
  2620 => x"C0C0C0C0A482A4C0",
  2621 => x"C0C0C0C0A482A4F9",
  2622 => x"C0C0C0C0A482A4A4",
  2623 => x"C0C0C0C0A482A4B0",
  2624 => x"C0C0C0C0A482A499",
  2625 => x"C0C0C0C0A482A492",
  2626 => x"C0C0C0C0A482A482",
  2627 => x"C0C0C0C0A482A4F8",
  2628 => x"C0C0C0C0A482A480",
  2629 => x"C0C0C0C0A482A490",
  2630 => x"C0C0C0C0A482B0C0",
  2631 => x"C0C0C0C0A482B0F9",
  2632 => x"C0C0C0C0A482B0A4",
  2633 => x"C0C0C0C0A482B0B0",
  2634 => x"C0C0C0C0A482B099",
  2635 => x"C0C0C0C0A482B092",
  2636 => x"C0C0C0C0A482B082",
  2637 => x"C0C0C0C0A482B0F8",
  2638 => x"C0C0C0C0A482B080",
  2639 => x"C0C0C0C0A482B090",
  2640 => x"C0C0C0C0A48299C0",
  2641 => x"C0C0C0C0A48299F9",
  2642 => x"C0C0C0C0A48299A4",
  2643 => x"C0C0C0C0A48299B0",
  2644 => x"C0C0C0C0A4829999",
  2645 => x"C0C0C0C0A4829992",
  2646 => x"C0C0C0C0A4829982",
  2647 => x"C0C0C0C0A48299F8",
  2648 => x"C0C0C0C0A4829980",
  2649 => x"C0C0C0C0A4829990",
  2650 => x"C0C0C0C0A48292C0",
  2651 => x"C0C0C0C0A48292F9",
  2652 => x"C0C0C0C0A48292A4",
  2653 => x"C0C0C0C0A48292B0",
  2654 => x"C0C0C0C0A4829299",
  2655 => x"C0C0C0C0A4829292",
  2656 => x"C0C0C0C0A4829282",
  2657 => x"C0C0C0C0A48292F8",
  2658 => x"C0C0C0C0A4829280",
  2659 => x"C0C0C0C0A4829290",
  2660 => x"C0C0C0C0A48282C0",
  2661 => x"C0C0C0C0A48282F9",
  2662 => x"C0C0C0C0A48282A4",
  2663 => x"C0C0C0C0A48282B0",
  2664 => x"C0C0C0C0A4828299",
  2665 => x"C0C0C0C0A4828292",
  2666 => x"C0C0C0C0A4828282",
  2667 => x"C0C0C0C0A48282F8",
  2668 => x"C0C0C0C0A4828280",
  2669 => x"C0C0C0C0A4828290",
  2670 => x"C0C0C0C0A482F8C0",
  2671 => x"C0C0C0C0A482F8F9",
  2672 => x"C0C0C0C0A482F8A4",
  2673 => x"C0C0C0C0A482F8B0",
  2674 => x"C0C0C0C0A482F899",
  2675 => x"C0C0C0C0A482F892",
  2676 => x"C0C0C0C0A482F882",
  2677 => x"C0C0C0C0A482F8F8",
  2678 => x"C0C0C0C0A482F880",
  2679 => x"C0C0C0C0A482F890",
  2680 => x"C0C0C0C0A48280C0",
  2681 => x"C0C0C0C0A48280F9",
  2682 => x"C0C0C0C0A48280A4",
  2683 => x"C0C0C0C0A48280B0",
  2684 => x"C0C0C0C0A4828099",
  2685 => x"C0C0C0C0A4828092",
  2686 => x"C0C0C0C0A4828082",
  2687 => x"C0C0C0C0A48280F8",
  2688 => x"C0C0C0C0A4828080",
  2689 => x"C0C0C0C0A4828090",
  2690 => x"C0C0C0C0A48290C0",
  2691 => x"C0C0C0C0A48290F9",
  2692 => x"C0C0C0C0A48290A4",
  2693 => x"C0C0C0C0A48290B0",
  2694 => x"C0C0C0C0A4829099",
  2695 => x"C0C0C0C0A4829092",
  2696 => x"C0C0C0C0A4829082",
  2697 => x"C0C0C0C0A48290F8",
  2698 => x"C0C0C0C0A4829080",
  2699 => x"C0C0C0C0A4829090",
  2700 => x"C0C0C0C0A4F8C0C0",
  2701 => x"C0C0C0C0A4F8C0F9",
  2702 => x"C0C0C0C0A4F8C0A4",
  2703 => x"C0C0C0C0A4F8C0B0",
  2704 => x"C0C0C0C0A4F8C099",
  2705 => x"C0C0C0C0A4F8C092",
  2706 => x"C0C0C0C0A4F8C082",
  2707 => x"C0C0C0C0A4F8C0F8",
  2708 => x"C0C0C0C0A4F8C080",
  2709 => x"C0C0C0C0A4F8C090",
  2710 => x"C0C0C0C0A4F8F9C0",
  2711 => x"C0C0C0C0A4F8F9F9",
  2712 => x"C0C0C0C0A4F8F9A4",
  2713 => x"C0C0C0C0A4F8F9B0",
  2714 => x"C0C0C0C0A4F8F999",
  2715 => x"C0C0C0C0A4F8F992",
  2716 => x"C0C0C0C0A4F8F982",
  2717 => x"C0C0C0C0A4F8F9F8",
  2718 => x"C0C0C0C0A4F8F980",
  2719 => x"C0C0C0C0A4F8F990",
  2720 => x"C0C0C0C0A4F8A4C0",
  2721 => x"C0C0C0C0A4F8A4F9",
  2722 => x"C0C0C0C0A4F8A4A4",
  2723 => x"C0C0C0C0A4F8A4B0",
  2724 => x"C0C0C0C0A4F8A499",
  2725 => x"C0C0C0C0A4F8A492",
  2726 => x"C0C0C0C0A4F8A482",
  2727 => x"C0C0C0C0A4F8A4F8",
  2728 => x"C0C0C0C0A4F8A480",
  2729 => x"C0C0C0C0A4F8A490",
  2730 => x"C0C0C0C0A4F8B0C0",
  2731 => x"C0C0C0C0A4F8B0F9",
  2732 => x"C0C0C0C0A4F8B0A4",
  2733 => x"C0C0C0C0A4F8B0B0",
  2734 => x"C0C0C0C0A4F8B099",
  2735 => x"C0C0C0C0A4F8B092",
  2736 => x"C0C0C0C0A4F8B082",
  2737 => x"C0C0C0C0A4F8B0F8",
  2738 => x"C0C0C0C0A4F8B080",
  2739 => x"C0C0C0C0A4F8B090",
  2740 => x"C0C0C0C0A4F899C0",
  2741 => x"C0C0C0C0A4F899F9",
  2742 => x"C0C0C0C0A4F899A4",
  2743 => x"C0C0C0C0A4F899B0",
  2744 => x"C0C0C0C0A4F89999",
  2745 => x"C0C0C0C0A4F89992",
  2746 => x"C0C0C0C0A4F89982",
  2747 => x"C0C0C0C0A4F899F8",
  2748 => x"C0C0C0C0A4F89980",
  2749 => x"C0C0C0C0A4F89990",
  2750 => x"C0C0C0C0A4F892C0",
  2751 => x"C0C0C0C0A4F892F9",
  2752 => x"C0C0C0C0A4F892A4",
  2753 => x"C0C0C0C0A4F892B0",
  2754 => x"C0C0C0C0A4F89299",
  2755 => x"C0C0C0C0A4F89292",
  2756 => x"C0C0C0C0A4F89282",
  2757 => x"C0C0C0C0A4F892F8",
  2758 => x"C0C0C0C0A4F89280",
  2759 => x"C0C0C0C0A4F89290",
  2760 => x"C0C0C0C0A4F882C0",
  2761 => x"C0C0C0C0A4F882F9",
  2762 => x"C0C0C0C0A4F882A4",
  2763 => x"C0C0C0C0A4F882B0",
  2764 => x"C0C0C0C0A4F88299",
  2765 => x"C0C0C0C0A4F88292",
  2766 => x"C0C0C0C0A4F88282",
  2767 => x"C0C0C0C0A4F882F8",
  2768 => x"C0C0C0C0A4F88280",
  2769 => x"C0C0C0C0A4F88290",
  2770 => x"C0C0C0C0A4F8F8C0",
  2771 => x"C0C0C0C0A4F8F8F9",
  2772 => x"C0C0C0C0A4F8F8A4",
  2773 => x"C0C0C0C0A4F8F8B0",
  2774 => x"C0C0C0C0A4F8F899",
  2775 => x"C0C0C0C0A4F8F892",
  2776 => x"C0C0C0C0A4F8F882",
  2777 => x"C0C0C0C0A4F8F8F8",
  2778 => x"C0C0C0C0A4F8F880",
  2779 => x"C0C0C0C0A4F8F890",
  2780 => x"C0C0C0C0A4F880C0",
  2781 => x"C0C0C0C0A4F880F9",
  2782 => x"C0C0C0C0A4F880A4",
  2783 => x"C0C0C0C0A4F880B0",
  2784 => x"C0C0C0C0A4F88099",
  2785 => x"C0C0C0C0A4F88092",
  2786 => x"C0C0C0C0A4F88082",
  2787 => x"C0C0C0C0A4F880F8",
  2788 => x"C0C0C0C0A4F88080",
  2789 => x"C0C0C0C0A4F88090",
  2790 => x"C0C0C0C0A4F890C0",
  2791 => x"C0C0C0C0A4F890F9",
  2792 => x"C0C0C0C0A4F890A4",
  2793 => x"C0C0C0C0A4F890B0",
  2794 => x"C0C0C0C0A4F89099",
  2795 => x"C0C0C0C0A4F89092",
  2796 => x"C0C0C0C0A4F89082",
  2797 => x"C0C0C0C0A4F890F8",
  2798 => x"C0C0C0C0A4F89080",
  2799 => x"C0C0C0C0A4F89090",
  2800 => x"C0C0C0C0A480C0C0",
  2801 => x"C0C0C0C0A480C0F9",
  2802 => x"C0C0C0C0A480C0A4",
  2803 => x"C0C0C0C0A480C0B0",
  2804 => x"C0C0C0C0A480C099",
  2805 => x"C0C0C0C0A480C092",
  2806 => x"C0C0C0C0A480C082",
  2807 => x"C0C0C0C0A480C0F8",
  2808 => x"C0C0C0C0A480C080",
  2809 => x"C0C0C0C0A480C090",
  2810 => x"C0C0C0C0A480F9C0",
  2811 => x"C0C0C0C0A480F9F9",
  2812 => x"C0C0C0C0A480F9A4",
  2813 => x"C0C0C0C0A480F9B0",
  2814 => x"C0C0C0C0A480F999",
  2815 => x"C0C0C0C0A480F992",
  2816 => x"C0C0C0C0A480F982",
  2817 => x"C0C0C0C0A480F9F8",
  2818 => x"C0C0C0C0A480F980",
  2819 => x"C0C0C0C0A480F990",
  2820 => x"C0C0C0C0A480A4C0",
  2821 => x"C0C0C0C0A480A4F9",
  2822 => x"C0C0C0C0A480A4A4",
  2823 => x"C0C0C0C0A480A4B0",
  2824 => x"C0C0C0C0A480A499",
  2825 => x"C0C0C0C0A480A492",
  2826 => x"C0C0C0C0A480A482",
  2827 => x"C0C0C0C0A480A4F8",
  2828 => x"C0C0C0C0A480A480",
  2829 => x"C0C0C0C0A480A490",
  2830 => x"C0C0C0C0A480B0C0",
  2831 => x"C0C0C0C0A480B0F9",
  2832 => x"C0C0C0C0A480B0A4",
  2833 => x"C0C0C0C0A480B0B0",
  2834 => x"C0C0C0C0A480B099",
  2835 => x"C0C0C0C0A480B092",
  2836 => x"C0C0C0C0A480B082",
  2837 => x"C0C0C0C0A480B0F8",
  2838 => x"C0C0C0C0A480B080",
  2839 => x"C0C0C0C0A480B090",
  2840 => x"C0C0C0C0A48099C0",
  2841 => x"C0C0C0C0A48099F9",
  2842 => x"C0C0C0C0A48099A4",
  2843 => x"C0C0C0C0A48099B0",
  2844 => x"C0C0C0C0A4809999",
  2845 => x"C0C0C0C0A4809992",
  2846 => x"C0C0C0C0A4809982",
  2847 => x"C0C0C0C0A48099F8",
  2848 => x"C0C0C0C0A4809980",
  2849 => x"C0C0C0C0A4809990",
  2850 => x"C0C0C0C0A48092C0",
  2851 => x"C0C0C0C0A48092F9",
  2852 => x"C0C0C0C0A48092A4",
  2853 => x"C0C0C0C0A48092B0",
  2854 => x"C0C0C0C0A4809299",
  2855 => x"C0C0C0C0A4809292",
  2856 => x"C0C0C0C0A4809282",
  2857 => x"C0C0C0C0A48092F8",
  2858 => x"C0C0C0C0A4809280",
  2859 => x"C0C0C0C0A4809290",
  2860 => x"C0C0C0C0A48082C0",
  2861 => x"C0C0C0C0A48082F9",
  2862 => x"C0C0C0C0A48082A4",
  2863 => x"C0C0C0C0A48082B0",
  2864 => x"C0C0C0C0A4808299",
  2865 => x"C0C0C0C0A4808292",
  2866 => x"C0C0C0C0A4808282",
  2867 => x"C0C0C0C0A48082F8",
  2868 => x"C0C0C0C0A4808280",
  2869 => x"C0C0C0C0A4808290",
  2870 => x"C0C0C0C0A480F8C0",
  2871 => x"C0C0C0C0A480F8F9",
  2872 => x"C0C0C0C0A480F8A4",
  2873 => x"C0C0C0C0A480F8B0",
  2874 => x"C0C0C0C0A480F899",
  2875 => x"C0C0C0C0A480F892",
  2876 => x"C0C0C0C0A480F882",
  2877 => x"C0C0C0C0A480F8F8",
  2878 => x"C0C0C0C0A480F880",
  2879 => x"C0C0C0C0A480F890",
  2880 => x"C0C0C0C0A48080C0",
  2881 => x"C0C0C0C0A48080F9",
  2882 => x"C0C0C0C0A48080A4",
  2883 => x"C0C0C0C0A48080B0",
  2884 => x"C0C0C0C0A4808099",
  2885 => x"C0C0C0C0A4808092",
  2886 => x"C0C0C0C0A4808082",
  2887 => x"C0C0C0C0A48080F8",
  2888 => x"C0C0C0C0A4808080",
  2889 => x"C0C0C0C0A4808090",
  2890 => x"C0C0C0C0A48090C0",
  2891 => x"C0C0C0C0A48090F9",
  2892 => x"C0C0C0C0A48090A4",
  2893 => x"C0C0C0C0A48090B0",
  2894 => x"C0C0C0C0A4809099",
  2895 => x"C0C0C0C0A4809092",
  2896 => x"C0C0C0C0A4809082",
  2897 => x"C0C0C0C0A48090F8",
  2898 => x"C0C0C0C0A4809080",
  2899 => x"C0C0C0C0A4809090",
  2900 => x"C0C0C0C0A490C0C0",
  2901 => x"C0C0C0C0A490C0F9",
  2902 => x"C0C0C0C0A490C0A4",
  2903 => x"C0C0C0C0A490C0B0",
  2904 => x"C0C0C0C0A490C099",
  2905 => x"C0C0C0C0A490C092",
  2906 => x"C0C0C0C0A490C082",
  2907 => x"C0C0C0C0A490C0F8",
  2908 => x"C0C0C0C0A490C080",
  2909 => x"C0C0C0C0A490C090",
  2910 => x"C0C0C0C0A490F9C0",
  2911 => x"C0C0C0C0A490F9F9",
  2912 => x"C0C0C0C0A490F9A4",
  2913 => x"C0C0C0C0A490F9B0",
  2914 => x"C0C0C0C0A490F999",
  2915 => x"C0C0C0C0A490F992",
  2916 => x"C0C0C0C0A490F982",
  2917 => x"C0C0C0C0A490F9F8",
  2918 => x"C0C0C0C0A490F980",
  2919 => x"C0C0C0C0A490F990",
  2920 => x"C0C0C0C0A490A4C0",
  2921 => x"C0C0C0C0A490A4F9",
  2922 => x"C0C0C0C0A490A4A4",
  2923 => x"C0C0C0C0A490A4B0",
  2924 => x"C0C0C0C0A490A499",
  2925 => x"C0C0C0C0A490A492",
  2926 => x"C0C0C0C0A490A482",
  2927 => x"C0C0C0C0A490A4F8",
  2928 => x"C0C0C0C0A490A480",
  2929 => x"C0C0C0C0A490A490",
  2930 => x"C0C0C0C0A490B0C0",
  2931 => x"C0C0C0C0A490B0F9",
  2932 => x"C0C0C0C0A490B0A4",
  2933 => x"C0C0C0C0A490B0B0",
  2934 => x"C0C0C0C0A490B099",
  2935 => x"C0C0C0C0A490B092",
  2936 => x"C0C0C0C0A490B082",
  2937 => x"C0C0C0C0A490B0F8",
  2938 => x"C0C0C0C0A490B080",
  2939 => x"C0C0C0C0A490B090",
  2940 => x"C0C0C0C0A49099C0",
  2941 => x"C0C0C0C0A49099F9",
  2942 => x"C0C0C0C0A49099A4",
  2943 => x"C0C0C0C0A49099B0",
  2944 => x"C0C0C0C0A4909999",
  2945 => x"C0C0C0C0A4909992",
  2946 => x"C0C0C0C0A4909982",
  2947 => x"C0C0C0C0A49099F8",
  2948 => x"C0C0C0C0A4909980",
  2949 => x"C0C0C0C0A4909990",
  2950 => x"C0C0C0C0A49092C0",
  2951 => x"C0C0C0C0A49092F9",
  2952 => x"C0C0C0C0A49092A4",
  2953 => x"C0C0C0C0A49092B0",
  2954 => x"C0C0C0C0A4909299",
  2955 => x"C0C0C0C0A4909292",
  2956 => x"C0C0C0C0A4909282",
  2957 => x"C0C0C0C0A49092F8",
  2958 => x"C0C0C0C0A4909280",
  2959 => x"C0C0C0C0A4909290",
  2960 => x"C0C0C0C0A49082C0",
  2961 => x"C0C0C0C0A49082F9",
  2962 => x"C0C0C0C0A49082A4",
  2963 => x"C0C0C0C0A49082B0",
  2964 => x"C0C0C0C0A4908299",
  2965 => x"C0C0C0C0A4908292",
  2966 => x"C0C0C0C0A4908282",
  2967 => x"C0C0C0C0A49082F8",
  2968 => x"C0C0C0C0A4908280",
  2969 => x"C0C0C0C0A4908290",
  2970 => x"C0C0C0C0A490F8C0",
  2971 => x"C0C0C0C0A490F8F9",
  2972 => x"C0C0C0C0A490F8A4",
  2973 => x"C0C0C0C0A490F8B0",
  2974 => x"C0C0C0C0A490F899",
  2975 => x"C0C0C0C0A490F892",
  2976 => x"C0C0C0C0A490F882",
  2977 => x"C0C0C0C0A490F8F8",
  2978 => x"C0C0C0C0A490F880",
  2979 => x"C0C0C0C0A490F890",
  2980 => x"C0C0C0C0A49080C0",
  2981 => x"C0C0C0C0A49080F9",
  2982 => x"C0C0C0C0A49080A4",
  2983 => x"C0C0C0C0A49080B0",
  2984 => x"C0C0C0C0A4908099",
  2985 => x"C0C0C0C0A4908092",
  2986 => x"C0C0C0C0A4908082",
  2987 => x"C0C0C0C0A49080F8",
  2988 => x"C0C0C0C0A4908080",
  2989 => x"C0C0C0C0A4908090",
  2990 => x"C0C0C0C0A49090C0",
  2991 => x"C0C0C0C0A49090F9",
  2992 => x"C0C0C0C0A49090A4",
  2993 => x"C0C0C0C0A49090B0",
  2994 => x"C0C0C0C0A4909099",
  2995 => x"C0C0C0C0A4909092",
  2996 => x"C0C0C0C0A4909082",
  2997 => x"C0C0C0C0A49090F8",
  2998 => x"C0C0C0C0A4909080",
  2999 => x"C0C0C0C0A4909090",
  3000 => x"C0C0C0C0B0C0C0C0",
  3001 => x"C0C0C0C0B0C0C0F9",
  3002 => x"C0C0C0C0B0C0C0A4",
  3003 => x"C0C0C0C0B0C0C0B0",
  3004 => x"C0C0C0C0B0C0C099",
  3005 => x"C0C0C0C0B0C0C092",
  3006 => x"C0C0C0C0B0C0C082",
  3007 => x"C0C0C0C0B0C0C0F8",
  3008 => x"C0C0C0C0B0C0C080",
  3009 => x"C0C0C0C0B0C0C090",
  3010 => x"C0C0C0C0B0C0F9C0",
  3011 => x"C0C0C0C0B0C0F9F9",
  3012 => x"C0C0C0C0B0C0F9A4",
  3013 => x"C0C0C0C0B0C0F9B0",
  3014 => x"C0C0C0C0B0C0F999",
  3015 => x"C0C0C0C0B0C0F992",
  3016 => x"C0C0C0C0B0C0F982",
  3017 => x"C0C0C0C0B0C0F9F8",
  3018 => x"C0C0C0C0B0C0F980",
  3019 => x"C0C0C0C0B0C0F990",
  3020 => x"C0C0C0C0B0C0A4C0",
  3021 => x"C0C0C0C0B0C0A4F9",
  3022 => x"C0C0C0C0B0C0A4A4",
  3023 => x"C0C0C0C0B0C0A4B0",
  3024 => x"C0C0C0C0B0C0A499",
  3025 => x"C0C0C0C0B0C0A492",
  3026 => x"C0C0C0C0B0C0A482",
  3027 => x"C0C0C0C0B0C0A4F8",
  3028 => x"C0C0C0C0B0C0A480",
  3029 => x"C0C0C0C0B0C0A490",
  3030 => x"C0C0C0C0B0C0B0C0",
  3031 => x"C0C0C0C0B0C0B0F9",
  3032 => x"C0C0C0C0B0C0B0A4",
  3033 => x"C0C0C0C0B0C0B0B0",
  3034 => x"C0C0C0C0B0C0B099",
  3035 => x"C0C0C0C0B0C0B092",
  3036 => x"C0C0C0C0B0C0B082",
  3037 => x"C0C0C0C0B0C0B0F8",
  3038 => x"C0C0C0C0B0C0B080",
  3039 => x"C0C0C0C0B0C0B090",
  3040 => x"C0C0C0C0B0C099C0",
  3041 => x"C0C0C0C0B0C099F9",
  3042 => x"C0C0C0C0B0C099A4",
  3043 => x"C0C0C0C0B0C099B0",
  3044 => x"C0C0C0C0B0C09999",
  3045 => x"C0C0C0C0B0C09992",
  3046 => x"C0C0C0C0B0C09982",
  3047 => x"C0C0C0C0B0C099F8",
  3048 => x"C0C0C0C0B0C09980",
  3049 => x"C0C0C0C0B0C09990",
  3050 => x"C0C0C0C0B0C092C0",
  3051 => x"C0C0C0C0B0C092F9",
  3052 => x"C0C0C0C0B0C092A4",
  3053 => x"C0C0C0C0B0C092B0",
  3054 => x"C0C0C0C0B0C09299",
  3055 => x"C0C0C0C0B0C09292",
  3056 => x"C0C0C0C0B0C09282",
  3057 => x"C0C0C0C0B0C092F8",
  3058 => x"C0C0C0C0B0C09280",
  3059 => x"C0C0C0C0B0C09290",
  3060 => x"C0C0C0C0B0C082C0",
  3061 => x"C0C0C0C0B0C082F9",
  3062 => x"C0C0C0C0B0C082A4",
  3063 => x"C0C0C0C0B0C082B0",
  3064 => x"C0C0C0C0B0C08299",
  3065 => x"C0C0C0C0B0C08292",
  3066 => x"C0C0C0C0B0C08282",
  3067 => x"C0C0C0C0B0C082F8",
  3068 => x"C0C0C0C0B0C08280",
  3069 => x"C0C0C0C0B0C08290",
  3070 => x"C0C0C0C0B0C0F8C0",
  3071 => x"C0C0C0C0B0C0F8F9",
  3072 => x"C0C0C0C0B0C0F8A4",
  3073 => x"C0C0C0C0B0C0F8B0",
  3074 => x"C0C0C0C0B0C0F899",
  3075 => x"C0C0C0C0B0C0F892",
  3076 => x"C0C0C0C0B0C0F882",
  3077 => x"C0C0C0C0B0C0F8F8",
  3078 => x"C0C0C0C0B0C0F880",
  3079 => x"C0C0C0C0B0C0F890",
  3080 => x"C0C0C0C0B0C080C0",
  3081 => x"C0C0C0C0B0C080F9",
  3082 => x"C0C0C0C0B0C080A4",
  3083 => x"C0C0C0C0B0C080B0",
  3084 => x"C0C0C0C0B0C08099",
  3085 => x"C0C0C0C0B0C08092",
  3086 => x"C0C0C0C0B0C08082",
  3087 => x"C0C0C0C0B0C080F8",
  3088 => x"C0C0C0C0B0C08080",
  3089 => x"C0C0C0C0B0C08090",
  3090 => x"C0C0C0C0B0C090C0",
  3091 => x"C0C0C0C0B0C090F9",
  3092 => x"C0C0C0C0B0C090A4",
  3093 => x"C0C0C0C0B0C090B0",
  3094 => x"C0C0C0C0B0C09099",
  3095 => x"C0C0C0C0B0C09092",
  3096 => x"C0C0C0C0B0C09082",
  3097 => x"C0C0C0C0B0C090F8",
  3098 => x"C0C0C0C0B0C09080",
  3099 => x"C0C0C0C0B0C09090",
  3100 => x"C0C0C0C0B0F9C0C0",
  3101 => x"C0C0C0C0B0F9C0F9",
  3102 => x"C0C0C0C0B0F9C0A4",
  3103 => x"C0C0C0C0B0F9C0B0",
  3104 => x"C0C0C0C0B0F9C099",
  3105 => x"C0C0C0C0B0F9C092",
  3106 => x"C0C0C0C0B0F9C082",
  3107 => x"C0C0C0C0B0F9C0F8",
  3108 => x"C0C0C0C0B0F9C080",
  3109 => x"C0C0C0C0B0F9C090",
  3110 => x"C0C0C0C0B0F9F9C0",
  3111 => x"C0C0C0C0B0F9F9F9",
  3112 => x"C0C0C0C0B0F9F9A4",
  3113 => x"C0C0C0C0B0F9F9B0",
  3114 => x"C0C0C0C0B0F9F999",
  3115 => x"C0C0C0C0B0F9F992",
  3116 => x"C0C0C0C0B0F9F982",
  3117 => x"C0C0C0C0B0F9F9F8",
  3118 => x"C0C0C0C0B0F9F980",
  3119 => x"C0C0C0C0B0F9F990",
  3120 => x"C0C0C0C0B0F9A4C0",
  3121 => x"C0C0C0C0B0F9A4F9",
  3122 => x"C0C0C0C0B0F9A4A4",
  3123 => x"C0C0C0C0B0F9A4B0",
  3124 => x"C0C0C0C0B0F9A499",
  3125 => x"C0C0C0C0B0F9A492",
  3126 => x"C0C0C0C0B0F9A482",
  3127 => x"C0C0C0C0B0F9A4F8",
  3128 => x"C0C0C0C0B0F9A480",
  3129 => x"C0C0C0C0B0F9A490",
  3130 => x"C0C0C0C0B0F9B0C0",
  3131 => x"C0C0C0C0B0F9B0F9",
  3132 => x"C0C0C0C0B0F9B0A4",
  3133 => x"C0C0C0C0B0F9B0B0",
  3134 => x"C0C0C0C0B0F9B099",
  3135 => x"C0C0C0C0B0F9B092",
  3136 => x"C0C0C0C0B0F9B082",
  3137 => x"C0C0C0C0B0F9B0F8",
  3138 => x"C0C0C0C0B0F9B080",
  3139 => x"C0C0C0C0B0F9B090",
  3140 => x"C0C0C0C0B0F999C0",
  3141 => x"C0C0C0C0B0F999F9",
  3142 => x"C0C0C0C0B0F999A4",
  3143 => x"C0C0C0C0B0F999B0",
  3144 => x"C0C0C0C0B0F99999",
  3145 => x"C0C0C0C0B0F99992",
  3146 => x"C0C0C0C0B0F99982",
  3147 => x"C0C0C0C0B0F999F8",
  3148 => x"C0C0C0C0B0F99980",
  3149 => x"C0C0C0C0B0F99990",
  3150 => x"C0C0C0C0B0F992C0",
  3151 => x"C0C0C0C0B0F992F9",
  3152 => x"C0C0C0C0B0F992A4",
  3153 => x"C0C0C0C0B0F992B0",
  3154 => x"C0C0C0C0B0F99299",
  3155 => x"C0C0C0C0B0F99292",
  3156 => x"C0C0C0C0B0F99282",
  3157 => x"C0C0C0C0B0F992F8",
  3158 => x"C0C0C0C0B0F99280",
  3159 => x"C0C0C0C0B0F99290",
  3160 => x"C0C0C0C0B0F982C0",
  3161 => x"C0C0C0C0B0F982F9",
  3162 => x"C0C0C0C0B0F982A4",
  3163 => x"C0C0C0C0B0F982B0",
  3164 => x"C0C0C0C0B0F98299",
  3165 => x"C0C0C0C0B0F98292",
  3166 => x"C0C0C0C0B0F98282",
  3167 => x"C0C0C0C0B0F982F8",
  3168 => x"C0C0C0C0B0F98280",
  3169 => x"C0C0C0C0B0F98290",
  3170 => x"C0C0C0C0B0F9F8C0",
  3171 => x"C0C0C0C0B0F9F8F9",
  3172 => x"C0C0C0C0B0F9F8A4",
  3173 => x"C0C0C0C0B0F9F8B0",
  3174 => x"C0C0C0C0B0F9F899",
  3175 => x"C0C0C0C0B0F9F892",
  3176 => x"C0C0C0C0B0F9F882",
  3177 => x"C0C0C0C0B0F9F8F8",
  3178 => x"C0C0C0C0B0F9F880",
  3179 => x"C0C0C0C0B0F9F890",
  3180 => x"C0C0C0C0B0F980C0",
  3181 => x"C0C0C0C0B0F980F9",
  3182 => x"C0C0C0C0B0F980A4",
  3183 => x"C0C0C0C0B0F980B0",
  3184 => x"C0C0C0C0B0F98099",
  3185 => x"C0C0C0C0B0F98092",
  3186 => x"C0C0C0C0B0F98082",
  3187 => x"C0C0C0C0B0F980F8",
  3188 => x"C0C0C0C0B0F98080",
  3189 => x"C0C0C0C0B0F98090",
  3190 => x"C0C0C0C0B0F990C0",
  3191 => x"C0C0C0C0B0F990F9",
  3192 => x"C0C0C0C0B0F990A4",
  3193 => x"C0C0C0C0B0F990B0",
  3194 => x"C0C0C0C0B0F99099",
  3195 => x"C0C0C0C0B0F99092",
  3196 => x"C0C0C0C0B0F99082",
  3197 => x"C0C0C0C0B0F990F8",
  3198 => x"C0C0C0C0B0F99080",
  3199 => x"C0C0C0C0B0F99090",
  3200 => x"C0C0C0C0B0A4C0C0",
  3201 => x"C0C0C0C0B0A4C0F9",
  3202 => x"C0C0C0C0B0A4C0A4",
  3203 => x"C0C0C0C0B0A4C0B0",
  3204 => x"C0C0C0C0B0A4C099",
  3205 => x"C0C0C0C0B0A4C092",
  3206 => x"C0C0C0C0B0A4C082",
  3207 => x"C0C0C0C0B0A4C0F8",
  3208 => x"C0C0C0C0B0A4C080",
  3209 => x"C0C0C0C0B0A4C090",
  3210 => x"C0C0C0C0B0A4F9C0",
  3211 => x"C0C0C0C0B0A4F9F9",
  3212 => x"C0C0C0C0B0A4F9A4",
  3213 => x"C0C0C0C0B0A4F9B0",
  3214 => x"C0C0C0C0B0A4F999",
  3215 => x"C0C0C0C0B0A4F992",
  3216 => x"C0C0C0C0B0A4F982",
  3217 => x"C0C0C0C0B0A4F9F8",
  3218 => x"C0C0C0C0B0A4F980",
  3219 => x"C0C0C0C0B0A4F990",
  3220 => x"C0C0C0C0B0A4A4C0",
  3221 => x"C0C0C0C0B0A4A4F9",
  3222 => x"C0C0C0C0B0A4A4A4",
  3223 => x"C0C0C0C0B0A4A4B0",
  3224 => x"C0C0C0C0B0A4A499",
  3225 => x"C0C0C0C0B0A4A492",
  3226 => x"C0C0C0C0B0A4A482",
  3227 => x"C0C0C0C0B0A4A4F8",
  3228 => x"C0C0C0C0B0A4A480",
  3229 => x"C0C0C0C0B0A4A490",
  3230 => x"C0C0C0C0B0A4B0C0",
  3231 => x"C0C0C0C0B0A4B0F9",
  3232 => x"C0C0C0C0B0A4B0A4",
  3233 => x"C0C0C0C0B0A4B0B0",
  3234 => x"C0C0C0C0B0A4B099",
  3235 => x"C0C0C0C0B0A4B092",
  3236 => x"C0C0C0C0B0A4B082",
  3237 => x"C0C0C0C0B0A4B0F8",
  3238 => x"C0C0C0C0B0A4B080",
  3239 => x"C0C0C0C0B0A4B090",
  3240 => x"C0C0C0C0B0A499C0",
  3241 => x"C0C0C0C0B0A499F9",
  3242 => x"C0C0C0C0B0A499A4",
  3243 => x"C0C0C0C0B0A499B0",
  3244 => x"C0C0C0C0B0A49999",
  3245 => x"C0C0C0C0B0A49992",
  3246 => x"C0C0C0C0B0A49982",
  3247 => x"C0C0C0C0B0A499F8",
  3248 => x"C0C0C0C0B0A49980",
  3249 => x"C0C0C0C0B0A49990",
  3250 => x"C0C0C0C0B0A492C0",
  3251 => x"C0C0C0C0B0A492F9",
  3252 => x"C0C0C0C0B0A492A4",
  3253 => x"C0C0C0C0B0A492B0",
  3254 => x"C0C0C0C0B0A49299",
  3255 => x"C0C0C0C0B0A49292",
  3256 => x"C0C0C0C0B0A49282",
  3257 => x"C0C0C0C0B0A492F8",
  3258 => x"C0C0C0C0B0A49280",
  3259 => x"C0C0C0C0B0A49290",
  3260 => x"C0C0C0C0B0A482C0",
  3261 => x"C0C0C0C0B0A482F9",
  3262 => x"C0C0C0C0B0A482A4",
  3263 => x"C0C0C0C0B0A482B0",
  3264 => x"C0C0C0C0B0A48299",
  3265 => x"C0C0C0C0B0A48292",
  3266 => x"C0C0C0C0B0A48282",
  3267 => x"C0C0C0C0B0A482F8",
  3268 => x"C0C0C0C0B0A48280",
  3269 => x"C0C0C0C0B0A48290",
  3270 => x"C0C0C0C0B0A4F8C0",
  3271 => x"C0C0C0C0B0A4F8F9",
  3272 => x"C0C0C0C0B0A4F8A4",
  3273 => x"C0C0C0C0B0A4F8B0",
  3274 => x"C0C0C0C0B0A4F899",
  3275 => x"C0C0C0C0B0A4F892",
  3276 => x"C0C0C0C0B0A4F882",
  3277 => x"C0C0C0C0B0A4F8F8",
  3278 => x"C0C0C0C0B0A4F880",
  3279 => x"C0C0C0C0B0A4F890",
  3280 => x"C0C0C0C0B0A480C0",
  3281 => x"C0C0C0C0B0A480F9",
  3282 => x"C0C0C0C0B0A480A4",
  3283 => x"C0C0C0C0B0A480B0",
  3284 => x"C0C0C0C0B0A48099",
  3285 => x"C0C0C0C0B0A48092",
  3286 => x"C0C0C0C0B0A48082",
  3287 => x"C0C0C0C0B0A480F8",
  3288 => x"C0C0C0C0B0A48080",
  3289 => x"C0C0C0C0B0A48090",
  3290 => x"C0C0C0C0B0A490C0",
  3291 => x"C0C0C0C0B0A490F9",
  3292 => x"C0C0C0C0B0A490A4",
  3293 => x"C0C0C0C0B0A490B0",
  3294 => x"C0C0C0C0B0A49099",
  3295 => x"C0C0C0C0B0A49092",
  3296 => x"C0C0C0C0B0A49082",
  3297 => x"C0C0C0C0B0A490F8",
  3298 => x"C0C0C0C0B0A49080",
  3299 => x"C0C0C0C0B0A49090",
  3300 => x"C0C0C0C0B0B0C0C0",
  3301 => x"C0C0C0C0B0B0C0F9",
  3302 => x"C0C0C0C0B0B0C0A4",
  3303 => x"C0C0C0C0B0B0C0B0",
  3304 => x"C0C0C0C0B0B0C099",
  3305 => x"C0C0C0C0B0B0C092",
  3306 => x"C0C0C0C0B0B0C082",
  3307 => x"C0C0C0C0B0B0C0F8",
  3308 => x"C0C0C0C0B0B0C080",
  3309 => x"C0C0C0C0B0B0C090",
  3310 => x"C0C0C0C0B0B0F9C0",
  3311 => x"C0C0C0C0B0B0F9F9",
  3312 => x"C0C0C0C0B0B0F9A4",
  3313 => x"C0C0C0C0B0B0F9B0",
  3314 => x"C0C0C0C0B0B0F999",
  3315 => x"C0C0C0C0B0B0F992",
  3316 => x"C0C0C0C0B0B0F982",
  3317 => x"C0C0C0C0B0B0F9F8",
  3318 => x"C0C0C0C0B0B0F980",
  3319 => x"C0C0C0C0B0B0F990",
  3320 => x"C0C0C0C0B0B0A4C0",
  3321 => x"C0C0C0C0B0B0A4F9",
  3322 => x"C0C0C0C0B0B0A4A4",
  3323 => x"C0C0C0C0B0B0A4B0",
  3324 => x"C0C0C0C0B0B0A499",
  3325 => x"C0C0C0C0B0B0A492",
  3326 => x"C0C0C0C0B0B0A482",
  3327 => x"C0C0C0C0B0B0A4F8",
  3328 => x"C0C0C0C0B0B0A480",
  3329 => x"C0C0C0C0B0B0A490",
  3330 => x"C0C0C0C0B0B0B0C0",
  3331 => x"C0C0C0C0B0B0B0F9",
  3332 => x"C0C0C0C0B0B0B0A4",
  3333 => x"C0C0C0C0B0B0B0B0",
  3334 => x"C0C0C0C0B0B0B099",
  3335 => x"C0C0C0C0B0B0B092",
  3336 => x"C0C0C0C0B0B0B082",
  3337 => x"C0C0C0C0B0B0B0F8",
  3338 => x"C0C0C0C0B0B0B080",
  3339 => x"C0C0C0C0B0B0B090",
  3340 => x"C0C0C0C0B0B099C0",
  3341 => x"C0C0C0C0B0B099F9",
  3342 => x"C0C0C0C0B0B099A4",
  3343 => x"C0C0C0C0B0B099B0",
  3344 => x"C0C0C0C0B0B09999",
  3345 => x"C0C0C0C0B0B09992",
  3346 => x"C0C0C0C0B0B09982",
  3347 => x"C0C0C0C0B0B099F8",
  3348 => x"C0C0C0C0B0B09980",
  3349 => x"C0C0C0C0B0B09990",
  3350 => x"C0C0C0C0B0B092C0",
  3351 => x"C0C0C0C0B0B092F9",
  3352 => x"C0C0C0C0B0B092A4",
  3353 => x"C0C0C0C0B0B092B0",
  3354 => x"C0C0C0C0B0B09299",
  3355 => x"C0C0C0C0B0B09292",
  3356 => x"C0C0C0C0B0B09282",
  3357 => x"C0C0C0C0B0B092F8",
  3358 => x"C0C0C0C0B0B09280",
  3359 => x"C0C0C0C0B0B09290",
  3360 => x"C0C0C0C0B0B082C0",
  3361 => x"C0C0C0C0B0B082F9",
  3362 => x"C0C0C0C0B0B082A4",
  3363 => x"C0C0C0C0B0B082B0",
  3364 => x"C0C0C0C0B0B08299",
  3365 => x"C0C0C0C0B0B08292",
  3366 => x"C0C0C0C0B0B08282",
  3367 => x"C0C0C0C0B0B082F8",
  3368 => x"C0C0C0C0B0B08280",
  3369 => x"C0C0C0C0B0B08290",
  3370 => x"C0C0C0C0B0B0F8C0",
  3371 => x"C0C0C0C0B0B0F8F9",
  3372 => x"C0C0C0C0B0B0F8A4",
  3373 => x"C0C0C0C0B0B0F8B0",
  3374 => x"C0C0C0C0B0B0F899",
  3375 => x"C0C0C0C0B0B0F892",
  3376 => x"C0C0C0C0B0B0F882",
  3377 => x"C0C0C0C0B0B0F8F8",
  3378 => x"C0C0C0C0B0B0F880",
  3379 => x"C0C0C0C0B0B0F890",
  3380 => x"C0C0C0C0B0B080C0",
  3381 => x"C0C0C0C0B0B080F9",
  3382 => x"C0C0C0C0B0B080A4",
  3383 => x"C0C0C0C0B0B080B0",
  3384 => x"C0C0C0C0B0B08099",
  3385 => x"C0C0C0C0B0B08092",
  3386 => x"C0C0C0C0B0B08082",
  3387 => x"C0C0C0C0B0B080F8",
  3388 => x"C0C0C0C0B0B08080",
  3389 => x"C0C0C0C0B0B08090",
  3390 => x"C0C0C0C0B0B090C0",
  3391 => x"C0C0C0C0B0B090F9",
  3392 => x"C0C0C0C0B0B090A4",
  3393 => x"C0C0C0C0B0B090B0",
  3394 => x"C0C0C0C0B0B09099",
  3395 => x"C0C0C0C0B0B09092",
  3396 => x"C0C0C0C0B0B09082",
  3397 => x"C0C0C0C0B0B090F8",
  3398 => x"C0C0C0C0B0B09080",
  3399 => x"C0C0C0C0B0B09090",
  3400 => x"C0C0C0C0B099C0C0",
  3401 => x"C0C0C0C0B099C0F9",
  3402 => x"C0C0C0C0B099C0A4",
  3403 => x"C0C0C0C0B099C0B0",
  3404 => x"C0C0C0C0B099C099",
  3405 => x"C0C0C0C0B099C092",
  3406 => x"C0C0C0C0B099C082",
  3407 => x"C0C0C0C0B099C0F8",
  3408 => x"C0C0C0C0B099C080",
  3409 => x"C0C0C0C0B099C090",
  3410 => x"C0C0C0C0B099F9C0",
  3411 => x"C0C0C0C0B099F9F9",
  3412 => x"C0C0C0C0B099F9A4",
  3413 => x"C0C0C0C0B099F9B0",
  3414 => x"C0C0C0C0B099F999",
  3415 => x"C0C0C0C0B099F992",
  3416 => x"C0C0C0C0B099F982",
  3417 => x"C0C0C0C0B099F9F8",
  3418 => x"C0C0C0C0B099F980",
  3419 => x"C0C0C0C0B099F990",
  3420 => x"C0C0C0C0B099A4C0",
  3421 => x"C0C0C0C0B099A4F9",
  3422 => x"C0C0C0C0B099A4A4",
  3423 => x"C0C0C0C0B099A4B0",
  3424 => x"C0C0C0C0B099A499",
  3425 => x"C0C0C0C0B099A492",
  3426 => x"C0C0C0C0B099A482",
  3427 => x"C0C0C0C0B099A4F8",
  3428 => x"C0C0C0C0B099A480",
  3429 => x"C0C0C0C0B099A490",
  3430 => x"C0C0C0C0B099B0C0",
  3431 => x"C0C0C0C0B099B0F9",
  3432 => x"C0C0C0C0B099B0A4",
  3433 => x"C0C0C0C0B099B0B0",
  3434 => x"C0C0C0C0B099B099",
  3435 => x"C0C0C0C0B099B092",
  3436 => x"C0C0C0C0B099B082",
  3437 => x"C0C0C0C0B099B0F8",
  3438 => x"C0C0C0C0B099B080",
  3439 => x"C0C0C0C0B099B090",
  3440 => x"C0C0C0C0B09999C0",
  3441 => x"C0C0C0C0B09999F9",
  3442 => x"C0C0C0C0B09999A4",
  3443 => x"C0C0C0C0B09999B0",
  3444 => x"C0C0C0C0B0999999",
  3445 => x"C0C0C0C0B0999992",
  3446 => x"C0C0C0C0B0999982",
  3447 => x"C0C0C0C0B09999F8",
  3448 => x"C0C0C0C0B0999980",
  3449 => x"C0C0C0C0B0999990",
  3450 => x"C0C0C0C0B09992C0",
  3451 => x"C0C0C0C0B09992F9",
  3452 => x"C0C0C0C0B09992A4",
  3453 => x"C0C0C0C0B09992B0",
  3454 => x"C0C0C0C0B0999299",
  3455 => x"C0C0C0C0B0999292",
  3456 => x"C0C0C0C0B0999282",
  3457 => x"C0C0C0C0B09992F8",
  3458 => x"C0C0C0C0B0999280",
  3459 => x"C0C0C0C0B0999290",
  3460 => x"C0C0C0C0B09982C0",
  3461 => x"C0C0C0C0B09982F9",
  3462 => x"C0C0C0C0B09982A4",
  3463 => x"C0C0C0C0B09982B0",
  3464 => x"C0C0C0C0B0998299",
  3465 => x"C0C0C0C0B0998292",
  3466 => x"C0C0C0C0B0998282",
  3467 => x"C0C0C0C0B09982F8",
  3468 => x"C0C0C0C0B0998280",
  3469 => x"C0C0C0C0B0998290",
  3470 => x"C0C0C0C0B099F8C0",
  3471 => x"C0C0C0C0B099F8F9",
  3472 => x"C0C0C0C0B099F8A4",
  3473 => x"C0C0C0C0B099F8B0",
  3474 => x"C0C0C0C0B099F899",
  3475 => x"C0C0C0C0B099F892",
  3476 => x"C0C0C0C0B099F882",
  3477 => x"C0C0C0C0B099F8F8",
  3478 => x"C0C0C0C0B099F880",
  3479 => x"C0C0C0C0B099F890",
  3480 => x"C0C0C0C0B09980C0",
  3481 => x"C0C0C0C0B09980F9",
  3482 => x"C0C0C0C0B09980A4",
  3483 => x"C0C0C0C0B09980B0",
  3484 => x"C0C0C0C0B0998099",
  3485 => x"C0C0C0C0B0998092",
  3486 => x"C0C0C0C0B0998082",
  3487 => x"C0C0C0C0B09980F8",
  3488 => x"C0C0C0C0B0998080",
  3489 => x"C0C0C0C0B0998090",
  3490 => x"C0C0C0C0B09990C0",
  3491 => x"C0C0C0C0B09990F9",
  3492 => x"C0C0C0C0B09990A4",
  3493 => x"C0C0C0C0B09990B0",
  3494 => x"C0C0C0C0B0999099",
  3495 => x"C0C0C0C0B0999092",
  3496 => x"C0C0C0C0B0999082",
  3497 => x"C0C0C0C0B09990F8",
  3498 => x"C0C0C0C0B0999080",
  3499 => x"C0C0C0C0B0999090",
  3500 => x"C0C0C0C0B092C0C0",
  3501 => x"C0C0C0C0B092C0F9",
  3502 => x"C0C0C0C0B092C0A4",
  3503 => x"C0C0C0C0B092C0B0",
  3504 => x"C0C0C0C0B092C099",
  3505 => x"C0C0C0C0B092C092",
  3506 => x"C0C0C0C0B092C082",
  3507 => x"C0C0C0C0B092C0F8",
  3508 => x"C0C0C0C0B092C080",
  3509 => x"C0C0C0C0B092C090",
  3510 => x"C0C0C0C0B092F9C0",
  3511 => x"C0C0C0C0B092F9F9",
  3512 => x"C0C0C0C0B092F9A4",
  3513 => x"C0C0C0C0B092F9B0",
  3514 => x"C0C0C0C0B092F999",
  3515 => x"C0C0C0C0B092F992",
  3516 => x"C0C0C0C0B092F982",
  3517 => x"C0C0C0C0B092F9F8",
  3518 => x"C0C0C0C0B092F980",
  3519 => x"C0C0C0C0B092F990",
  3520 => x"C0C0C0C0B092A4C0",
  3521 => x"C0C0C0C0B092A4F9",
  3522 => x"C0C0C0C0B092A4A4",
  3523 => x"C0C0C0C0B092A4B0",
  3524 => x"C0C0C0C0B092A499",
  3525 => x"C0C0C0C0B092A492",
  3526 => x"C0C0C0C0B092A482",
  3527 => x"C0C0C0C0B092A4F8",
  3528 => x"C0C0C0C0B092A480",
  3529 => x"C0C0C0C0B092A490",
  3530 => x"C0C0C0C0B092B0C0",
  3531 => x"C0C0C0C0B092B0F9",
  3532 => x"C0C0C0C0B092B0A4",
  3533 => x"C0C0C0C0B092B0B0",
  3534 => x"C0C0C0C0B092B099",
  3535 => x"C0C0C0C0B092B092",
  3536 => x"C0C0C0C0B092B082",
  3537 => x"C0C0C0C0B092B0F8",
  3538 => x"C0C0C0C0B092B080",
  3539 => x"C0C0C0C0B092B090",
  3540 => x"C0C0C0C0B09299C0",
  3541 => x"C0C0C0C0B09299F9",
  3542 => x"C0C0C0C0B09299A4",
  3543 => x"C0C0C0C0B09299B0",
  3544 => x"C0C0C0C0B0929999",
  3545 => x"C0C0C0C0B0929992",
  3546 => x"C0C0C0C0B0929982",
  3547 => x"C0C0C0C0B09299F8",
  3548 => x"C0C0C0C0B0929980",
  3549 => x"C0C0C0C0B0929990",
  3550 => x"C0C0C0C0B09292C0",
  3551 => x"C0C0C0C0B09292F9",
  3552 => x"C0C0C0C0B09292A4",
  3553 => x"C0C0C0C0B09292B0",
  3554 => x"C0C0C0C0B0929299",
  3555 => x"C0C0C0C0B0929292",
  3556 => x"C0C0C0C0B0929282",
  3557 => x"C0C0C0C0B09292F8",
  3558 => x"C0C0C0C0B0929280",
  3559 => x"C0C0C0C0B0929290",
  3560 => x"C0C0C0C0B09282C0",
  3561 => x"C0C0C0C0B09282F9",
  3562 => x"C0C0C0C0B09282A4",
  3563 => x"C0C0C0C0B09282B0",
  3564 => x"C0C0C0C0B0928299",
  3565 => x"C0C0C0C0B0928292",
  3566 => x"C0C0C0C0B0928282",
  3567 => x"C0C0C0C0B09282F8",
  3568 => x"C0C0C0C0B0928280",
  3569 => x"C0C0C0C0B0928290",
  3570 => x"C0C0C0C0B092F8C0",
  3571 => x"C0C0C0C0B092F8F9",
  3572 => x"C0C0C0C0B092F8A4",
  3573 => x"C0C0C0C0B092F8B0",
  3574 => x"C0C0C0C0B092F899",
  3575 => x"C0C0C0C0B092F892",
  3576 => x"C0C0C0C0B092F882",
  3577 => x"C0C0C0C0B092F8F8",
  3578 => x"C0C0C0C0B092F880",
  3579 => x"C0C0C0C0B092F890",
  3580 => x"C0C0C0C0B09280C0",
  3581 => x"C0C0C0C0B09280F9",
  3582 => x"C0C0C0C0B09280A4",
  3583 => x"C0C0C0C0B09280B0",
  3584 => x"C0C0C0C0B0928099",
  3585 => x"C0C0C0C0B0928092",
  3586 => x"C0C0C0C0B0928082",
  3587 => x"C0C0C0C0B09280F8",
  3588 => x"C0C0C0C0B0928080",
  3589 => x"C0C0C0C0B0928090",
  3590 => x"C0C0C0C0B09290C0",
  3591 => x"C0C0C0C0B09290F9",
  3592 => x"C0C0C0C0B09290A4",
  3593 => x"C0C0C0C0B09290B0",
  3594 => x"C0C0C0C0B0929099",
  3595 => x"C0C0C0C0B0929092",
  3596 => x"C0C0C0C0B0929082",
  3597 => x"C0C0C0C0B09290F8",
  3598 => x"C0C0C0C0B0929080",
  3599 => x"C0C0C0C0B0929090",
  3600 => x"C0C0C0C0B082C0C0",
  3601 => x"C0C0C0C0B082C0F9",
  3602 => x"C0C0C0C0B082C0A4",
  3603 => x"C0C0C0C0B082C0B0",
  3604 => x"C0C0C0C0B082C099",
  3605 => x"C0C0C0C0B082C092",
  3606 => x"C0C0C0C0B082C082",
  3607 => x"C0C0C0C0B082C0F8",
  3608 => x"C0C0C0C0B082C080",
  3609 => x"C0C0C0C0B082C090",
  3610 => x"C0C0C0C0B082F9C0",
  3611 => x"C0C0C0C0B082F9F9",
  3612 => x"C0C0C0C0B082F9A4",
  3613 => x"C0C0C0C0B082F9B0",
  3614 => x"C0C0C0C0B082F999",
  3615 => x"C0C0C0C0B082F992",
  3616 => x"C0C0C0C0B082F982",
  3617 => x"C0C0C0C0B082F9F8",
  3618 => x"C0C0C0C0B082F980",
  3619 => x"C0C0C0C0B082F990",
  3620 => x"C0C0C0C0B082A4C0",
  3621 => x"C0C0C0C0B082A4F9",
  3622 => x"C0C0C0C0B082A4A4",
  3623 => x"C0C0C0C0B082A4B0",
  3624 => x"C0C0C0C0B082A499",
  3625 => x"C0C0C0C0B082A492",
  3626 => x"C0C0C0C0B082A482",
  3627 => x"C0C0C0C0B082A4F8",
  3628 => x"C0C0C0C0B082A480",
  3629 => x"C0C0C0C0B082A490",
  3630 => x"C0C0C0C0B082B0C0",
  3631 => x"C0C0C0C0B082B0F9",
  3632 => x"C0C0C0C0B082B0A4",
  3633 => x"C0C0C0C0B082B0B0",
  3634 => x"C0C0C0C0B082B099",
  3635 => x"C0C0C0C0B082B092",
  3636 => x"C0C0C0C0B082B082",
  3637 => x"C0C0C0C0B082B0F8",
  3638 => x"C0C0C0C0B082B080",
  3639 => x"C0C0C0C0B082B090",
  3640 => x"C0C0C0C0B08299C0",
  3641 => x"C0C0C0C0B08299F9",
  3642 => x"C0C0C0C0B08299A4",
  3643 => x"C0C0C0C0B08299B0",
  3644 => x"C0C0C0C0B0829999",
  3645 => x"C0C0C0C0B0829992",
  3646 => x"C0C0C0C0B0829982",
  3647 => x"C0C0C0C0B08299F8",
  3648 => x"C0C0C0C0B0829980",
  3649 => x"C0C0C0C0B0829990",
  3650 => x"C0C0C0C0B08292C0",
  3651 => x"C0C0C0C0B08292F9",
  3652 => x"C0C0C0C0B08292A4",
  3653 => x"C0C0C0C0B08292B0",
  3654 => x"C0C0C0C0B0829299",
  3655 => x"C0C0C0C0B0829292",
  3656 => x"C0C0C0C0B0829282",
  3657 => x"C0C0C0C0B08292F8",
  3658 => x"C0C0C0C0B0829280",
  3659 => x"C0C0C0C0B0829290",
  3660 => x"C0C0C0C0B08282C0",
  3661 => x"C0C0C0C0B08282F9",
  3662 => x"C0C0C0C0B08282A4",
  3663 => x"C0C0C0C0B08282B0",
  3664 => x"C0C0C0C0B0828299",
  3665 => x"C0C0C0C0B0828292",
  3666 => x"C0C0C0C0B0828282",
  3667 => x"C0C0C0C0B08282F8",
  3668 => x"C0C0C0C0B0828280",
  3669 => x"C0C0C0C0B0828290",
  3670 => x"C0C0C0C0B082F8C0",
  3671 => x"C0C0C0C0B082F8F9",
  3672 => x"C0C0C0C0B082F8A4",
  3673 => x"C0C0C0C0B082F8B0",
  3674 => x"C0C0C0C0B082F899",
  3675 => x"C0C0C0C0B082F892",
  3676 => x"C0C0C0C0B082F882",
  3677 => x"C0C0C0C0B082F8F8",
  3678 => x"C0C0C0C0B082F880",
  3679 => x"C0C0C0C0B082F890",
  3680 => x"C0C0C0C0B08280C0",
  3681 => x"C0C0C0C0B08280F9",
  3682 => x"C0C0C0C0B08280A4",
  3683 => x"C0C0C0C0B08280B0",
  3684 => x"C0C0C0C0B0828099",
  3685 => x"C0C0C0C0B0828092",
  3686 => x"C0C0C0C0B0828082",
  3687 => x"C0C0C0C0B08280F8",
  3688 => x"C0C0C0C0B0828080",
  3689 => x"C0C0C0C0B0828090",
  3690 => x"C0C0C0C0B08290C0",
  3691 => x"C0C0C0C0B08290F9",
  3692 => x"C0C0C0C0B08290A4",
  3693 => x"C0C0C0C0B08290B0",
  3694 => x"C0C0C0C0B0829099",
  3695 => x"C0C0C0C0B0829092",
  3696 => x"C0C0C0C0B0829082",
  3697 => x"C0C0C0C0B08290F8",
  3698 => x"C0C0C0C0B0829080",
  3699 => x"C0C0C0C0B0829090",
  3700 => x"C0C0C0C0B0F8C0C0",
  3701 => x"C0C0C0C0B0F8C0F9",
  3702 => x"C0C0C0C0B0F8C0A4",
  3703 => x"C0C0C0C0B0F8C0B0",
  3704 => x"C0C0C0C0B0F8C099",
  3705 => x"C0C0C0C0B0F8C092",
  3706 => x"C0C0C0C0B0F8C082",
  3707 => x"C0C0C0C0B0F8C0F8",
  3708 => x"C0C0C0C0B0F8C080",
  3709 => x"C0C0C0C0B0F8C090",
  3710 => x"C0C0C0C0B0F8F9C0",
  3711 => x"C0C0C0C0B0F8F9F9",
  3712 => x"C0C0C0C0B0F8F9A4",
  3713 => x"C0C0C0C0B0F8F9B0",
  3714 => x"C0C0C0C0B0F8F999",
  3715 => x"C0C0C0C0B0F8F992",
  3716 => x"C0C0C0C0B0F8F982",
  3717 => x"C0C0C0C0B0F8F9F8",
  3718 => x"C0C0C0C0B0F8F980",
  3719 => x"C0C0C0C0B0F8F990",
  3720 => x"C0C0C0C0B0F8A4C0",
  3721 => x"C0C0C0C0B0F8A4F9",
  3722 => x"C0C0C0C0B0F8A4A4",
  3723 => x"C0C0C0C0B0F8A4B0",
  3724 => x"C0C0C0C0B0F8A499",
  3725 => x"C0C0C0C0B0F8A492",
  3726 => x"C0C0C0C0B0F8A482",
  3727 => x"C0C0C0C0B0F8A4F8",
  3728 => x"C0C0C0C0B0F8A480",
  3729 => x"C0C0C0C0B0F8A490",
  3730 => x"C0C0C0C0B0F8B0C0",
  3731 => x"C0C0C0C0B0F8B0F9",
  3732 => x"C0C0C0C0B0F8B0A4",
  3733 => x"C0C0C0C0B0F8B0B0",
  3734 => x"C0C0C0C0B0F8B099",
  3735 => x"C0C0C0C0B0F8B092",
  3736 => x"C0C0C0C0B0F8B082",
  3737 => x"C0C0C0C0B0F8B0F8",
  3738 => x"C0C0C0C0B0F8B080",
  3739 => x"C0C0C0C0B0F8B090",
  3740 => x"C0C0C0C0B0F899C0",
  3741 => x"C0C0C0C0B0F899F9",
  3742 => x"C0C0C0C0B0F899A4",
  3743 => x"C0C0C0C0B0F899B0",
  3744 => x"C0C0C0C0B0F89999",
  3745 => x"C0C0C0C0B0F89992",
  3746 => x"C0C0C0C0B0F89982",
  3747 => x"C0C0C0C0B0F899F8",
  3748 => x"C0C0C0C0B0F89980",
  3749 => x"C0C0C0C0B0F89990",
  3750 => x"C0C0C0C0B0F892C0",
  3751 => x"C0C0C0C0B0F892F9",
  3752 => x"C0C0C0C0B0F892A4",
  3753 => x"C0C0C0C0B0F892B0",
  3754 => x"C0C0C0C0B0F89299",
  3755 => x"C0C0C0C0B0F89292",
  3756 => x"C0C0C0C0B0F89282",
  3757 => x"C0C0C0C0B0F892F8",
  3758 => x"C0C0C0C0B0F89280",
  3759 => x"C0C0C0C0B0F89290",
  3760 => x"C0C0C0C0B0F882C0",
  3761 => x"C0C0C0C0B0F882F9",
  3762 => x"C0C0C0C0B0F882A4",
  3763 => x"C0C0C0C0B0F882B0",
  3764 => x"C0C0C0C0B0F88299",
  3765 => x"C0C0C0C0B0F88292",
  3766 => x"C0C0C0C0B0F88282",
  3767 => x"C0C0C0C0B0F882F8",
  3768 => x"C0C0C0C0B0F88280",
  3769 => x"C0C0C0C0B0F88290",
  3770 => x"C0C0C0C0B0F8F8C0",
  3771 => x"C0C0C0C0B0F8F8F9",
  3772 => x"C0C0C0C0B0F8F8A4",
  3773 => x"C0C0C0C0B0F8F8B0",
  3774 => x"C0C0C0C0B0F8F899",
  3775 => x"C0C0C0C0B0F8F892",
  3776 => x"C0C0C0C0B0F8F882",
  3777 => x"C0C0C0C0B0F8F8F8",
  3778 => x"C0C0C0C0B0F8F880",
  3779 => x"C0C0C0C0B0F8F890",
  3780 => x"C0C0C0C0B0F880C0",
  3781 => x"C0C0C0C0B0F880F9",
  3782 => x"C0C0C0C0B0F880A4",
  3783 => x"C0C0C0C0B0F880B0",
  3784 => x"C0C0C0C0B0F88099",
  3785 => x"C0C0C0C0B0F88092",
  3786 => x"C0C0C0C0B0F88082",
  3787 => x"C0C0C0C0B0F880F8",
  3788 => x"C0C0C0C0B0F88080",
  3789 => x"C0C0C0C0B0F88090",
  3790 => x"C0C0C0C0B0F890C0",
  3791 => x"C0C0C0C0B0F890F9",
  3792 => x"C0C0C0C0B0F890A4",
  3793 => x"C0C0C0C0B0F890B0",
  3794 => x"C0C0C0C0B0F89099",
  3795 => x"C0C0C0C0B0F89092",
  3796 => x"C0C0C0C0B0F89082",
  3797 => x"C0C0C0C0B0F890F8",
  3798 => x"C0C0C0C0B0F89080",
  3799 => x"C0C0C0C0B0F89090",
  3800 => x"C0C0C0C0B080C0C0",
  3801 => x"C0C0C0C0B080C0F9",
  3802 => x"C0C0C0C0B080C0A4",
  3803 => x"C0C0C0C0B080C0B0",
  3804 => x"C0C0C0C0B080C099",
  3805 => x"C0C0C0C0B080C092",
  3806 => x"C0C0C0C0B080C082",
  3807 => x"C0C0C0C0B080C0F8",
  3808 => x"C0C0C0C0B080C080",
  3809 => x"C0C0C0C0B080C090",
  3810 => x"C0C0C0C0B080F9C0",
  3811 => x"C0C0C0C0B080F9F9",
  3812 => x"C0C0C0C0B080F9A4",
  3813 => x"C0C0C0C0B080F9B0",
  3814 => x"C0C0C0C0B080F999",
  3815 => x"C0C0C0C0B080F992",
  3816 => x"C0C0C0C0B080F982",
  3817 => x"C0C0C0C0B080F9F8",
  3818 => x"C0C0C0C0B080F980",
  3819 => x"C0C0C0C0B080F990",
  3820 => x"C0C0C0C0B080A4C0",
  3821 => x"C0C0C0C0B080A4F9",
  3822 => x"C0C0C0C0B080A4A4",
  3823 => x"C0C0C0C0B080A4B0",
  3824 => x"C0C0C0C0B080A499",
  3825 => x"C0C0C0C0B080A492",
  3826 => x"C0C0C0C0B080A482",
  3827 => x"C0C0C0C0B080A4F8",
  3828 => x"C0C0C0C0B080A480",
  3829 => x"C0C0C0C0B080A490",
  3830 => x"C0C0C0C0B080B0C0",
  3831 => x"C0C0C0C0B080B0F9",
  3832 => x"C0C0C0C0B080B0A4",
  3833 => x"C0C0C0C0B080B0B0",
  3834 => x"C0C0C0C0B080B099",
  3835 => x"C0C0C0C0B080B092",
  3836 => x"C0C0C0C0B080B082",
  3837 => x"C0C0C0C0B080B0F8",
  3838 => x"C0C0C0C0B080B080",
  3839 => x"C0C0C0C0B080B090",
  3840 => x"C0C0C0C0B08099C0",
  3841 => x"C0C0C0C0B08099F9",
  3842 => x"C0C0C0C0B08099A4",
  3843 => x"C0C0C0C0B08099B0",
  3844 => x"C0C0C0C0B0809999",
  3845 => x"C0C0C0C0B0809992",
  3846 => x"C0C0C0C0B0809982",
  3847 => x"C0C0C0C0B08099F8",
  3848 => x"C0C0C0C0B0809980",
  3849 => x"C0C0C0C0B0809990",
  3850 => x"C0C0C0C0B08092C0",
  3851 => x"C0C0C0C0B08092F9",
  3852 => x"C0C0C0C0B08092A4",
  3853 => x"C0C0C0C0B08092B0",
  3854 => x"C0C0C0C0B0809299",
  3855 => x"C0C0C0C0B0809292",
  3856 => x"C0C0C0C0B0809282",
  3857 => x"C0C0C0C0B08092F8",
  3858 => x"C0C0C0C0B0809280",
  3859 => x"C0C0C0C0B0809290",
  3860 => x"C0C0C0C0B08082C0",
  3861 => x"C0C0C0C0B08082F9",
  3862 => x"C0C0C0C0B08082A4",
  3863 => x"C0C0C0C0B08082B0",
  3864 => x"C0C0C0C0B0808299",
  3865 => x"C0C0C0C0B0808292",
  3866 => x"C0C0C0C0B0808282",
  3867 => x"C0C0C0C0B08082F8",
  3868 => x"C0C0C0C0B0808280",
  3869 => x"C0C0C0C0B0808290",
  3870 => x"C0C0C0C0B080F8C0",
  3871 => x"C0C0C0C0B080F8F9",
  3872 => x"C0C0C0C0B080F8A4",
  3873 => x"C0C0C0C0B080F8B0",
  3874 => x"C0C0C0C0B080F899",
  3875 => x"C0C0C0C0B080F892",
  3876 => x"C0C0C0C0B080F882",
  3877 => x"C0C0C0C0B080F8F8",
  3878 => x"C0C0C0C0B080F880",
  3879 => x"C0C0C0C0B080F890",
  3880 => x"C0C0C0C0B08080C0",
  3881 => x"C0C0C0C0B08080F9",
  3882 => x"C0C0C0C0B08080A4",
  3883 => x"C0C0C0C0B08080B0",
  3884 => x"C0C0C0C0B0808099",
  3885 => x"C0C0C0C0B0808092",
  3886 => x"C0C0C0C0B0808082",
  3887 => x"C0C0C0C0B08080F8",
  3888 => x"C0C0C0C0B0808080",
  3889 => x"C0C0C0C0B0808090",
  3890 => x"C0C0C0C0B08090C0",
  3891 => x"C0C0C0C0B08090F9",
  3892 => x"C0C0C0C0B08090A4",
  3893 => x"C0C0C0C0B08090B0",
  3894 => x"C0C0C0C0B0809099",
  3895 => x"C0C0C0C0B0809092",
  3896 => x"C0C0C0C0B0809082",
  3897 => x"C0C0C0C0B08090F8",
  3898 => x"C0C0C0C0B0809080",
  3899 => x"C0C0C0C0B0809090",
  3900 => x"C0C0C0C0B090C0C0",
  3901 => x"C0C0C0C0B090C0F9",
  3902 => x"C0C0C0C0B090C0A4",
  3903 => x"C0C0C0C0B090C0B0",
  3904 => x"C0C0C0C0B090C099",
  3905 => x"C0C0C0C0B090C092",
  3906 => x"C0C0C0C0B090C082",
  3907 => x"C0C0C0C0B090C0F8",
  3908 => x"C0C0C0C0B090C080",
  3909 => x"C0C0C0C0B090C090",
  3910 => x"C0C0C0C0B090F9C0",
  3911 => x"C0C0C0C0B090F9F9",
  3912 => x"C0C0C0C0B090F9A4",
  3913 => x"C0C0C0C0B090F9B0",
  3914 => x"C0C0C0C0B090F999",
  3915 => x"C0C0C0C0B090F992",
  3916 => x"C0C0C0C0B090F982",
  3917 => x"C0C0C0C0B090F9F8",
  3918 => x"C0C0C0C0B090F980",
  3919 => x"C0C0C0C0B090F990",
  3920 => x"C0C0C0C0B090A4C0",
  3921 => x"C0C0C0C0B090A4F9",
  3922 => x"C0C0C0C0B090A4A4",
  3923 => x"C0C0C0C0B090A4B0",
  3924 => x"C0C0C0C0B090A499",
  3925 => x"C0C0C0C0B090A492",
  3926 => x"C0C0C0C0B090A482",
  3927 => x"C0C0C0C0B090A4F8",
  3928 => x"C0C0C0C0B090A480",
  3929 => x"C0C0C0C0B090A490",
  3930 => x"C0C0C0C0B090B0C0",
  3931 => x"C0C0C0C0B090B0F9",
  3932 => x"C0C0C0C0B090B0A4",
  3933 => x"C0C0C0C0B090B0B0",
  3934 => x"C0C0C0C0B090B099",
  3935 => x"C0C0C0C0B090B092",
  3936 => x"C0C0C0C0B090B082",
  3937 => x"C0C0C0C0B090B0F8",
  3938 => x"C0C0C0C0B090B080",
  3939 => x"C0C0C0C0B090B090",
  3940 => x"C0C0C0C0B09099C0",
  3941 => x"C0C0C0C0B09099F9",
  3942 => x"C0C0C0C0B09099A4",
  3943 => x"C0C0C0C0B09099B0",
  3944 => x"C0C0C0C0B0909999",
  3945 => x"C0C0C0C0B0909992",
  3946 => x"C0C0C0C0B0909982",
  3947 => x"C0C0C0C0B09099F8",
  3948 => x"C0C0C0C0B0909980",
  3949 => x"C0C0C0C0B0909990",
  3950 => x"C0C0C0C0B09092C0",
  3951 => x"C0C0C0C0B09092F9",
  3952 => x"C0C0C0C0B09092A4",
  3953 => x"C0C0C0C0B09092B0",
  3954 => x"C0C0C0C0B0909299",
  3955 => x"C0C0C0C0B0909292",
  3956 => x"C0C0C0C0B0909282",
  3957 => x"C0C0C0C0B09092F8",
  3958 => x"C0C0C0C0B0909280",
  3959 => x"C0C0C0C0B0909290",
  3960 => x"C0C0C0C0B09082C0",
  3961 => x"C0C0C0C0B09082F9",
  3962 => x"C0C0C0C0B09082A4",
  3963 => x"C0C0C0C0B09082B0",
  3964 => x"C0C0C0C0B0908299",
  3965 => x"C0C0C0C0B0908292",
  3966 => x"C0C0C0C0B0908282",
  3967 => x"C0C0C0C0B09082F8",
  3968 => x"C0C0C0C0B0908280",
  3969 => x"C0C0C0C0B0908290",
  3970 => x"C0C0C0C0B090F8C0",
  3971 => x"C0C0C0C0B090F8F9",
  3972 => x"C0C0C0C0B090F8A4",
  3973 => x"C0C0C0C0B090F8B0",
  3974 => x"C0C0C0C0B090F899",
  3975 => x"C0C0C0C0B090F892",
  3976 => x"C0C0C0C0B090F882",
  3977 => x"C0C0C0C0B090F8F8",
  3978 => x"C0C0C0C0B090F880",
  3979 => x"C0C0C0C0B090F890",
  3980 => x"C0C0C0C0B09080C0",
  3981 => x"C0C0C0C0B09080F9",
  3982 => x"C0C0C0C0B09080A4",
  3983 => x"C0C0C0C0B09080B0",
  3984 => x"C0C0C0C0B0908099",
  3985 => x"C0C0C0C0B0908092",
  3986 => x"C0C0C0C0B0908082",
  3987 => x"C0C0C0C0B09080F8",
  3988 => x"C0C0C0C0B0908080",
  3989 => x"C0C0C0C0B0908090",
  3990 => x"C0C0C0C0B09090C0",
  3991 => x"C0C0C0C0B09090F9",
  3992 => x"C0C0C0C0B09090A4",
  3993 => x"C0C0C0C0B09090B0",
  3994 => x"C0C0C0C0B0909099",
  3995 => x"C0C0C0C0B0909092",
  3996 => x"C0C0C0C0B0909082",
  3997 => x"C0C0C0C0B09090F8",
  3998 => x"C0C0C0C0B0909080",
  3999 => x"C0C0C0C0B0909090",
  4000 => x"C0C0C0C099C0C0C0",
  4001 => x"C0C0C0C099C0C0F9",
  4002 => x"C0C0C0C099C0C0A4",
  4003 => x"C0C0C0C099C0C0B0",
  4004 => x"C0C0C0C099C0C099",
  4005 => x"C0C0C0C099C0C092",
  4006 => x"C0C0C0C099C0C082",
  4007 => x"C0C0C0C099C0C0F8",
  4008 => x"C0C0C0C099C0C080",
  4009 => x"C0C0C0C099C0C090",
  4010 => x"C0C0C0C099C0F9C0",
  4011 => x"C0C0C0C099C0F9F9",
  4012 => x"C0C0C0C099C0F9A4",
  4013 => x"C0C0C0C099C0F9B0",
  4014 => x"C0C0C0C099C0F999",
  4015 => x"C0C0C0C099C0F992",
  4016 => x"C0C0C0C099C0F982",
  4017 => x"C0C0C0C099C0F9F8",
  4018 => x"C0C0C0C099C0F980",
  4019 => x"C0C0C0C099C0F990",
  4020 => x"C0C0C0C099C0A4C0",
  4021 => x"C0C0C0C099C0A4F9",
  4022 => x"C0C0C0C099C0A4A4",
  4023 => x"C0C0C0C099C0A4B0",
  4024 => x"C0C0C0C099C0A499",
  4025 => x"C0C0C0C099C0A492",
  4026 => x"C0C0C0C099C0A482",
  4027 => x"C0C0C0C099C0A4F8",
  4028 => x"C0C0C0C099C0A480",
  4029 => x"C0C0C0C099C0A490",
  4030 => x"C0C0C0C099C0B0C0",
  4031 => x"C0C0C0C099C0B0F9",
  4032 => x"C0C0C0C099C0B0A4",
  4033 => x"C0C0C0C099C0B0B0",
  4034 => x"C0C0C0C099C0B099",
  4035 => x"C0C0C0C099C0B092",
  4036 => x"C0C0C0C099C0B082",
  4037 => x"C0C0C0C099C0B0F8",
  4038 => x"C0C0C0C099C0B080",
  4039 => x"C0C0C0C099C0B090",
  4040 => x"C0C0C0C099C099C0",
  4041 => x"C0C0C0C099C099F9",
  4042 => x"C0C0C0C099C099A4",
  4043 => x"C0C0C0C099C099B0",
  4044 => x"C0C0C0C099C09999",
  4045 => x"C0C0C0C099C09992",
  4046 => x"C0C0C0C099C09982",
  4047 => x"C0C0C0C099C099F8",
  4048 => x"C0C0C0C099C09980",
  4049 => x"C0C0C0C099C09990",
  4050 => x"C0C0C0C099C092C0",
  4051 => x"C0C0C0C099C092F9",
  4052 => x"C0C0C0C099C092A4",
  4053 => x"C0C0C0C099C092B0",
  4054 => x"C0C0C0C099C09299",
  4055 => x"C0C0C0C099C09292",
  4056 => x"C0C0C0C099C09282",
  4057 => x"C0C0C0C099C092F8",
  4058 => x"C0C0C0C099C09280",
  4059 => x"C0C0C0C099C09290",
  4060 => x"C0C0C0C099C082C0",
  4061 => x"C0C0C0C099C082F9",
  4062 => x"C0C0C0C099C082A4",
  4063 => x"C0C0C0C099C082B0",
  4064 => x"C0C0C0C099C08299",
  4065 => x"C0C0C0C099C08292",
  4066 => x"C0C0C0C099C08282",
  4067 => x"C0C0C0C099C082F8",
  4068 => x"C0C0C0C099C08280",
  4069 => x"C0C0C0C099C08290",
  4070 => x"C0C0C0C099C0F8C0",
  4071 => x"C0C0C0C099C0F8F9",
  4072 => x"C0C0C0C099C0F8A4",
  4073 => x"C0C0C0C099C0F8B0",
  4074 => x"C0C0C0C099C0F899",
  4075 => x"C0C0C0C099C0F892",
  4076 => x"C0C0C0C099C0F882",
  4077 => x"C0C0C0C099C0F8F8",
  4078 => x"C0C0C0C099C0F880",
  4079 => x"C0C0C0C099C0F890",
  4080 => x"C0C0C0C099C080C0",
  4081 => x"C0C0C0C099C080F9",
  4082 => x"C0C0C0C099C080A4",
  4083 => x"C0C0C0C099C080B0",
  4084 => x"C0C0C0C099C08099",
  4085 => x"C0C0C0C099C08092",
  4086 => x"C0C0C0C099C08082",
  4087 => x"C0C0C0C099C080F8",
  4088 => x"C0C0C0C099C08080",
  4089 => x"C0C0C0C099C08090",
  4090 => x"C0C0C0C099C090C0",
  4091 => x"C0C0C0C099C090F9",
  4092 => x"C0C0C0C099C090A4",
  4093 => x"C0C0C0C099C090B0",
  4094 => x"C0C0C0C099C09099",
  4095 => x"C0C0C0C099C09092",
  4096 => x"C0C0C0C099C09082",
  4097 => x"C0C0C0C099C090F8",
  4098 => x"C0C0C0C099C09080",
  4099 => x"C0C0C0C099C09090",
  4100 => x"C0C0C0C099F9C0C0",
  4101 => x"C0C0C0C099F9C0F9",
  4102 => x"C0C0C0C099F9C0A4",
  4103 => x"C0C0C0C099F9C0B0",
  4104 => x"C0C0C0C099F9C099",
  4105 => x"C0C0C0C099F9C092",
  4106 => x"C0C0C0C099F9C082",
  4107 => x"C0C0C0C099F9C0F8",
  4108 => x"C0C0C0C099F9C080",
  4109 => x"C0C0C0C099F9C090",
  4110 => x"C0C0C0C099F9F9C0",
  4111 => x"C0C0C0C099F9F9F9",
  4112 => x"C0C0C0C099F9F9A4",
  4113 => x"C0C0C0C099F9F9B0",
  4114 => x"C0C0C0C099F9F999",
  4115 => x"C0C0C0C099F9F992",
  4116 => x"C0C0C0C099F9F982",
  4117 => x"C0C0C0C099F9F9F8",
  4118 => x"C0C0C0C099F9F980",
  4119 => x"C0C0C0C099F9F990",
  4120 => x"C0C0C0C099F9A4C0",
  4121 => x"C0C0C0C099F9A4F9",
  4122 => x"C0C0C0C099F9A4A4",
  4123 => x"C0C0C0C099F9A4B0",
  4124 => x"C0C0C0C099F9A499",
  4125 => x"C0C0C0C099F9A492",
  4126 => x"C0C0C0C099F9A482",
  4127 => x"C0C0C0C099F9A4F8",
  4128 => x"C0C0C0C099F9A480",
  4129 => x"C0C0C0C099F9A490",
  4130 => x"C0C0C0C099F9B0C0",
  4131 => x"C0C0C0C099F9B0F9",
  4132 => x"C0C0C0C099F9B0A4",
  4133 => x"C0C0C0C099F9B0B0",
  4134 => x"C0C0C0C099F9B099",
  4135 => x"C0C0C0C099F9B092",
  4136 => x"C0C0C0C099F9B082",
  4137 => x"C0C0C0C099F9B0F8",
  4138 => x"C0C0C0C099F9B080",
  4139 => x"C0C0C0C099F9B090",
  4140 => x"C0C0C0C099F999C0",
  4141 => x"C0C0C0C099F999F9",
  4142 => x"C0C0C0C099F999A4",
  4143 => x"C0C0C0C099F999B0",
  4144 => x"C0C0C0C099F99999",
  4145 => x"C0C0C0C099F99992",
  4146 => x"C0C0C0C099F99982",
  4147 => x"C0C0C0C099F999F8",
  4148 => x"C0C0C0C099F99980",
  4149 => x"C0C0C0C099F99990",
  4150 => x"C0C0C0C099F992C0",
  4151 => x"C0C0C0C099F992F9",
  4152 => x"C0C0C0C099F992A4",
  4153 => x"C0C0C0C099F992B0",
  4154 => x"C0C0C0C099F99299",
  4155 => x"C0C0C0C099F99292",
  4156 => x"C0C0C0C099F99282",
  4157 => x"C0C0C0C099F992F8",
  4158 => x"C0C0C0C099F99280",
  4159 => x"C0C0C0C099F99290",
  4160 => x"C0C0C0C099F982C0",
  4161 => x"C0C0C0C099F982F9",
  4162 => x"C0C0C0C099F982A4",
  4163 => x"C0C0C0C099F982B0",
  4164 => x"C0C0C0C099F98299",
  4165 => x"C0C0C0C099F98292",
  4166 => x"C0C0C0C099F98282",
  4167 => x"C0C0C0C099F982F8",
  4168 => x"C0C0C0C099F98280",
  4169 => x"C0C0C0C099F98290",
  4170 => x"C0C0C0C099F9F8C0",
  4171 => x"C0C0C0C099F9F8F9",
  4172 => x"C0C0C0C099F9F8A4",
  4173 => x"C0C0C0C099F9F8B0",
  4174 => x"C0C0C0C099F9F899",
  4175 => x"C0C0C0C099F9F892",
  4176 => x"C0C0C0C099F9F882",
  4177 => x"C0C0C0C099F9F8F8",
  4178 => x"C0C0C0C099F9F880",
  4179 => x"C0C0C0C099F9F890",
  4180 => x"C0C0C0C099F980C0",
  4181 => x"C0C0C0C099F980F9",
  4182 => x"C0C0C0C099F980A4",
  4183 => x"C0C0C0C099F980B0",
  4184 => x"C0C0C0C099F98099",
  4185 => x"C0C0C0C099F98092",
  4186 => x"C0C0C0C099F98082",
  4187 => x"C0C0C0C099F980F8",
  4188 => x"C0C0C0C099F98080",
  4189 => x"C0C0C0C099F98090",
  4190 => x"C0C0C0C099F990C0",
  4191 => x"C0C0C0C099F990F9",
  4192 => x"C0C0C0C099F990A4",
  4193 => x"C0C0C0C099F990B0",
  4194 => x"C0C0C0C099F99099",
  4195 => x"C0C0C0C099F99092",
  4196 => x"C0C0C0C099F99082",
  4197 => x"C0C0C0C099F990F8",
  4198 => x"C0C0C0C099F99080",
  4199 => x"C0C0C0C099F99090",
  4200 => x"C0C0C0C099A4C0C0",
  4201 => x"C0C0C0C099A4C0F9",
  4202 => x"C0C0C0C099A4C0A4",
  4203 => x"C0C0C0C099A4C0B0",
  4204 => x"C0C0C0C099A4C099",
  4205 => x"C0C0C0C099A4C092",
  4206 => x"C0C0C0C099A4C082",
  4207 => x"C0C0C0C099A4C0F8",
  4208 => x"C0C0C0C099A4C080",
  4209 => x"C0C0C0C099A4C090",
  4210 => x"C0C0C0C099A4F9C0",
  4211 => x"C0C0C0C099A4F9F9",
  4212 => x"C0C0C0C099A4F9A4",
  4213 => x"C0C0C0C099A4F9B0",
  4214 => x"C0C0C0C099A4F999",
  4215 => x"C0C0C0C099A4F992",
  4216 => x"C0C0C0C099A4F982",
  4217 => x"C0C0C0C099A4F9F8",
  4218 => x"C0C0C0C099A4F980",
  4219 => x"C0C0C0C099A4F990",
  4220 => x"C0C0C0C099A4A4C0",
  4221 => x"C0C0C0C099A4A4F9",
  4222 => x"C0C0C0C099A4A4A4",
  4223 => x"C0C0C0C099A4A4B0",
  4224 => x"C0C0C0C099A4A499",
  4225 => x"C0C0C0C099A4A492",
  4226 => x"C0C0C0C099A4A482",
  4227 => x"C0C0C0C099A4A4F8",
  4228 => x"C0C0C0C099A4A480",
  4229 => x"C0C0C0C099A4A490",
  4230 => x"C0C0C0C099A4B0C0",
  4231 => x"C0C0C0C099A4B0F9",
  4232 => x"C0C0C0C099A4B0A4",
  4233 => x"C0C0C0C099A4B0B0",
  4234 => x"C0C0C0C099A4B099",
  4235 => x"C0C0C0C099A4B092",
  4236 => x"C0C0C0C099A4B082",
  4237 => x"C0C0C0C099A4B0F8",
  4238 => x"C0C0C0C099A4B080",
  4239 => x"C0C0C0C099A4B090",
  4240 => x"C0C0C0C099A499C0",
  4241 => x"C0C0C0C099A499F9",
  4242 => x"C0C0C0C099A499A4",
  4243 => x"C0C0C0C099A499B0",
  4244 => x"C0C0C0C099A49999",
  4245 => x"C0C0C0C099A49992",
  4246 => x"C0C0C0C099A49982",
  4247 => x"C0C0C0C099A499F8",
  4248 => x"C0C0C0C099A49980",
  4249 => x"C0C0C0C099A49990",
  4250 => x"C0C0C0C099A492C0",
  4251 => x"C0C0C0C099A492F9",
  4252 => x"C0C0C0C099A492A4",
  4253 => x"C0C0C0C099A492B0",
  4254 => x"C0C0C0C099A49299",
  4255 => x"C0C0C0C099A49292",
  4256 => x"C0C0C0C099A49282",
  4257 => x"C0C0C0C099A492F8",
  4258 => x"C0C0C0C099A49280",
  4259 => x"C0C0C0C099A49290",
  4260 => x"C0C0C0C099A482C0",
  4261 => x"C0C0C0C099A482F9",
  4262 => x"C0C0C0C099A482A4",
  4263 => x"C0C0C0C099A482B0",
  4264 => x"C0C0C0C099A48299",
  4265 => x"C0C0C0C099A48292",
  4266 => x"C0C0C0C099A48282",
  4267 => x"C0C0C0C099A482F8",
  4268 => x"C0C0C0C099A48280",
  4269 => x"C0C0C0C099A48290",
  4270 => x"C0C0C0C099A4F8C0",
  4271 => x"C0C0C0C099A4F8F9",
  4272 => x"C0C0C0C099A4F8A4",
  4273 => x"C0C0C0C099A4F8B0",
  4274 => x"C0C0C0C099A4F899",
  4275 => x"C0C0C0C099A4F892",
  4276 => x"C0C0C0C099A4F882",
  4277 => x"C0C0C0C099A4F8F8",
  4278 => x"C0C0C0C099A4F880",
  4279 => x"C0C0C0C099A4F890",
  4280 => x"C0C0C0C099A480C0",
  4281 => x"C0C0C0C099A480F9",
  4282 => x"C0C0C0C099A480A4",
  4283 => x"C0C0C0C099A480B0",
  4284 => x"C0C0C0C099A48099",
  4285 => x"C0C0C0C099A48092",
  4286 => x"C0C0C0C099A48082",
  4287 => x"C0C0C0C099A480F8",
  4288 => x"C0C0C0C099A48080",
  4289 => x"C0C0C0C099A48090",
  4290 => x"C0C0C0C099A490C0",
  4291 => x"C0C0C0C099A490F9",
  4292 => x"C0C0C0C099A490A4",
  4293 => x"C0C0C0C099A490B0",
  4294 => x"C0C0C0C099A49099",
  4295 => x"C0C0C0C099A49092",
  4296 => x"C0C0C0C099A49082",
  4297 => x"C0C0C0C099A490F8",
  4298 => x"C0C0C0C099A49080",
  4299 => x"C0C0C0C099A49090",
  4300 => x"C0C0C0C099B0C0C0",
  4301 => x"C0C0C0C099B0C0F9",
  4302 => x"C0C0C0C099B0C0A4",
  4303 => x"C0C0C0C099B0C0B0",
  4304 => x"C0C0C0C099B0C099",
  4305 => x"C0C0C0C099B0C092",
  4306 => x"C0C0C0C099B0C082",
  4307 => x"C0C0C0C099B0C0F8",
  4308 => x"C0C0C0C099B0C080",
  4309 => x"C0C0C0C099B0C090",
  4310 => x"C0C0C0C099B0F9C0",
  4311 => x"C0C0C0C099B0F9F9",
  4312 => x"C0C0C0C099B0F9A4",
  4313 => x"C0C0C0C099B0F9B0",
  4314 => x"C0C0C0C099B0F999",
  4315 => x"C0C0C0C099B0F992",
  4316 => x"C0C0C0C099B0F982",
  4317 => x"C0C0C0C099B0F9F8",
  4318 => x"C0C0C0C099B0F980",
  4319 => x"C0C0C0C099B0F990",
  4320 => x"C0C0C0C099B0A4C0",
  4321 => x"C0C0C0C099B0A4F9",
  4322 => x"C0C0C0C099B0A4A4",
  4323 => x"C0C0C0C099B0A4B0",
  4324 => x"C0C0C0C099B0A499",
  4325 => x"C0C0C0C099B0A492",
  4326 => x"C0C0C0C099B0A482",
  4327 => x"C0C0C0C099B0A4F8",
  4328 => x"C0C0C0C099B0A480",
  4329 => x"C0C0C0C099B0A490",
  4330 => x"C0C0C0C099B0B0C0",
  4331 => x"C0C0C0C099B0B0F9",
  4332 => x"C0C0C0C099B0B0A4",
  4333 => x"C0C0C0C099B0B0B0",
  4334 => x"C0C0C0C099B0B099",
  4335 => x"C0C0C0C099B0B092",
  4336 => x"C0C0C0C099B0B082",
  4337 => x"C0C0C0C099B0B0F8",
  4338 => x"C0C0C0C099B0B080",
  4339 => x"C0C0C0C099B0B090",
  4340 => x"C0C0C0C099B099C0",
  4341 => x"C0C0C0C099B099F9",
  4342 => x"C0C0C0C099B099A4",
  4343 => x"C0C0C0C099B099B0",
  4344 => x"C0C0C0C099B09999",
  4345 => x"C0C0C0C099B09992",
  4346 => x"C0C0C0C099B09982",
  4347 => x"C0C0C0C099B099F8",
  4348 => x"C0C0C0C099B09980",
  4349 => x"C0C0C0C099B09990",
  4350 => x"C0C0C0C099B092C0",
  4351 => x"C0C0C0C099B092F9",
  4352 => x"C0C0C0C099B092A4",
  4353 => x"C0C0C0C099B092B0",
  4354 => x"C0C0C0C099B09299",
  4355 => x"C0C0C0C099B09292",
  4356 => x"C0C0C0C099B09282",
  4357 => x"C0C0C0C099B092F8",
  4358 => x"C0C0C0C099B09280",
  4359 => x"C0C0C0C099B09290",
  4360 => x"C0C0C0C099B082C0",
  4361 => x"C0C0C0C099B082F9",
  4362 => x"C0C0C0C099B082A4",
  4363 => x"C0C0C0C099B082B0",
  4364 => x"C0C0C0C099B08299",
  4365 => x"C0C0C0C099B08292",
  4366 => x"C0C0C0C099B08282",
  4367 => x"C0C0C0C099B082F8",
  4368 => x"C0C0C0C099B08280",
  4369 => x"C0C0C0C099B08290",
  4370 => x"C0C0C0C099B0F8C0",
  4371 => x"C0C0C0C099B0F8F9",
  4372 => x"C0C0C0C099B0F8A4",
  4373 => x"C0C0C0C099B0F8B0",
  4374 => x"C0C0C0C099B0F899",
  4375 => x"C0C0C0C099B0F892",
  4376 => x"C0C0C0C099B0F882",
  4377 => x"C0C0C0C099B0F8F8",
  4378 => x"C0C0C0C099B0F880",
  4379 => x"C0C0C0C099B0F890",
  4380 => x"C0C0C0C099B080C0",
  4381 => x"C0C0C0C099B080F9",
  4382 => x"C0C0C0C099B080A4",
  4383 => x"C0C0C0C099B080B0",
  4384 => x"C0C0C0C099B08099",
  4385 => x"C0C0C0C099B08092",
  4386 => x"C0C0C0C099B08082",
  4387 => x"C0C0C0C099B080F8",
  4388 => x"C0C0C0C099B08080",
  4389 => x"C0C0C0C099B08090",
  4390 => x"C0C0C0C099B090C0",
  4391 => x"C0C0C0C099B090F9",
  4392 => x"C0C0C0C099B090A4",
  4393 => x"C0C0C0C099B090B0",
  4394 => x"C0C0C0C099B09099",
  4395 => x"C0C0C0C099B09092",
  4396 => x"C0C0C0C099B09082",
  4397 => x"C0C0C0C099B090F8",
  4398 => x"C0C0C0C099B09080",
  4399 => x"C0C0C0C099B09090",
  4400 => x"C0C0C0C09999C0C0",
  4401 => x"C0C0C0C09999C0F9",
  4402 => x"C0C0C0C09999C0A4",
  4403 => x"C0C0C0C09999C0B0",
  4404 => x"C0C0C0C09999C099",
  4405 => x"C0C0C0C09999C092",
  4406 => x"C0C0C0C09999C082",
  4407 => x"C0C0C0C09999C0F8",
  4408 => x"C0C0C0C09999C080",
  4409 => x"C0C0C0C09999C090",
  4410 => x"C0C0C0C09999F9C0",
  4411 => x"C0C0C0C09999F9F9",
  4412 => x"C0C0C0C09999F9A4",
  4413 => x"C0C0C0C09999F9B0",
  4414 => x"C0C0C0C09999F999",
  4415 => x"C0C0C0C09999F992",
  4416 => x"C0C0C0C09999F982",
  4417 => x"C0C0C0C09999F9F8",
  4418 => x"C0C0C0C09999F980",
  4419 => x"C0C0C0C09999F990",
  4420 => x"C0C0C0C09999A4C0",
  4421 => x"C0C0C0C09999A4F9",
  4422 => x"C0C0C0C09999A4A4",
  4423 => x"C0C0C0C09999A4B0",
  4424 => x"C0C0C0C09999A499",
  4425 => x"C0C0C0C09999A492",
  4426 => x"C0C0C0C09999A482",
  4427 => x"C0C0C0C09999A4F8",
  4428 => x"C0C0C0C09999A480",
  4429 => x"C0C0C0C09999A490",
  4430 => x"C0C0C0C09999B0C0",
  4431 => x"C0C0C0C09999B0F9",
  4432 => x"C0C0C0C09999B0A4",
  4433 => x"C0C0C0C09999B0B0",
  4434 => x"C0C0C0C09999B099",
  4435 => x"C0C0C0C09999B092",
  4436 => x"C0C0C0C09999B082",
  4437 => x"C0C0C0C09999B0F8",
  4438 => x"C0C0C0C09999B080",
  4439 => x"C0C0C0C09999B090",
  4440 => x"C0C0C0C0999999C0",
  4441 => x"C0C0C0C0999999F9",
  4442 => x"C0C0C0C0999999A4",
  4443 => x"C0C0C0C0999999B0",
  4444 => x"C0C0C0C099999999",
  4445 => x"C0C0C0C099999992",
  4446 => x"C0C0C0C099999982",
  4447 => x"C0C0C0C0999999F8",
  4448 => x"C0C0C0C099999980",
  4449 => x"C0C0C0C099999990",
  4450 => x"C0C0C0C0999992C0",
  4451 => x"C0C0C0C0999992F9",
  4452 => x"C0C0C0C0999992A4",
  4453 => x"C0C0C0C0999992B0",
  4454 => x"C0C0C0C099999299",
  4455 => x"C0C0C0C099999292",
  4456 => x"C0C0C0C099999282",
  4457 => x"C0C0C0C0999992F8",
  4458 => x"C0C0C0C099999280",
  4459 => x"C0C0C0C099999290",
  4460 => x"C0C0C0C0999982C0",
  4461 => x"C0C0C0C0999982F9",
  4462 => x"C0C0C0C0999982A4",
  4463 => x"C0C0C0C0999982B0",
  4464 => x"C0C0C0C099998299",
  4465 => x"C0C0C0C099998292",
  4466 => x"C0C0C0C099998282",
  4467 => x"C0C0C0C0999982F8",
  4468 => x"C0C0C0C099998280",
  4469 => x"C0C0C0C099998290",
  4470 => x"C0C0C0C09999F8C0",
  4471 => x"C0C0C0C09999F8F9",
  4472 => x"C0C0C0C09999F8A4",
  4473 => x"C0C0C0C09999F8B0",
  4474 => x"C0C0C0C09999F899",
  4475 => x"C0C0C0C09999F892",
  4476 => x"C0C0C0C09999F882",
  4477 => x"C0C0C0C09999F8F8",
  4478 => x"C0C0C0C09999F880",
  4479 => x"C0C0C0C09999F890",
  4480 => x"C0C0C0C0999980C0",
  4481 => x"C0C0C0C0999980F9",
  4482 => x"C0C0C0C0999980A4",
  4483 => x"C0C0C0C0999980B0",
  4484 => x"C0C0C0C099998099",
  4485 => x"C0C0C0C099998092",
  4486 => x"C0C0C0C099998082",
  4487 => x"C0C0C0C0999980F8",
  4488 => x"C0C0C0C099998080",
  4489 => x"C0C0C0C099998090",
  4490 => x"C0C0C0C0999990C0",
  4491 => x"C0C0C0C0999990F9",
  4492 => x"C0C0C0C0999990A4",
  4493 => x"C0C0C0C0999990B0",
  4494 => x"C0C0C0C099999099",
  4495 => x"C0C0C0C099999092",
  4496 => x"C0C0C0C099999082",
  4497 => x"C0C0C0C0999990F8",
  4498 => x"C0C0C0C099999080",
  4499 => x"C0C0C0C099999090",
  4500 => x"C0C0C0C09992C0C0",
  4501 => x"C0C0C0C09992C0F9",
  4502 => x"C0C0C0C09992C0A4",
  4503 => x"C0C0C0C09992C0B0",
  4504 => x"C0C0C0C09992C099",
  4505 => x"C0C0C0C09992C092",
  4506 => x"C0C0C0C09992C082",
  4507 => x"C0C0C0C09992C0F8",
  4508 => x"C0C0C0C09992C080",
  4509 => x"C0C0C0C09992C090",
  4510 => x"C0C0C0C09992F9C0",
  4511 => x"C0C0C0C09992F9F9",
  4512 => x"C0C0C0C09992F9A4",
  4513 => x"C0C0C0C09992F9B0",
  4514 => x"C0C0C0C09992F999",
  4515 => x"C0C0C0C09992F992",
  4516 => x"C0C0C0C09992F982",
  4517 => x"C0C0C0C09992F9F8",
  4518 => x"C0C0C0C09992F980",
  4519 => x"C0C0C0C09992F990",
  4520 => x"C0C0C0C09992A4C0",
  4521 => x"C0C0C0C09992A4F9",
  4522 => x"C0C0C0C09992A4A4",
  4523 => x"C0C0C0C09992A4B0",
  4524 => x"C0C0C0C09992A499",
  4525 => x"C0C0C0C09992A492",
  4526 => x"C0C0C0C09992A482",
  4527 => x"C0C0C0C09992A4F8",
  4528 => x"C0C0C0C09992A480",
  4529 => x"C0C0C0C09992A490",
  4530 => x"C0C0C0C09992B0C0",
  4531 => x"C0C0C0C09992B0F9",
  4532 => x"C0C0C0C09992B0A4",
  4533 => x"C0C0C0C09992B0B0",
  4534 => x"C0C0C0C09992B099",
  4535 => x"C0C0C0C09992B092",
  4536 => x"C0C0C0C09992B082",
  4537 => x"C0C0C0C09992B0F8",
  4538 => x"C0C0C0C09992B080",
  4539 => x"C0C0C0C09992B090",
  4540 => x"C0C0C0C0999299C0",
  4541 => x"C0C0C0C0999299F9",
  4542 => x"C0C0C0C0999299A4",
  4543 => x"C0C0C0C0999299B0",
  4544 => x"C0C0C0C099929999",
  4545 => x"C0C0C0C099929992",
  4546 => x"C0C0C0C099929982",
  4547 => x"C0C0C0C0999299F8",
  4548 => x"C0C0C0C099929980",
  4549 => x"C0C0C0C099929990",
  4550 => x"C0C0C0C0999292C0",
  4551 => x"C0C0C0C0999292F9",
  4552 => x"C0C0C0C0999292A4",
  4553 => x"C0C0C0C0999292B0",
  4554 => x"C0C0C0C099929299",
  4555 => x"C0C0C0C099929292",
  4556 => x"C0C0C0C099929282",
  4557 => x"C0C0C0C0999292F8",
  4558 => x"C0C0C0C099929280",
  4559 => x"C0C0C0C099929290",
  4560 => x"C0C0C0C0999282C0",
  4561 => x"C0C0C0C0999282F9",
  4562 => x"C0C0C0C0999282A4",
  4563 => x"C0C0C0C0999282B0",
  4564 => x"C0C0C0C099928299",
  4565 => x"C0C0C0C099928292",
  4566 => x"C0C0C0C099928282",
  4567 => x"C0C0C0C0999282F8",
  4568 => x"C0C0C0C099928280",
  4569 => x"C0C0C0C099928290",
  4570 => x"C0C0C0C09992F8C0",
  4571 => x"C0C0C0C09992F8F9",
  4572 => x"C0C0C0C09992F8A4",
  4573 => x"C0C0C0C09992F8B0",
  4574 => x"C0C0C0C09992F899",
  4575 => x"C0C0C0C09992F892",
  4576 => x"C0C0C0C09992F882",
  4577 => x"C0C0C0C09992F8F8",
  4578 => x"C0C0C0C09992F880",
  4579 => x"C0C0C0C09992F890",
  4580 => x"C0C0C0C0999280C0",
  4581 => x"C0C0C0C0999280F9",
  4582 => x"C0C0C0C0999280A4",
  4583 => x"C0C0C0C0999280B0",
  4584 => x"C0C0C0C099928099",
  4585 => x"C0C0C0C099928092",
  4586 => x"C0C0C0C099928082",
  4587 => x"C0C0C0C0999280F8",
  4588 => x"C0C0C0C099928080",
  4589 => x"C0C0C0C099928090",
  4590 => x"C0C0C0C0999290C0",
  4591 => x"C0C0C0C0999290F9",
  4592 => x"C0C0C0C0999290A4",
  4593 => x"C0C0C0C0999290B0",
  4594 => x"C0C0C0C099929099",
  4595 => x"C0C0C0C099929092",
  4596 => x"C0C0C0C099929082",
  4597 => x"C0C0C0C0999290F8",
  4598 => x"C0C0C0C099929080",
  4599 => x"C0C0C0C099929090",
  4600 => x"C0C0C0C09982C0C0",
  4601 => x"C0C0C0C09982C0F9",
  4602 => x"C0C0C0C09982C0A4",
  4603 => x"C0C0C0C09982C0B0",
  4604 => x"C0C0C0C09982C099",
  4605 => x"C0C0C0C09982C092",
  4606 => x"C0C0C0C09982C082",
  4607 => x"C0C0C0C09982C0F8",
  4608 => x"C0C0C0C09982C080",
  4609 => x"C0C0C0C09982C090",
  4610 => x"C0C0C0C09982F9C0",
  4611 => x"C0C0C0C09982F9F9",
  4612 => x"C0C0C0C09982F9A4",
  4613 => x"C0C0C0C09982F9B0",
  4614 => x"C0C0C0C09982F999",
  4615 => x"C0C0C0C09982F992",
  4616 => x"C0C0C0C09982F982",
  4617 => x"C0C0C0C09982F9F8",
  4618 => x"C0C0C0C09982F980",
  4619 => x"C0C0C0C09982F990",
  4620 => x"C0C0C0C09982A4C0",
  4621 => x"C0C0C0C09982A4F9",
  4622 => x"C0C0C0C09982A4A4",
  4623 => x"C0C0C0C09982A4B0",
  4624 => x"C0C0C0C09982A499",
  4625 => x"C0C0C0C09982A492",
  4626 => x"C0C0C0C09982A482",
  4627 => x"C0C0C0C09982A4F8",
  4628 => x"C0C0C0C09982A480",
  4629 => x"C0C0C0C09982A490",
  4630 => x"C0C0C0C09982B0C0",
  4631 => x"C0C0C0C09982B0F9",
  4632 => x"C0C0C0C09982B0A4",
  4633 => x"C0C0C0C09982B0B0",
  4634 => x"C0C0C0C09982B099",
  4635 => x"C0C0C0C09982B092",
  4636 => x"C0C0C0C09982B082",
  4637 => x"C0C0C0C09982B0F8",
  4638 => x"C0C0C0C09982B080",
  4639 => x"C0C0C0C09982B090",
  4640 => x"C0C0C0C0998299C0",
  4641 => x"C0C0C0C0998299F9",
  4642 => x"C0C0C0C0998299A4",
  4643 => x"C0C0C0C0998299B0",
  4644 => x"C0C0C0C099829999",
  4645 => x"C0C0C0C099829992",
  4646 => x"C0C0C0C099829982",
  4647 => x"C0C0C0C0998299F8",
  4648 => x"C0C0C0C099829980",
  4649 => x"C0C0C0C099829990",
  4650 => x"C0C0C0C0998292C0",
  4651 => x"C0C0C0C0998292F9",
  4652 => x"C0C0C0C0998292A4",
  4653 => x"C0C0C0C0998292B0",
  4654 => x"C0C0C0C099829299",
  4655 => x"C0C0C0C099829292",
  4656 => x"C0C0C0C099829282",
  4657 => x"C0C0C0C0998292F8",
  4658 => x"C0C0C0C099829280",
  4659 => x"C0C0C0C099829290",
  4660 => x"C0C0C0C0998282C0",
  4661 => x"C0C0C0C0998282F9",
  4662 => x"C0C0C0C0998282A4",
  4663 => x"C0C0C0C0998282B0",
  4664 => x"C0C0C0C099828299",
  4665 => x"C0C0C0C099828292",
  4666 => x"C0C0C0C099828282",
  4667 => x"C0C0C0C0998282F8",
  4668 => x"C0C0C0C099828280",
  4669 => x"C0C0C0C099828290",
  4670 => x"C0C0C0C09982F8C0",
  4671 => x"C0C0C0C09982F8F9",
  4672 => x"C0C0C0C09982F8A4",
  4673 => x"C0C0C0C09982F8B0",
  4674 => x"C0C0C0C09982F899",
  4675 => x"C0C0C0C09982F892",
  4676 => x"C0C0C0C09982F882",
  4677 => x"C0C0C0C09982F8F8",
  4678 => x"C0C0C0C09982F880",
  4679 => x"C0C0C0C09982F890",
  4680 => x"C0C0C0C0998280C0",
  4681 => x"C0C0C0C0998280F9",
  4682 => x"C0C0C0C0998280A4",
  4683 => x"C0C0C0C0998280B0",
  4684 => x"C0C0C0C099828099",
  4685 => x"C0C0C0C099828092",
  4686 => x"C0C0C0C099828082",
  4687 => x"C0C0C0C0998280F8",
  4688 => x"C0C0C0C099828080",
  4689 => x"C0C0C0C099828090",
  4690 => x"C0C0C0C0998290C0",
  4691 => x"C0C0C0C0998290F9",
  4692 => x"C0C0C0C0998290A4",
  4693 => x"C0C0C0C0998290B0",
  4694 => x"C0C0C0C099829099",
  4695 => x"C0C0C0C099829092",
  4696 => x"C0C0C0C099829082",
  4697 => x"C0C0C0C0998290F8",
  4698 => x"C0C0C0C099829080",
  4699 => x"C0C0C0C099829090",
  4700 => x"C0C0C0C099F8C0C0",
  4701 => x"C0C0C0C099F8C0F9",
  4702 => x"C0C0C0C099F8C0A4",
  4703 => x"C0C0C0C099F8C0B0",
  4704 => x"C0C0C0C099F8C099",
  4705 => x"C0C0C0C099F8C092",
  4706 => x"C0C0C0C099F8C082",
  4707 => x"C0C0C0C099F8C0F8",
  4708 => x"C0C0C0C099F8C080",
  4709 => x"C0C0C0C099F8C090",
  4710 => x"C0C0C0C099F8F9C0",
  4711 => x"C0C0C0C099F8F9F9",
  4712 => x"C0C0C0C099F8F9A4",
  4713 => x"C0C0C0C099F8F9B0",
  4714 => x"C0C0C0C099F8F999",
  4715 => x"C0C0C0C099F8F992",
  4716 => x"C0C0C0C099F8F982",
  4717 => x"C0C0C0C099F8F9F8",
  4718 => x"C0C0C0C099F8F980",
  4719 => x"C0C0C0C099F8F990",
  4720 => x"C0C0C0C099F8A4C0",
  4721 => x"C0C0C0C099F8A4F9",
  4722 => x"C0C0C0C099F8A4A4",
  4723 => x"C0C0C0C099F8A4B0",
  4724 => x"C0C0C0C099F8A499",
  4725 => x"C0C0C0C099F8A492",
  4726 => x"C0C0C0C099F8A482",
  4727 => x"C0C0C0C099F8A4F8",
  4728 => x"C0C0C0C099F8A480",
  4729 => x"C0C0C0C099F8A490",
  4730 => x"C0C0C0C099F8B0C0",
  4731 => x"C0C0C0C099F8B0F9",
  4732 => x"C0C0C0C099F8B0A4",
  4733 => x"C0C0C0C099F8B0B0",
  4734 => x"C0C0C0C099F8B099",
  4735 => x"C0C0C0C099F8B092",
  4736 => x"C0C0C0C099F8B082",
  4737 => x"C0C0C0C099F8B0F8",
  4738 => x"C0C0C0C099F8B080",
  4739 => x"C0C0C0C099F8B090",
  4740 => x"C0C0C0C099F899C0",
  4741 => x"C0C0C0C099F899F9",
  4742 => x"C0C0C0C099F899A4",
  4743 => x"C0C0C0C099F899B0",
  4744 => x"C0C0C0C099F89999",
  4745 => x"C0C0C0C099F89992",
  4746 => x"C0C0C0C099F89982",
  4747 => x"C0C0C0C099F899F8",
  4748 => x"C0C0C0C099F89980",
  4749 => x"C0C0C0C099F89990",
  4750 => x"C0C0C0C099F892C0",
  4751 => x"C0C0C0C099F892F9",
  4752 => x"C0C0C0C099F892A4",
  4753 => x"C0C0C0C099F892B0",
  4754 => x"C0C0C0C099F89299",
  4755 => x"C0C0C0C099F89292",
  4756 => x"C0C0C0C099F89282",
  4757 => x"C0C0C0C099F892F8",
  4758 => x"C0C0C0C099F89280",
  4759 => x"C0C0C0C099F89290",
  4760 => x"C0C0C0C099F882C0",
  4761 => x"C0C0C0C099F882F9",
  4762 => x"C0C0C0C099F882A4",
  4763 => x"C0C0C0C099F882B0",
  4764 => x"C0C0C0C099F88299",
  4765 => x"C0C0C0C099F88292",
  4766 => x"C0C0C0C099F88282",
  4767 => x"C0C0C0C099F882F8",
  4768 => x"C0C0C0C099F88280",
  4769 => x"C0C0C0C099F88290",
  4770 => x"C0C0C0C099F8F8C0",
  4771 => x"C0C0C0C099F8F8F9",
  4772 => x"C0C0C0C099F8F8A4",
  4773 => x"C0C0C0C099F8F8B0",
  4774 => x"C0C0C0C099F8F899",
  4775 => x"C0C0C0C099F8F892",
  4776 => x"C0C0C0C099F8F882",
  4777 => x"C0C0C0C099F8F8F8",
  4778 => x"C0C0C0C099F8F880",
  4779 => x"C0C0C0C099F8F890",
  4780 => x"C0C0C0C099F880C0",
  4781 => x"C0C0C0C099F880F9",
  4782 => x"C0C0C0C099F880A4",
  4783 => x"C0C0C0C099F880B0",
  4784 => x"C0C0C0C099F88099",
  4785 => x"C0C0C0C099F88092",
  4786 => x"C0C0C0C099F88082",
  4787 => x"C0C0C0C099F880F8",
  4788 => x"C0C0C0C099F88080",
  4789 => x"C0C0C0C099F88090",
  4790 => x"C0C0C0C099F890C0",
  4791 => x"C0C0C0C099F890F9",
  4792 => x"C0C0C0C099F890A4",
  4793 => x"C0C0C0C099F890B0",
  4794 => x"C0C0C0C099F89099",
  4795 => x"C0C0C0C099F89092",
  4796 => x"C0C0C0C099F89082",
  4797 => x"C0C0C0C099F890F8",
  4798 => x"C0C0C0C099F89080",
  4799 => x"C0C0C0C099F89090",
  4800 => x"C0C0C0C09980C0C0",
  4801 => x"C0C0C0C09980C0F9",
  4802 => x"C0C0C0C09980C0A4",
  4803 => x"C0C0C0C09980C0B0",
  4804 => x"C0C0C0C09980C099",
  4805 => x"C0C0C0C09980C092",
  4806 => x"C0C0C0C09980C082",
  4807 => x"C0C0C0C09980C0F8",
  4808 => x"C0C0C0C09980C080",
  4809 => x"C0C0C0C09980C090",
  4810 => x"C0C0C0C09980F9C0",
  4811 => x"C0C0C0C09980F9F9",
  4812 => x"C0C0C0C09980F9A4",
  4813 => x"C0C0C0C09980F9B0",
  4814 => x"C0C0C0C09980F999",
  4815 => x"C0C0C0C09980F992",
  4816 => x"C0C0C0C09980F982",
  4817 => x"C0C0C0C09980F9F8",
  4818 => x"C0C0C0C09980F980",
  4819 => x"C0C0C0C09980F990",
  4820 => x"C0C0C0C09980A4C0",
  4821 => x"C0C0C0C09980A4F9",
  4822 => x"C0C0C0C09980A4A4",
  4823 => x"C0C0C0C09980A4B0",
  4824 => x"C0C0C0C09980A499",
  4825 => x"C0C0C0C09980A492",
  4826 => x"C0C0C0C09980A482",
  4827 => x"C0C0C0C09980A4F8",
  4828 => x"C0C0C0C09980A480",
  4829 => x"C0C0C0C09980A490",
  4830 => x"C0C0C0C09980B0C0",
  4831 => x"C0C0C0C09980B0F9",
  4832 => x"C0C0C0C09980B0A4",
  4833 => x"C0C0C0C09980B0B0",
  4834 => x"C0C0C0C09980B099",
  4835 => x"C0C0C0C09980B092",
  4836 => x"C0C0C0C09980B082",
  4837 => x"C0C0C0C09980B0F8",
  4838 => x"C0C0C0C09980B080",
  4839 => x"C0C0C0C09980B090",
  4840 => x"C0C0C0C0998099C0",
  4841 => x"C0C0C0C0998099F9",
  4842 => x"C0C0C0C0998099A4",
  4843 => x"C0C0C0C0998099B0",
  4844 => x"C0C0C0C099809999",
  4845 => x"C0C0C0C099809992",
  4846 => x"C0C0C0C099809982",
  4847 => x"C0C0C0C0998099F8",
  4848 => x"C0C0C0C099809980",
  4849 => x"C0C0C0C099809990",
  4850 => x"C0C0C0C0998092C0",
  4851 => x"C0C0C0C0998092F9",
  4852 => x"C0C0C0C0998092A4",
  4853 => x"C0C0C0C0998092B0",
  4854 => x"C0C0C0C099809299",
  4855 => x"C0C0C0C099809292",
  4856 => x"C0C0C0C099809282",
  4857 => x"C0C0C0C0998092F8",
  4858 => x"C0C0C0C099809280",
  4859 => x"C0C0C0C099809290",
  4860 => x"C0C0C0C0998082C0",
  4861 => x"C0C0C0C0998082F9",
  4862 => x"C0C0C0C0998082A4",
  4863 => x"C0C0C0C0998082B0",
  4864 => x"C0C0C0C099808299",
  4865 => x"C0C0C0C099808292",
  4866 => x"C0C0C0C099808282",
  4867 => x"C0C0C0C0998082F8",
  4868 => x"C0C0C0C099808280",
  4869 => x"C0C0C0C099808290",
  4870 => x"C0C0C0C09980F8C0",
  4871 => x"C0C0C0C09980F8F9",
  4872 => x"C0C0C0C09980F8A4",
  4873 => x"C0C0C0C09980F8B0",
  4874 => x"C0C0C0C09980F899",
  4875 => x"C0C0C0C09980F892",
  4876 => x"C0C0C0C09980F882",
  4877 => x"C0C0C0C09980F8F8",
  4878 => x"C0C0C0C09980F880",
  4879 => x"C0C0C0C09980F890",
  4880 => x"C0C0C0C0998080C0",
  4881 => x"C0C0C0C0998080F9",
  4882 => x"C0C0C0C0998080A4",
  4883 => x"C0C0C0C0998080B0",
  4884 => x"C0C0C0C099808099",
  4885 => x"C0C0C0C099808092",
  4886 => x"C0C0C0C099808082",
  4887 => x"C0C0C0C0998080F8",
  4888 => x"C0C0C0C099808080",
  4889 => x"C0C0C0C099808090",
  4890 => x"C0C0C0C0998090C0",
  4891 => x"C0C0C0C0998090F9",
  4892 => x"C0C0C0C0998090A4",
  4893 => x"C0C0C0C0998090B0",
  4894 => x"C0C0C0C099809099",
  4895 => x"C0C0C0C099809092",
  4896 => x"C0C0C0C099809082",
  4897 => x"C0C0C0C0998090F8",
  4898 => x"C0C0C0C099809080",
  4899 => x"C0C0C0C099809090",
  4900 => x"C0C0C0C09990C0C0",
  4901 => x"C0C0C0C09990C0F9",
  4902 => x"C0C0C0C09990C0A4",
  4903 => x"C0C0C0C09990C0B0",
  4904 => x"C0C0C0C09990C099",
  4905 => x"C0C0C0C09990C092",
  4906 => x"C0C0C0C09990C082",
  4907 => x"C0C0C0C09990C0F8",
  4908 => x"C0C0C0C09990C080",
  4909 => x"C0C0C0C09990C090",
  4910 => x"C0C0C0C09990F9C0",
  4911 => x"C0C0C0C09990F9F9",
  4912 => x"C0C0C0C09990F9A4",
  4913 => x"C0C0C0C09990F9B0",
  4914 => x"C0C0C0C09990F999",
  4915 => x"C0C0C0C09990F992",
  4916 => x"C0C0C0C09990F982",
  4917 => x"C0C0C0C09990F9F8",
  4918 => x"C0C0C0C09990F980",
  4919 => x"C0C0C0C09990F990",
  4920 => x"C0C0C0C09990A4C0",
  4921 => x"C0C0C0C09990A4F9",
  4922 => x"C0C0C0C09990A4A4",
  4923 => x"C0C0C0C09990A4B0",
  4924 => x"C0C0C0C09990A499",
  4925 => x"C0C0C0C09990A492",
  4926 => x"C0C0C0C09990A482",
  4927 => x"C0C0C0C09990A4F8",
  4928 => x"C0C0C0C09990A480",
  4929 => x"C0C0C0C09990A490",
  4930 => x"C0C0C0C09990B0C0",
  4931 => x"C0C0C0C09990B0F9",
  4932 => x"C0C0C0C09990B0A4",
  4933 => x"C0C0C0C09990B0B0",
  4934 => x"C0C0C0C09990B099",
  4935 => x"C0C0C0C09990B092",
  4936 => x"C0C0C0C09990B082",
  4937 => x"C0C0C0C09990B0F8",
  4938 => x"C0C0C0C09990B080",
  4939 => x"C0C0C0C09990B090",
  4940 => x"C0C0C0C0999099C0",
  4941 => x"C0C0C0C0999099F9",
  4942 => x"C0C0C0C0999099A4",
  4943 => x"C0C0C0C0999099B0",
  4944 => x"C0C0C0C099909999",
  4945 => x"C0C0C0C099909992",
  4946 => x"C0C0C0C099909982",
  4947 => x"C0C0C0C0999099F8",
  4948 => x"C0C0C0C099909980",
  4949 => x"C0C0C0C099909990",
  4950 => x"C0C0C0C0999092C0",
  4951 => x"C0C0C0C0999092F9",
  4952 => x"C0C0C0C0999092A4",
  4953 => x"C0C0C0C0999092B0",
  4954 => x"C0C0C0C099909299",
  4955 => x"C0C0C0C099909292",
  4956 => x"C0C0C0C099909282",
  4957 => x"C0C0C0C0999092F8",
  4958 => x"C0C0C0C099909280",
  4959 => x"C0C0C0C099909290",
  4960 => x"C0C0C0C0999082C0",
  4961 => x"C0C0C0C0999082F9",
  4962 => x"C0C0C0C0999082A4",
  4963 => x"C0C0C0C0999082B0",
  4964 => x"C0C0C0C099908299",
  4965 => x"C0C0C0C099908292",
  4966 => x"C0C0C0C099908282",
  4967 => x"C0C0C0C0999082F8",
  4968 => x"C0C0C0C099908280",
  4969 => x"C0C0C0C099908290",
  4970 => x"C0C0C0C09990F8C0",
  4971 => x"C0C0C0C09990F8F9",
  4972 => x"C0C0C0C09990F8A4",
  4973 => x"C0C0C0C09990F8B0",
  4974 => x"C0C0C0C09990F899",
  4975 => x"C0C0C0C09990F892",
  4976 => x"C0C0C0C09990F882",
  4977 => x"C0C0C0C09990F8F8",
  4978 => x"C0C0C0C09990F880",
  4979 => x"C0C0C0C09990F890",
  4980 => x"C0C0C0C0999080C0",
  4981 => x"C0C0C0C0999080F9",
  4982 => x"C0C0C0C0999080A4",
  4983 => x"C0C0C0C0999080B0",
  4984 => x"C0C0C0C099908099",
  4985 => x"C0C0C0C099908092",
  4986 => x"C0C0C0C099908082",
  4987 => x"C0C0C0C0999080F8",
  4988 => x"C0C0C0C099908080",
  4989 => x"C0C0C0C099908090",
  4990 => x"C0C0C0C0999090C0",
  4991 => x"C0C0C0C0999090F9",
  4992 => x"C0C0C0C0999090A4",
  4993 => x"C0C0C0C0999090B0",
  4994 => x"C0C0C0C099909099",
  4995 => x"C0C0C0C099909092",
  4996 => x"C0C0C0C099909082",
  4997 => x"C0C0C0C0999090F8",
  4998 => x"C0C0C0C099909080",
  4999 => x"C0C0C0C099909090",
  5000 => x"C0C0C0C092C0C0C0",
  5001 => x"C0C0C0C092C0C0F9",
  5002 => x"C0C0C0C092C0C0A4",
  5003 => x"C0C0C0C092C0C0B0",
  5004 => x"C0C0C0C092C0C099",
  5005 => x"C0C0C0C092C0C092",
  5006 => x"C0C0C0C092C0C082",
  5007 => x"C0C0C0C092C0C0F8",
  5008 => x"C0C0C0C092C0C080",
  5009 => x"C0C0C0C092C0C090",
  5010 => x"C0C0C0C092C0F9C0",
  5011 => x"C0C0C0C092C0F9F9",
  5012 => x"C0C0C0C092C0F9A4",
  5013 => x"C0C0C0C092C0F9B0",
  5014 => x"C0C0C0C092C0F999",
  5015 => x"C0C0C0C092C0F992",
  5016 => x"C0C0C0C092C0F982",
  5017 => x"C0C0C0C092C0F9F8",
  5018 => x"C0C0C0C092C0F980",
  5019 => x"C0C0C0C092C0F990",
  5020 => x"C0C0C0C092C0A4C0",
  5021 => x"C0C0C0C092C0A4F9",
  5022 => x"C0C0C0C092C0A4A4",
  5023 => x"C0C0C0C092C0A4B0",
  5024 => x"C0C0C0C092C0A499",
  5025 => x"C0C0C0C092C0A492",
  5026 => x"C0C0C0C092C0A482",
  5027 => x"C0C0C0C092C0A4F8",
  5028 => x"C0C0C0C092C0A480",
  5029 => x"C0C0C0C092C0A490",
  5030 => x"C0C0C0C092C0B0C0",
  5031 => x"C0C0C0C092C0B0F9",
  5032 => x"C0C0C0C092C0B0A4",
  5033 => x"C0C0C0C092C0B0B0",
  5034 => x"C0C0C0C092C0B099",
  5035 => x"C0C0C0C092C0B092",
  5036 => x"C0C0C0C092C0B082",
  5037 => x"C0C0C0C092C0B0F8",
  5038 => x"C0C0C0C092C0B080",
  5039 => x"C0C0C0C092C0B090",
  5040 => x"C0C0C0C092C099C0",
  5041 => x"C0C0C0C092C099F9",
  5042 => x"C0C0C0C092C099A4",
  5043 => x"C0C0C0C092C099B0",
  5044 => x"C0C0C0C092C09999",
  5045 => x"C0C0C0C092C09992",
  5046 => x"C0C0C0C092C09982",
  5047 => x"C0C0C0C092C099F8",
  5048 => x"C0C0C0C092C09980",
  5049 => x"C0C0C0C092C09990",
  5050 => x"C0C0C0C092C092C0",
  5051 => x"C0C0C0C092C092F9",
  5052 => x"C0C0C0C092C092A4",
  5053 => x"C0C0C0C092C092B0",
  5054 => x"C0C0C0C092C09299",
  5055 => x"C0C0C0C092C09292",
  5056 => x"C0C0C0C092C09282",
  5057 => x"C0C0C0C092C092F8",
  5058 => x"C0C0C0C092C09280",
  5059 => x"C0C0C0C092C09290",
  5060 => x"C0C0C0C092C082C0",
  5061 => x"C0C0C0C092C082F9",
  5062 => x"C0C0C0C092C082A4",
  5063 => x"C0C0C0C092C082B0",
  5064 => x"C0C0C0C092C08299",
  5065 => x"C0C0C0C092C08292",
  5066 => x"C0C0C0C092C08282",
  5067 => x"C0C0C0C092C082F8",
  5068 => x"C0C0C0C092C08280",
  5069 => x"C0C0C0C092C08290",
  5070 => x"C0C0C0C092C0F8C0",
  5071 => x"C0C0C0C092C0F8F9",
  5072 => x"C0C0C0C092C0F8A4",
  5073 => x"C0C0C0C092C0F8B0",
  5074 => x"C0C0C0C092C0F899",
  5075 => x"C0C0C0C092C0F892",
  5076 => x"C0C0C0C092C0F882",
  5077 => x"C0C0C0C092C0F8F8",
  5078 => x"C0C0C0C092C0F880",
  5079 => x"C0C0C0C092C0F890",
  5080 => x"C0C0C0C092C080C0",
  5081 => x"C0C0C0C092C080F9",
  5082 => x"C0C0C0C092C080A4",
  5083 => x"C0C0C0C092C080B0",
  5084 => x"C0C0C0C092C08099",
  5085 => x"C0C0C0C092C08092",
  5086 => x"C0C0C0C092C08082",
  5087 => x"C0C0C0C092C080F8",
  5088 => x"C0C0C0C092C08080",
  5089 => x"C0C0C0C092C08090",
  5090 => x"C0C0C0C092C090C0",
  5091 => x"C0C0C0C092C090F9",
  5092 => x"C0C0C0C092C090A4",
  5093 => x"C0C0C0C092C090B0",
  5094 => x"C0C0C0C092C09099",
  5095 => x"C0C0C0C092C09092",
  5096 => x"C0C0C0C092C09082",
  5097 => x"C0C0C0C092C090F8",
  5098 => x"C0C0C0C092C09080",
  5099 => x"C0C0C0C092C09090",
  5100 => x"C0C0C0C092F9C0C0",
  5101 => x"C0C0C0C092F9C0F9",
  5102 => x"C0C0C0C092F9C0A4",
  5103 => x"C0C0C0C092F9C0B0",
  5104 => x"C0C0C0C092F9C099",
  5105 => x"C0C0C0C092F9C092",
  5106 => x"C0C0C0C092F9C082",
  5107 => x"C0C0C0C092F9C0F8",
  5108 => x"C0C0C0C092F9C080",
  5109 => x"C0C0C0C092F9C090",
  5110 => x"C0C0C0C092F9F9C0",
  5111 => x"C0C0C0C092F9F9F9",
  5112 => x"C0C0C0C092F9F9A4",
  5113 => x"C0C0C0C092F9F9B0",
  5114 => x"C0C0C0C092F9F999",
  5115 => x"C0C0C0C092F9F992",
  5116 => x"C0C0C0C092F9F982",
  5117 => x"C0C0C0C092F9F9F8",
  5118 => x"C0C0C0C092F9F980",
  5119 => x"C0C0C0C092F9F990",
  5120 => x"C0C0C0C092F9A4C0",
  5121 => x"C0C0C0C092F9A4F9",
  5122 => x"C0C0C0C092F9A4A4",
  5123 => x"C0C0C0C092F9A4B0",
  5124 => x"C0C0C0C092F9A499",
  5125 => x"C0C0C0C092F9A492",
  5126 => x"C0C0C0C092F9A482",
  5127 => x"C0C0C0C092F9A4F8",
  5128 => x"C0C0C0C092F9A480",
  5129 => x"C0C0C0C092F9A490",
  5130 => x"C0C0C0C092F9B0C0",
  5131 => x"C0C0C0C092F9B0F9",
  5132 => x"C0C0C0C092F9B0A4",
  5133 => x"C0C0C0C092F9B0B0",
  5134 => x"C0C0C0C092F9B099",
  5135 => x"C0C0C0C092F9B092",
  5136 => x"C0C0C0C092F9B082",
  5137 => x"C0C0C0C092F9B0F8",
  5138 => x"C0C0C0C092F9B080",
  5139 => x"C0C0C0C092F9B090",
  5140 => x"C0C0C0C092F999C0",
  5141 => x"C0C0C0C092F999F9",
  5142 => x"C0C0C0C092F999A4",
  5143 => x"C0C0C0C092F999B0",
  5144 => x"C0C0C0C092F99999",
  5145 => x"C0C0C0C092F99992",
  5146 => x"C0C0C0C092F99982",
  5147 => x"C0C0C0C092F999F8",
  5148 => x"C0C0C0C092F99980",
  5149 => x"C0C0C0C092F99990",
  5150 => x"C0C0C0C092F992C0",
  5151 => x"C0C0C0C092F992F9",
  5152 => x"C0C0C0C092F992A4",
  5153 => x"C0C0C0C092F992B0",
  5154 => x"C0C0C0C092F99299",
  5155 => x"C0C0C0C092F99292",
  5156 => x"C0C0C0C092F99282",
  5157 => x"C0C0C0C092F992F8",
  5158 => x"C0C0C0C092F99280",
  5159 => x"C0C0C0C092F99290",
  5160 => x"C0C0C0C092F982C0",
  5161 => x"C0C0C0C092F982F9",
  5162 => x"C0C0C0C092F982A4",
  5163 => x"C0C0C0C092F982B0",
  5164 => x"C0C0C0C092F98299",
  5165 => x"C0C0C0C092F98292",
  5166 => x"C0C0C0C092F98282",
  5167 => x"C0C0C0C092F982F8",
  5168 => x"C0C0C0C092F98280",
  5169 => x"C0C0C0C092F98290",
  5170 => x"C0C0C0C092F9F8C0",
  5171 => x"C0C0C0C092F9F8F9",
  5172 => x"C0C0C0C092F9F8A4",
  5173 => x"C0C0C0C092F9F8B0",
  5174 => x"C0C0C0C092F9F899",
  5175 => x"C0C0C0C092F9F892",
  5176 => x"C0C0C0C092F9F882",
  5177 => x"C0C0C0C092F9F8F8",
  5178 => x"C0C0C0C092F9F880",
  5179 => x"C0C0C0C092F9F890",
  5180 => x"C0C0C0C092F980C0",
  5181 => x"C0C0C0C092F980F9",
  5182 => x"C0C0C0C092F980A4",
  5183 => x"C0C0C0C092F980B0",
  5184 => x"C0C0C0C092F98099",
  5185 => x"C0C0C0C092F98092",
  5186 => x"C0C0C0C092F98082",
  5187 => x"C0C0C0C092F980F8",
  5188 => x"C0C0C0C092F98080",
  5189 => x"C0C0C0C092F98090",
  5190 => x"C0C0C0C092F990C0",
  5191 => x"C0C0C0C092F990F9",
  5192 => x"C0C0C0C092F990A4",
  5193 => x"C0C0C0C092F990B0",
  5194 => x"C0C0C0C092F99099",
  5195 => x"C0C0C0C092F99092",
  5196 => x"C0C0C0C092F99082",
  5197 => x"C0C0C0C092F990F8",
  5198 => x"C0C0C0C092F99080",
  5199 => x"C0C0C0C092F99090",
  5200 => x"C0C0C0C092A4C0C0",
  5201 => x"C0C0C0C092A4C0F9",
  5202 => x"C0C0C0C092A4C0A4",
  5203 => x"C0C0C0C092A4C0B0",
  5204 => x"C0C0C0C092A4C099",
  5205 => x"C0C0C0C092A4C092",
  5206 => x"C0C0C0C092A4C082",
  5207 => x"C0C0C0C092A4C0F8",
  5208 => x"C0C0C0C092A4C080",
  5209 => x"C0C0C0C092A4C090",
  5210 => x"C0C0C0C092A4F9C0",
  5211 => x"C0C0C0C092A4F9F9",
  5212 => x"C0C0C0C092A4F9A4",
  5213 => x"C0C0C0C092A4F9B0",
  5214 => x"C0C0C0C092A4F999",
  5215 => x"C0C0C0C092A4F992",
  5216 => x"C0C0C0C092A4F982",
  5217 => x"C0C0C0C092A4F9F8",
  5218 => x"C0C0C0C092A4F980",
  5219 => x"C0C0C0C092A4F990",
  5220 => x"C0C0C0C092A4A4C0",
  5221 => x"C0C0C0C092A4A4F9",
  5222 => x"C0C0C0C092A4A4A4",
  5223 => x"C0C0C0C092A4A4B0",
  5224 => x"C0C0C0C092A4A499",
  5225 => x"C0C0C0C092A4A492",
  5226 => x"C0C0C0C092A4A482",
  5227 => x"C0C0C0C092A4A4F8",
  5228 => x"C0C0C0C092A4A480",
  5229 => x"C0C0C0C092A4A490",
  5230 => x"C0C0C0C092A4B0C0",
  5231 => x"C0C0C0C092A4B0F9",
  5232 => x"C0C0C0C092A4B0A4",
  5233 => x"C0C0C0C092A4B0B0",
  5234 => x"C0C0C0C092A4B099",
  5235 => x"C0C0C0C092A4B092",
  5236 => x"C0C0C0C092A4B082",
  5237 => x"C0C0C0C092A4B0F8",
  5238 => x"C0C0C0C092A4B080",
  5239 => x"C0C0C0C092A4B090",
  5240 => x"C0C0C0C092A499C0",
  5241 => x"C0C0C0C092A499F9",
  5242 => x"C0C0C0C092A499A4",
  5243 => x"C0C0C0C092A499B0",
  5244 => x"C0C0C0C092A49999",
  5245 => x"C0C0C0C092A49992",
  5246 => x"C0C0C0C092A49982",
  5247 => x"C0C0C0C092A499F8",
  5248 => x"C0C0C0C092A49980",
  5249 => x"C0C0C0C092A49990",
  5250 => x"C0C0C0C092A492C0",
  5251 => x"C0C0C0C092A492F9",
  5252 => x"C0C0C0C092A492A4",
  5253 => x"C0C0C0C092A492B0",
  5254 => x"C0C0C0C092A49299",
  5255 => x"C0C0C0C092A49292",
  5256 => x"C0C0C0C092A49282",
  5257 => x"C0C0C0C092A492F8",
  5258 => x"C0C0C0C092A49280",
  5259 => x"C0C0C0C092A49290",
  5260 => x"C0C0C0C092A482C0",
  5261 => x"C0C0C0C092A482F9",
  5262 => x"C0C0C0C092A482A4",
  5263 => x"C0C0C0C092A482B0",
  5264 => x"C0C0C0C092A48299",
  5265 => x"C0C0C0C092A48292",
  5266 => x"C0C0C0C092A48282",
  5267 => x"C0C0C0C092A482F8",
  5268 => x"C0C0C0C092A48280",
  5269 => x"C0C0C0C092A48290",
  5270 => x"C0C0C0C092A4F8C0",
  5271 => x"C0C0C0C092A4F8F9",
  5272 => x"C0C0C0C092A4F8A4",
  5273 => x"C0C0C0C092A4F8B0",
  5274 => x"C0C0C0C092A4F899",
  5275 => x"C0C0C0C092A4F892",
  5276 => x"C0C0C0C092A4F882",
  5277 => x"C0C0C0C092A4F8F8",
  5278 => x"C0C0C0C092A4F880",
  5279 => x"C0C0C0C092A4F890",
  5280 => x"C0C0C0C092A480C0",
  5281 => x"C0C0C0C092A480F9",
  5282 => x"C0C0C0C092A480A4",
  5283 => x"C0C0C0C092A480B0",
  5284 => x"C0C0C0C092A48099",
  5285 => x"C0C0C0C092A48092",
  5286 => x"C0C0C0C092A48082",
  5287 => x"C0C0C0C092A480F8",
  5288 => x"C0C0C0C092A48080",
  5289 => x"C0C0C0C092A48090",
  5290 => x"C0C0C0C092A490C0",
  5291 => x"C0C0C0C092A490F9",
  5292 => x"C0C0C0C092A490A4",
  5293 => x"C0C0C0C092A490B0",
  5294 => x"C0C0C0C092A49099",
  5295 => x"C0C0C0C092A49092",
  5296 => x"C0C0C0C092A49082",
  5297 => x"C0C0C0C092A490F8",
  5298 => x"C0C0C0C092A49080",
  5299 => x"C0C0C0C092A49090",
  5300 => x"C0C0C0C092B0C0C0",
  5301 => x"C0C0C0C092B0C0F9",
  5302 => x"C0C0C0C092B0C0A4",
  5303 => x"C0C0C0C092B0C0B0",
  5304 => x"C0C0C0C092B0C099",
  5305 => x"C0C0C0C092B0C092",
  5306 => x"C0C0C0C092B0C082",
  5307 => x"C0C0C0C092B0C0F8",
  5308 => x"C0C0C0C092B0C080",
  5309 => x"C0C0C0C092B0C090",
  5310 => x"C0C0C0C092B0F9C0",
  5311 => x"C0C0C0C092B0F9F9",
  5312 => x"C0C0C0C092B0F9A4",
  5313 => x"C0C0C0C092B0F9B0",
  5314 => x"C0C0C0C092B0F999",
  5315 => x"C0C0C0C092B0F992",
  5316 => x"C0C0C0C092B0F982",
  5317 => x"C0C0C0C092B0F9F8",
  5318 => x"C0C0C0C092B0F980",
  5319 => x"C0C0C0C092B0F990",
  5320 => x"C0C0C0C092B0A4C0",
  5321 => x"C0C0C0C092B0A4F9",
  5322 => x"C0C0C0C092B0A4A4",
  5323 => x"C0C0C0C092B0A4B0",
  5324 => x"C0C0C0C092B0A499",
  5325 => x"C0C0C0C092B0A492",
  5326 => x"C0C0C0C092B0A482",
  5327 => x"C0C0C0C092B0A4F8",
  5328 => x"C0C0C0C092B0A480",
  5329 => x"C0C0C0C092B0A490",
  5330 => x"C0C0C0C092B0B0C0",
  5331 => x"C0C0C0C092B0B0F9",
  5332 => x"C0C0C0C092B0B0A4",
  5333 => x"C0C0C0C092B0B0B0",
  5334 => x"C0C0C0C092B0B099",
  5335 => x"C0C0C0C092B0B092",
  5336 => x"C0C0C0C092B0B082",
  5337 => x"C0C0C0C092B0B0F8",
  5338 => x"C0C0C0C092B0B080",
  5339 => x"C0C0C0C092B0B090",
  5340 => x"C0C0C0C092B099C0",
  5341 => x"C0C0C0C092B099F9",
  5342 => x"C0C0C0C092B099A4",
  5343 => x"C0C0C0C092B099B0",
  5344 => x"C0C0C0C092B09999",
  5345 => x"C0C0C0C092B09992",
  5346 => x"C0C0C0C092B09982",
  5347 => x"C0C0C0C092B099F8",
  5348 => x"C0C0C0C092B09980",
  5349 => x"C0C0C0C092B09990",
  5350 => x"C0C0C0C092B092C0",
  5351 => x"C0C0C0C092B092F9",
  5352 => x"C0C0C0C092B092A4",
  5353 => x"C0C0C0C092B092B0",
  5354 => x"C0C0C0C092B09299",
  5355 => x"C0C0C0C092B09292",
  5356 => x"C0C0C0C092B09282",
  5357 => x"C0C0C0C092B092F8",
  5358 => x"C0C0C0C092B09280",
  5359 => x"C0C0C0C092B09290",
  5360 => x"C0C0C0C092B082C0",
  5361 => x"C0C0C0C092B082F9",
  5362 => x"C0C0C0C092B082A4",
  5363 => x"C0C0C0C092B082B0",
  5364 => x"C0C0C0C092B08299",
  5365 => x"C0C0C0C092B08292",
  5366 => x"C0C0C0C092B08282",
  5367 => x"C0C0C0C092B082F8",
  5368 => x"C0C0C0C092B08280",
  5369 => x"C0C0C0C092B08290",
  5370 => x"C0C0C0C092B0F8C0",
  5371 => x"C0C0C0C092B0F8F9",
  5372 => x"C0C0C0C092B0F8A4",
  5373 => x"C0C0C0C092B0F8B0",
  5374 => x"C0C0C0C092B0F899",
  5375 => x"C0C0C0C092B0F892",
  5376 => x"C0C0C0C092B0F882",
  5377 => x"C0C0C0C092B0F8F8",
  5378 => x"C0C0C0C092B0F880",
  5379 => x"C0C0C0C092B0F890",
  5380 => x"C0C0C0C092B080C0",
  5381 => x"C0C0C0C092B080F9",
  5382 => x"C0C0C0C092B080A4",
  5383 => x"C0C0C0C092B080B0",
  5384 => x"C0C0C0C092B08099",
  5385 => x"C0C0C0C092B08092",
  5386 => x"C0C0C0C092B08082",
  5387 => x"C0C0C0C092B080F8",
  5388 => x"C0C0C0C092B08080",
  5389 => x"C0C0C0C092B08090",
  5390 => x"C0C0C0C092B090C0",
  5391 => x"C0C0C0C092B090F9",
  5392 => x"C0C0C0C092B090A4",
  5393 => x"C0C0C0C092B090B0",
  5394 => x"C0C0C0C092B09099",
  5395 => x"C0C0C0C092B09092",
  5396 => x"C0C0C0C092B09082",
  5397 => x"C0C0C0C092B090F8",
  5398 => x"C0C0C0C092B09080",
  5399 => x"C0C0C0C092B09090",
  5400 => x"C0C0C0C09299C0C0",
  5401 => x"C0C0C0C09299C0F9",
  5402 => x"C0C0C0C09299C0A4",
  5403 => x"C0C0C0C09299C0B0",
  5404 => x"C0C0C0C09299C099",
  5405 => x"C0C0C0C09299C092",
  5406 => x"C0C0C0C09299C082",
  5407 => x"C0C0C0C09299C0F8",
  5408 => x"C0C0C0C09299C080",
  5409 => x"C0C0C0C09299C090",
  5410 => x"C0C0C0C09299F9C0",
  5411 => x"C0C0C0C09299F9F9",
  5412 => x"C0C0C0C09299F9A4",
  5413 => x"C0C0C0C09299F9B0",
  5414 => x"C0C0C0C09299F999",
  5415 => x"C0C0C0C09299F992",
  5416 => x"C0C0C0C09299F982",
  5417 => x"C0C0C0C09299F9F8",
  5418 => x"C0C0C0C09299F980",
  5419 => x"C0C0C0C09299F990",
  5420 => x"C0C0C0C09299A4C0",
  5421 => x"C0C0C0C09299A4F9",
  5422 => x"C0C0C0C09299A4A4",
  5423 => x"C0C0C0C09299A4B0",
  5424 => x"C0C0C0C09299A499",
  5425 => x"C0C0C0C09299A492",
  5426 => x"C0C0C0C09299A482",
  5427 => x"C0C0C0C09299A4F8",
  5428 => x"C0C0C0C09299A480",
  5429 => x"C0C0C0C09299A490",
  5430 => x"C0C0C0C09299B0C0",
  5431 => x"C0C0C0C09299B0F9",
  5432 => x"C0C0C0C09299B0A4",
  5433 => x"C0C0C0C09299B0B0",
  5434 => x"C0C0C0C09299B099",
  5435 => x"C0C0C0C09299B092",
  5436 => x"C0C0C0C09299B082",
  5437 => x"C0C0C0C09299B0F8",
  5438 => x"C0C0C0C09299B080",
  5439 => x"C0C0C0C09299B090",
  5440 => x"C0C0C0C0929999C0",
  5441 => x"C0C0C0C0929999F9",
  5442 => x"C0C0C0C0929999A4",
  5443 => x"C0C0C0C0929999B0",
  5444 => x"C0C0C0C092999999",
  5445 => x"C0C0C0C092999992",
  5446 => x"C0C0C0C092999982",
  5447 => x"C0C0C0C0929999F8",
  5448 => x"C0C0C0C092999980",
  5449 => x"C0C0C0C092999990",
  5450 => x"C0C0C0C0929992C0",
  5451 => x"C0C0C0C0929992F9",
  5452 => x"C0C0C0C0929992A4",
  5453 => x"C0C0C0C0929992B0",
  5454 => x"C0C0C0C092999299",
  5455 => x"C0C0C0C092999292",
  5456 => x"C0C0C0C092999282",
  5457 => x"C0C0C0C0929992F8",
  5458 => x"C0C0C0C092999280",
  5459 => x"C0C0C0C092999290",
  5460 => x"C0C0C0C0929982C0",
  5461 => x"C0C0C0C0929982F9",
  5462 => x"C0C0C0C0929982A4",
  5463 => x"C0C0C0C0929982B0",
  5464 => x"C0C0C0C092998299",
  5465 => x"C0C0C0C092998292",
  5466 => x"C0C0C0C092998282",
  5467 => x"C0C0C0C0929982F8",
  5468 => x"C0C0C0C092998280",
  5469 => x"C0C0C0C092998290",
  5470 => x"C0C0C0C09299F8C0",
  5471 => x"C0C0C0C09299F8F9",
  5472 => x"C0C0C0C09299F8A4",
  5473 => x"C0C0C0C09299F8B0",
  5474 => x"C0C0C0C09299F899",
  5475 => x"C0C0C0C09299F892",
  5476 => x"C0C0C0C09299F882",
  5477 => x"C0C0C0C09299F8F8",
  5478 => x"C0C0C0C09299F880",
  5479 => x"C0C0C0C09299F890",
  5480 => x"C0C0C0C0929980C0",
  5481 => x"C0C0C0C0929980F9",
  5482 => x"C0C0C0C0929980A4",
  5483 => x"C0C0C0C0929980B0",
  5484 => x"C0C0C0C092998099",
  5485 => x"C0C0C0C092998092",
  5486 => x"C0C0C0C092998082",
  5487 => x"C0C0C0C0929980F8",
  5488 => x"C0C0C0C092998080",
  5489 => x"C0C0C0C092998090",
  5490 => x"C0C0C0C0929990C0",
  5491 => x"C0C0C0C0929990F9",
  5492 => x"C0C0C0C0929990A4",
  5493 => x"C0C0C0C0929990B0",
  5494 => x"C0C0C0C092999099",
  5495 => x"C0C0C0C092999092",
  5496 => x"C0C0C0C092999082",
  5497 => x"C0C0C0C0929990F8",
  5498 => x"C0C0C0C092999080",
  5499 => x"C0C0C0C092999090",
  5500 => x"C0C0C0C09292C0C0",
  5501 => x"C0C0C0C09292C0F9",
  5502 => x"C0C0C0C09292C0A4",
  5503 => x"C0C0C0C09292C0B0",
  5504 => x"C0C0C0C09292C099",
  5505 => x"C0C0C0C09292C092",
  5506 => x"C0C0C0C09292C082",
  5507 => x"C0C0C0C09292C0F8",
  5508 => x"C0C0C0C09292C080",
  5509 => x"C0C0C0C09292C090",
  5510 => x"C0C0C0C09292F9C0",
  5511 => x"C0C0C0C09292F9F9",
  5512 => x"C0C0C0C09292F9A4",
  5513 => x"C0C0C0C09292F9B0",
  5514 => x"C0C0C0C09292F999",
  5515 => x"C0C0C0C09292F992",
  5516 => x"C0C0C0C09292F982",
  5517 => x"C0C0C0C09292F9F8",
  5518 => x"C0C0C0C09292F980",
  5519 => x"C0C0C0C09292F990",
  5520 => x"C0C0C0C09292A4C0",
  5521 => x"C0C0C0C09292A4F9",
  5522 => x"C0C0C0C09292A4A4",
  5523 => x"C0C0C0C09292A4B0",
  5524 => x"C0C0C0C09292A499",
  5525 => x"C0C0C0C09292A492",
  5526 => x"C0C0C0C09292A482",
  5527 => x"C0C0C0C09292A4F8",
  5528 => x"C0C0C0C09292A480",
  5529 => x"C0C0C0C09292A490",
  5530 => x"C0C0C0C09292B0C0",
  5531 => x"C0C0C0C09292B0F9",
  5532 => x"C0C0C0C09292B0A4",
  5533 => x"C0C0C0C09292B0B0",
  5534 => x"C0C0C0C09292B099",
  5535 => x"C0C0C0C09292B092",
  5536 => x"C0C0C0C09292B082",
  5537 => x"C0C0C0C09292B0F8",
  5538 => x"C0C0C0C09292B080",
  5539 => x"C0C0C0C09292B090",
  5540 => x"C0C0C0C0929299C0",
  5541 => x"C0C0C0C0929299F9",
  5542 => x"C0C0C0C0929299A4",
  5543 => x"C0C0C0C0929299B0",
  5544 => x"C0C0C0C092929999",
  5545 => x"C0C0C0C092929992",
  5546 => x"C0C0C0C092929982",
  5547 => x"C0C0C0C0929299F8",
  5548 => x"C0C0C0C092929980",
  5549 => x"C0C0C0C092929990",
  5550 => x"C0C0C0C0929292C0",
  5551 => x"C0C0C0C0929292F9",
  5552 => x"C0C0C0C0929292A4",
  5553 => x"C0C0C0C0929292B0",
  5554 => x"C0C0C0C092929299",
  5555 => x"C0C0C0C092929292",
  5556 => x"C0C0C0C092929282",
  5557 => x"C0C0C0C0929292F8",
  5558 => x"C0C0C0C092929280",
  5559 => x"C0C0C0C092929290",
  5560 => x"C0C0C0C0929282C0",
  5561 => x"C0C0C0C0929282F9",
  5562 => x"C0C0C0C0929282A4",
  5563 => x"C0C0C0C0929282B0",
  5564 => x"C0C0C0C092928299",
  5565 => x"C0C0C0C092928292",
  5566 => x"C0C0C0C092928282",
  5567 => x"C0C0C0C0929282F8",
  5568 => x"C0C0C0C092928280",
  5569 => x"C0C0C0C092928290",
  5570 => x"C0C0C0C09292F8C0",
  5571 => x"C0C0C0C09292F8F9",
  5572 => x"C0C0C0C09292F8A4",
  5573 => x"C0C0C0C09292F8B0",
  5574 => x"C0C0C0C09292F899",
  5575 => x"C0C0C0C09292F892",
  5576 => x"C0C0C0C09292F882",
  5577 => x"C0C0C0C09292F8F8",
  5578 => x"C0C0C0C09292F880",
  5579 => x"C0C0C0C09292F890",
  5580 => x"C0C0C0C0929280C0",
  5581 => x"C0C0C0C0929280F9",
  5582 => x"C0C0C0C0929280A4",
  5583 => x"C0C0C0C0929280B0",
  5584 => x"C0C0C0C092928099",
  5585 => x"C0C0C0C092928092",
  5586 => x"C0C0C0C092928082",
  5587 => x"C0C0C0C0929280F8",
  5588 => x"C0C0C0C092928080",
  5589 => x"C0C0C0C092928090",
  5590 => x"C0C0C0C0929290C0",
  5591 => x"C0C0C0C0929290F9",
  5592 => x"C0C0C0C0929290A4",
  5593 => x"C0C0C0C0929290B0",
  5594 => x"C0C0C0C092929099",
  5595 => x"C0C0C0C092929092",
  5596 => x"C0C0C0C092929082",
  5597 => x"C0C0C0C0929290F8",
  5598 => x"C0C0C0C092929080",
  5599 => x"C0C0C0C092929090",
  5600 => x"C0C0C0C09282C0C0",
  5601 => x"C0C0C0C09282C0F9",
  5602 => x"C0C0C0C09282C0A4",
  5603 => x"C0C0C0C09282C0B0",
  5604 => x"C0C0C0C09282C099",
  5605 => x"C0C0C0C09282C092",
  5606 => x"C0C0C0C09282C082",
  5607 => x"C0C0C0C09282C0F8",
  5608 => x"C0C0C0C09282C080",
  5609 => x"C0C0C0C09282C090",
  5610 => x"C0C0C0C09282F9C0",
  5611 => x"C0C0C0C09282F9F9",
  5612 => x"C0C0C0C09282F9A4",
  5613 => x"C0C0C0C09282F9B0",
  5614 => x"C0C0C0C09282F999",
  5615 => x"C0C0C0C09282F992",
  5616 => x"C0C0C0C09282F982",
  5617 => x"C0C0C0C09282F9F8",
  5618 => x"C0C0C0C09282F980",
  5619 => x"C0C0C0C09282F990",
  5620 => x"C0C0C0C09282A4C0",
  5621 => x"C0C0C0C09282A4F9",
  5622 => x"C0C0C0C09282A4A4",
  5623 => x"C0C0C0C09282A4B0",
  5624 => x"C0C0C0C09282A499",
  5625 => x"C0C0C0C09282A492",
  5626 => x"C0C0C0C09282A482",
  5627 => x"C0C0C0C09282A4F8",
  5628 => x"C0C0C0C09282A480",
  5629 => x"C0C0C0C09282A490",
  5630 => x"C0C0C0C09282B0C0",
  5631 => x"C0C0C0C09282B0F9",
  5632 => x"C0C0C0C09282B0A4",
  5633 => x"C0C0C0C09282B0B0",
  5634 => x"C0C0C0C09282B099",
  5635 => x"C0C0C0C09282B092",
  5636 => x"C0C0C0C09282B082",
  5637 => x"C0C0C0C09282B0F8",
  5638 => x"C0C0C0C09282B080",
  5639 => x"C0C0C0C09282B090",
  5640 => x"C0C0C0C0928299C0",
  5641 => x"C0C0C0C0928299F9",
  5642 => x"C0C0C0C0928299A4",
  5643 => x"C0C0C0C0928299B0",
  5644 => x"C0C0C0C092829999",
  5645 => x"C0C0C0C092829992",
  5646 => x"C0C0C0C092829982",
  5647 => x"C0C0C0C0928299F8",
  5648 => x"C0C0C0C092829980",
  5649 => x"C0C0C0C092829990",
  5650 => x"C0C0C0C0928292C0",
  5651 => x"C0C0C0C0928292F9",
  5652 => x"C0C0C0C0928292A4",
  5653 => x"C0C0C0C0928292B0",
  5654 => x"C0C0C0C092829299",
  5655 => x"C0C0C0C092829292",
  5656 => x"C0C0C0C092829282",
  5657 => x"C0C0C0C0928292F8",
  5658 => x"C0C0C0C092829280",
  5659 => x"C0C0C0C092829290",
  5660 => x"C0C0C0C0928282C0",
  5661 => x"C0C0C0C0928282F9",
  5662 => x"C0C0C0C0928282A4",
  5663 => x"C0C0C0C0928282B0",
  5664 => x"C0C0C0C092828299",
  5665 => x"C0C0C0C092828292",
  5666 => x"C0C0C0C092828282",
  5667 => x"C0C0C0C0928282F8",
  5668 => x"C0C0C0C092828280",
  5669 => x"C0C0C0C092828290",
  5670 => x"C0C0C0C09282F8C0",
  5671 => x"C0C0C0C09282F8F9",
  5672 => x"C0C0C0C09282F8A4",
  5673 => x"C0C0C0C09282F8B0",
  5674 => x"C0C0C0C09282F899",
  5675 => x"C0C0C0C09282F892",
  5676 => x"C0C0C0C09282F882",
  5677 => x"C0C0C0C09282F8F8",
  5678 => x"C0C0C0C09282F880",
  5679 => x"C0C0C0C09282F890",
  5680 => x"C0C0C0C0928280C0",
  5681 => x"C0C0C0C0928280F9",
  5682 => x"C0C0C0C0928280A4",
  5683 => x"C0C0C0C0928280B0",
  5684 => x"C0C0C0C092828099",
  5685 => x"C0C0C0C092828092",
  5686 => x"C0C0C0C092828082",
  5687 => x"C0C0C0C0928280F8",
  5688 => x"C0C0C0C092828080",
  5689 => x"C0C0C0C092828090",
  5690 => x"C0C0C0C0928290C0",
  5691 => x"C0C0C0C0928290F9",
  5692 => x"C0C0C0C0928290A4",
  5693 => x"C0C0C0C0928290B0",
  5694 => x"C0C0C0C092829099",
  5695 => x"C0C0C0C092829092",
  5696 => x"C0C0C0C092829082",
  5697 => x"C0C0C0C0928290F8",
  5698 => x"C0C0C0C092829080",
  5699 => x"C0C0C0C092829090",
  5700 => x"C0C0C0C092F8C0C0",
  5701 => x"C0C0C0C092F8C0F9",
  5702 => x"C0C0C0C092F8C0A4",
  5703 => x"C0C0C0C092F8C0B0",
  5704 => x"C0C0C0C092F8C099",
  5705 => x"C0C0C0C092F8C092",
  5706 => x"C0C0C0C092F8C082",
  5707 => x"C0C0C0C092F8C0F8",
  5708 => x"C0C0C0C092F8C080",
  5709 => x"C0C0C0C092F8C090",
  5710 => x"C0C0C0C092F8F9C0",
  5711 => x"C0C0C0C092F8F9F9",
  5712 => x"C0C0C0C092F8F9A4",
  5713 => x"C0C0C0C092F8F9B0",
  5714 => x"C0C0C0C092F8F999",
  5715 => x"C0C0C0C092F8F992",
  5716 => x"C0C0C0C092F8F982",
  5717 => x"C0C0C0C092F8F9F8",
  5718 => x"C0C0C0C092F8F980",
  5719 => x"C0C0C0C092F8F990",
  5720 => x"C0C0C0C092F8A4C0",
  5721 => x"C0C0C0C092F8A4F9",
  5722 => x"C0C0C0C092F8A4A4",
  5723 => x"C0C0C0C092F8A4B0",
  5724 => x"C0C0C0C092F8A499",
  5725 => x"C0C0C0C092F8A492",
  5726 => x"C0C0C0C092F8A482",
  5727 => x"C0C0C0C092F8A4F8",
  5728 => x"C0C0C0C092F8A480",
  5729 => x"C0C0C0C092F8A490",
  5730 => x"C0C0C0C092F8B0C0",
  5731 => x"C0C0C0C092F8B0F9",
  5732 => x"C0C0C0C092F8B0A4",
  5733 => x"C0C0C0C092F8B0B0",
  5734 => x"C0C0C0C092F8B099",
  5735 => x"C0C0C0C092F8B092",
  5736 => x"C0C0C0C092F8B082",
  5737 => x"C0C0C0C092F8B0F8",
  5738 => x"C0C0C0C092F8B080",
  5739 => x"C0C0C0C092F8B090",
  5740 => x"C0C0C0C092F899C0",
  5741 => x"C0C0C0C092F899F9",
  5742 => x"C0C0C0C092F899A4",
  5743 => x"C0C0C0C092F899B0",
  5744 => x"C0C0C0C092F89999",
  5745 => x"C0C0C0C092F89992",
  5746 => x"C0C0C0C092F89982",
  5747 => x"C0C0C0C092F899F8",
  5748 => x"C0C0C0C092F89980",
  5749 => x"C0C0C0C092F89990",
  5750 => x"C0C0C0C092F892C0",
  5751 => x"C0C0C0C092F892F9",
  5752 => x"C0C0C0C092F892A4",
  5753 => x"C0C0C0C092F892B0",
  5754 => x"C0C0C0C092F89299",
  5755 => x"C0C0C0C092F89292",
  5756 => x"C0C0C0C092F89282",
  5757 => x"C0C0C0C092F892F8",
  5758 => x"C0C0C0C092F89280",
  5759 => x"C0C0C0C092F89290",
  5760 => x"C0C0C0C092F882C0",
  5761 => x"C0C0C0C092F882F9",
  5762 => x"C0C0C0C092F882A4",
  5763 => x"C0C0C0C092F882B0",
  5764 => x"C0C0C0C092F88299",
  5765 => x"C0C0C0C092F88292",
  5766 => x"C0C0C0C092F88282",
  5767 => x"C0C0C0C092F882F8",
  5768 => x"C0C0C0C092F88280",
  5769 => x"C0C0C0C092F88290",
  5770 => x"C0C0C0C092F8F8C0",
  5771 => x"C0C0C0C092F8F8F9",
  5772 => x"C0C0C0C092F8F8A4",
  5773 => x"C0C0C0C092F8F8B0",
  5774 => x"C0C0C0C092F8F899",
  5775 => x"C0C0C0C092F8F892",
  5776 => x"C0C0C0C092F8F882",
  5777 => x"C0C0C0C092F8F8F8",
  5778 => x"C0C0C0C092F8F880",
  5779 => x"C0C0C0C092F8F890",
  5780 => x"C0C0C0C092F880C0",
  5781 => x"C0C0C0C092F880F9",
  5782 => x"C0C0C0C092F880A4",
  5783 => x"C0C0C0C092F880B0",
  5784 => x"C0C0C0C092F88099",
  5785 => x"C0C0C0C092F88092",
  5786 => x"C0C0C0C092F88082",
  5787 => x"C0C0C0C092F880F8",
  5788 => x"C0C0C0C092F88080",
  5789 => x"C0C0C0C092F88090",
  5790 => x"C0C0C0C092F890C0",
  5791 => x"C0C0C0C092F890F9",
  5792 => x"C0C0C0C092F890A4",
  5793 => x"C0C0C0C092F890B0",
  5794 => x"C0C0C0C092F89099",
  5795 => x"C0C0C0C092F89092",
  5796 => x"C0C0C0C092F89082",
  5797 => x"C0C0C0C092F890F8",
  5798 => x"C0C0C0C092F89080",
  5799 => x"C0C0C0C092F89090",
  5800 => x"C0C0C0C09280C0C0",
  5801 => x"C0C0C0C09280C0F9",
  5802 => x"C0C0C0C09280C0A4",
  5803 => x"C0C0C0C09280C0B0",
  5804 => x"C0C0C0C09280C099",
  5805 => x"C0C0C0C09280C092",
  5806 => x"C0C0C0C09280C082",
  5807 => x"C0C0C0C09280C0F8",
  5808 => x"C0C0C0C09280C080",
  5809 => x"C0C0C0C09280C090",
  5810 => x"C0C0C0C09280F9C0",
  5811 => x"C0C0C0C09280F9F9",
  5812 => x"C0C0C0C09280F9A4",
  5813 => x"C0C0C0C09280F9B0",
  5814 => x"C0C0C0C09280F999",
  5815 => x"C0C0C0C09280F992",
  5816 => x"C0C0C0C09280F982",
  5817 => x"C0C0C0C09280F9F8",
  5818 => x"C0C0C0C09280F980",
  5819 => x"C0C0C0C09280F990",
  5820 => x"C0C0C0C09280A4C0",
  5821 => x"C0C0C0C09280A4F9",
  5822 => x"C0C0C0C09280A4A4",
  5823 => x"C0C0C0C09280A4B0",
  5824 => x"C0C0C0C09280A499",
  5825 => x"C0C0C0C09280A492",
  5826 => x"C0C0C0C09280A482",
  5827 => x"C0C0C0C09280A4F8",
  5828 => x"C0C0C0C09280A480",
  5829 => x"C0C0C0C09280A490",
  5830 => x"C0C0C0C09280B0C0",
  5831 => x"C0C0C0C09280B0F9",
  5832 => x"C0C0C0C09280B0A4",
  5833 => x"C0C0C0C09280B0B0",
  5834 => x"C0C0C0C09280B099",
  5835 => x"C0C0C0C09280B092",
  5836 => x"C0C0C0C09280B082",
  5837 => x"C0C0C0C09280B0F8",
  5838 => x"C0C0C0C09280B080",
  5839 => x"C0C0C0C09280B090",
  5840 => x"C0C0C0C0928099C0",
  5841 => x"C0C0C0C0928099F9",
  5842 => x"C0C0C0C0928099A4",
  5843 => x"C0C0C0C0928099B0",
  5844 => x"C0C0C0C092809999",
  5845 => x"C0C0C0C092809992",
  5846 => x"C0C0C0C092809982",
  5847 => x"C0C0C0C0928099F8",
  5848 => x"C0C0C0C092809980",
  5849 => x"C0C0C0C092809990",
  5850 => x"C0C0C0C0928092C0",
  5851 => x"C0C0C0C0928092F9",
  5852 => x"C0C0C0C0928092A4",
  5853 => x"C0C0C0C0928092B0",
  5854 => x"C0C0C0C092809299",
  5855 => x"C0C0C0C092809292",
  5856 => x"C0C0C0C092809282",
  5857 => x"C0C0C0C0928092F8",
  5858 => x"C0C0C0C092809280",
  5859 => x"C0C0C0C092809290",
  5860 => x"C0C0C0C0928082C0",
  5861 => x"C0C0C0C0928082F9",
  5862 => x"C0C0C0C0928082A4",
  5863 => x"C0C0C0C0928082B0",
  5864 => x"C0C0C0C092808299",
  5865 => x"C0C0C0C092808292",
  5866 => x"C0C0C0C092808282",
  5867 => x"C0C0C0C0928082F8",
  5868 => x"C0C0C0C092808280",
  5869 => x"C0C0C0C092808290",
  5870 => x"C0C0C0C09280F8C0",
  5871 => x"C0C0C0C09280F8F9",
  5872 => x"C0C0C0C09280F8A4",
  5873 => x"C0C0C0C09280F8B0",
  5874 => x"C0C0C0C09280F899",
  5875 => x"C0C0C0C09280F892",
  5876 => x"C0C0C0C09280F882",
  5877 => x"C0C0C0C09280F8F8",
  5878 => x"C0C0C0C09280F880",
  5879 => x"C0C0C0C09280F890",
  5880 => x"C0C0C0C0928080C0",
  5881 => x"C0C0C0C0928080F9",
  5882 => x"C0C0C0C0928080A4",
  5883 => x"C0C0C0C0928080B0",
  5884 => x"C0C0C0C092808099",
  5885 => x"C0C0C0C092808092",
  5886 => x"C0C0C0C092808082",
  5887 => x"C0C0C0C0928080F8",
  5888 => x"C0C0C0C092808080",
  5889 => x"C0C0C0C092808090",
  5890 => x"C0C0C0C0928090C0",
  5891 => x"C0C0C0C0928090F9",
  5892 => x"C0C0C0C0928090A4",
  5893 => x"C0C0C0C0928090B0",
  5894 => x"C0C0C0C092809099",
  5895 => x"C0C0C0C092809092",
  5896 => x"C0C0C0C092809082",
  5897 => x"C0C0C0C0928090F8",
  5898 => x"C0C0C0C092809080",
  5899 => x"C0C0C0C092809090",
  5900 => x"C0C0C0C09290C0C0",
  5901 => x"C0C0C0C09290C0F9",
  5902 => x"C0C0C0C09290C0A4",
  5903 => x"C0C0C0C09290C0B0",
  5904 => x"C0C0C0C09290C099",
  5905 => x"C0C0C0C09290C092",
  5906 => x"C0C0C0C09290C082",
  5907 => x"C0C0C0C09290C0F8",
  5908 => x"C0C0C0C09290C080",
  5909 => x"C0C0C0C09290C090",
  5910 => x"C0C0C0C09290F9C0",
  5911 => x"C0C0C0C09290F9F9",
  5912 => x"C0C0C0C09290F9A4",
  5913 => x"C0C0C0C09290F9B0",
  5914 => x"C0C0C0C09290F999",
  5915 => x"C0C0C0C09290F992",
  5916 => x"C0C0C0C09290F982",
  5917 => x"C0C0C0C09290F9F8",
  5918 => x"C0C0C0C09290F980",
  5919 => x"C0C0C0C09290F990",
  5920 => x"C0C0C0C09290A4C0",
  5921 => x"C0C0C0C09290A4F9",
  5922 => x"C0C0C0C09290A4A4",
  5923 => x"C0C0C0C09290A4B0",
  5924 => x"C0C0C0C09290A499",
  5925 => x"C0C0C0C09290A492",
  5926 => x"C0C0C0C09290A482",
  5927 => x"C0C0C0C09290A4F8",
  5928 => x"C0C0C0C09290A480",
  5929 => x"C0C0C0C09290A490",
  5930 => x"C0C0C0C09290B0C0",
  5931 => x"C0C0C0C09290B0F9",
  5932 => x"C0C0C0C09290B0A4",
  5933 => x"C0C0C0C09290B0B0",
  5934 => x"C0C0C0C09290B099",
  5935 => x"C0C0C0C09290B092",
  5936 => x"C0C0C0C09290B082",
  5937 => x"C0C0C0C09290B0F8",
  5938 => x"C0C0C0C09290B080",
  5939 => x"C0C0C0C09290B090",
  5940 => x"C0C0C0C0929099C0",
  5941 => x"C0C0C0C0929099F9",
  5942 => x"C0C0C0C0929099A4",
  5943 => x"C0C0C0C0929099B0",
  5944 => x"C0C0C0C092909999",
  5945 => x"C0C0C0C092909992",
  5946 => x"C0C0C0C092909982",
  5947 => x"C0C0C0C0929099F8",
  5948 => x"C0C0C0C092909980",
  5949 => x"C0C0C0C092909990",
  5950 => x"C0C0C0C0929092C0",
  5951 => x"C0C0C0C0929092F9",
  5952 => x"C0C0C0C0929092A4",
  5953 => x"C0C0C0C0929092B0",
  5954 => x"C0C0C0C092909299",
  5955 => x"C0C0C0C092909292",
  5956 => x"C0C0C0C092909282",
  5957 => x"C0C0C0C0929092F8",
  5958 => x"C0C0C0C092909280",
  5959 => x"C0C0C0C092909290",
  5960 => x"C0C0C0C0929082C0",
  5961 => x"C0C0C0C0929082F9",
  5962 => x"C0C0C0C0929082A4",
  5963 => x"C0C0C0C0929082B0",
  5964 => x"C0C0C0C092908299",
  5965 => x"C0C0C0C092908292",
  5966 => x"C0C0C0C092908282",
  5967 => x"C0C0C0C0929082F8",
  5968 => x"C0C0C0C092908280",
  5969 => x"C0C0C0C092908290",
  5970 => x"C0C0C0C09290F8C0",
  5971 => x"C0C0C0C09290F8F9",
  5972 => x"C0C0C0C09290F8A4",
  5973 => x"C0C0C0C09290F8B0",
  5974 => x"C0C0C0C09290F899",
  5975 => x"C0C0C0C09290F892",
  5976 => x"C0C0C0C09290F882",
  5977 => x"C0C0C0C09290F8F8",
  5978 => x"C0C0C0C09290F880",
  5979 => x"C0C0C0C09290F890",
  5980 => x"C0C0C0C0929080C0",
  5981 => x"C0C0C0C0929080F9",
  5982 => x"C0C0C0C0929080A4",
  5983 => x"C0C0C0C0929080B0",
  5984 => x"C0C0C0C092908099",
  5985 => x"C0C0C0C092908092",
  5986 => x"C0C0C0C092908082",
  5987 => x"C0C0C0C0929080F8",
  5988 => x"C0C0C0C092908080",
  5989 => x"C0C0C0C092908090",
  5990 => x"C0C0C0C0929090C0",
  5991 => x"C0C0C0C0929090F9",
  5992 => x"C0C0C0C0929090A4",
  5993 => x"C0C0C0C0929090B0",
  5994 => x"C0C0C0C092909099",
  5995 => x"C0C0C0C092909092",
  5996 => x"C0C0C0C092909082",
  5997 => x"C0C0C0C0929090F8",
  5998 => x"C0C0C0C092909080",
  5999 => x"C0C0C0C092909090",
  6000 => x"C0C0C0C082C0C0C0",
  6001 => x"C0C0C0C082C0C0F9",
  6002 => x"C0C0C0C082C0C0A4",
  6003 => x"C0C0C0C082C0C0B0",
  6004 => x"C0C0C0C082C0C099",
  6005 => x"C0C0C0C082C0C092",
  6006 => x"C0C0C0C082C0C082",
  6007 => x"C0C0C0C082C0C0F8",
  6008 => x"C0C0C0C082C0C080",
  6009 => x"C0C0C0C082C0C090",
  6010 => x"C0C0C0C082C0F9C0",
  6011 => x"C0C0C0C082C0F9F9",
  6012 => x"C0C0C0C082C0F9A4",
  6013 => x"C0C0C0C082C0F9B0",
  6014 => x"C0C0C0C082C0F999",
  6015 => x"C0C0C0C082C0F992",
  6016 => x"C0C0C0C082C0F982",
  6017 => x"C0C0C0C082C0F9F8",
  6018 => x"C0C0C0C082C0F980",
  6019 => x"C0C0C0C082C0F990",
  6020 => x"C0C0C0C082C0A4C0",
  6021 => x"C0C0C0C082C0A4F9",
  6022 => x"C0C0C0C082C0A4A4",
  6023 => x"C0C0C0C082C0A4B0",
  6024 => x"C0C0C0C082C0A499",
  6025 => x"C0C0C0C082C0A492",
  6026 => x"C0C0C0C082C0A482",
  6027 => x"C0C0C0C082C0A4F8",
  6028 => x"C0C0C0C082C0A480",
  6029 => x"C0C0C0C082C0A490",
  6030 => x"C0C0C0C082C0B0C0",
  6031 => x"C0C0C0C082C0B0F9",
  6032 => x"C0C0C0C082C0B0A4",
  6033 => x"C0C0C0C082C0B0B0",
  6034 => x"C0C0C0C082C0B099",
  6035 => x"C0C0C0C082C0B092",
  6036 => x"C0C0C0C082C0B082",
  6037 => x"C0C0C0C082C0B0F8",
  6038 => x"C0C0C0C082C0B080",
  6039 => x"C0C0C0C082C0B090",
  6040 => x"C0C0C0C082C099C0",
  6041 => x"C0C0C0C082C099F9",
  6042 => x"C0C0C0C082C099A4",
  6043 => x"C0C0C0C082C099B0",
  6044 => x"C0C0C0C082C09999",
  6045 => x"C0C0C0C082C09992",
  6046 => x"C0C0C0C082C09982",
  6047 => x"C0C0C0C082C099F8",
  6048 => x"C0C0C0C082C09980",
  6049 => x"C0C0C0C082C09990",
  6050 => x"C0C0C0C082C092C0",
  6051 => x"C0C0C0C082C092F9",
  6052 => x"C0C0C0C082C092A4",
  6053 => x"C0C0C0C082C092B0",
  6054 => x"C0C0C0C082C09299",
  6055 => x"C0C0C0C082C09292",
  6056 => x"C0C0C0C082C09282",
  6057 => x"C0C0C0C082C092F8",
  6058 => x"C0C0C0C082C09280",
  6059 => x"C0C0C0C082C09290",
  6060 => x"C0C0C0C082C082C0",
  6061 => x"C0C0C0C082C082F9",
  6062 => x"C0C0C0C082C082A4",
  6063 => x"C0C0C0C082C082B0",
  6064 => x"C0C0C0C082C08299",
  6065 => x"C0C0C0C082C08292",
  6066 => x"C0C0C0C082C08282",
  6067 => x"C0C0C0C082C082F8",
  6068 => x"C0C0C0C082C08280",
  6069 => x"C0C0C0C082C08290",
  6070 => x"C0C0C0C082C0F8C0",
  6071 => x"C0C0C0C082C0F8F9",
  6072 => x"C0C0C0C082C0F8A4",
  6073 => x"C0C0C0C082C0F8B0",
  6074 => x"C0C0C0C082C0F899",
  6075 => x"C0C0C0C082C0F892",
  6076 => x"C0C0C0C082C0F882",
  6077 => x"C0C0C0C082C0F8F8",
  6078 => x"C0C0C0C082C0F880",
  6079 => x"C0C0C0C082C0F890",
  6080 => x"C0C0C0C082C080C0",
  6081 => x"C0C0C0C082C080F9",
  6082 => x"C0C0C0C082C080A4",
  6083 => x"C0C0C0C082C080B0",
  6084 => x"C0C0C0C082C08099",
  6085 => x"C0C0C0C082C08092",
  6086 => x"C0C0C0C082C08082",
  6087 => x"C0C0C0C082C080F8",
  6088 => x"C0C0C0C082C08080",
  6089 => x"C0C0C0C082C08090",
  6090 => x"C0C0C0C082C090C0",
  6091 => x"C0C0C0C082C090F9",
  6092 => x"C0C0C0C082C090A4",
  6093 => x"C0C0C0C082C090B0",
  6094 => x"C0C0C0C082C09099",
  6095 => x"C0C0C0C082C09092",
  6096 => x"C0C0C0C082C09082",
  6097 => x"C0C0C0C082C090F8",
  6098 => x"C0C0C0C082C09080",
  6099 => x"C0C0C0C082C09090",
  6100 => x"C0C0C0C082F9C0C0",
  6101 => x"C0C0C0C082F9C0F9",
  6102 => x"C0C0C0C082F9C0A4",
  6103 => x"C0C0C0C082F9C0B0",
  6104 => x"C0C0C0C082F9C099",
  6105 => x"C0C0C0C082F9C092",
  6106 => x"C0C0C0C082F9C082",
  6107 => x"C0C0C0C082F9C0F8",
  6108 => x"C0C0C0C082F9C080",
  6109 => x"C0C0C0C082F9C090",
  6110 => x"C0C0C0C082F9F9C0",
  6111 => x"C0C0C0C082F9F9F9",
  6112 => x"C0C0C0C082F9F9A4",
  6113 => x"C0C0C0C082F9F9B0",
  6114 => x"C0C0C0C082F9F999",
  6115 => x"C0C0C0C082F9F992",
  6116 => x"C0C0C0C082F9F982",
  6117 => x"C0C0C0C082F9F9F8",
  6118 => x"C0C0C0C082F9F980",
  6119 => x"C0C0C0C082F9F990",
  6120 => x"C0C0C0C082F9A4C0",
  6121 => x"C0C0C0C082F9A4F9",
  6122 => x"C0C0C0C082F9A4A4",
  6123 => x"C0C0C0C082F9A4B0",
  6124 => x"C0C0C0C082F9A499",
  6125 => x"C0C0C0C082F9A492",
  6126 => x"C0C0C0C082F9A482",
  6127 => x"C0C0C0C082F9A4F8",
  6128 => x"C0C0C0C082F9A480",
  6129 => x"C0C0C0C082F9A490",
  6130 => x"C0C0C0C082F9B0C0",
  6131 => x"C0C0C0C082F9B0F9",
  6132 => x"C0C0C0C082F9B0A4",
  6133 => x"C0C0C0C082F9B0B0",
  6134 => x"C0C0C0C082F9B099",
  6135 => x"C0C0C0C082F9B092",
  6136 => x"C0C0C0C082F9B082",
  6137 => x"C0C0C0C082F9B0F8",
  6138 => x"C0C0C0C082F9B080",
  6139 => x"C0C0C0C082F9B090",
  6140 => x"C0C0C0C082F999C0",
  6141 => x"C0C0C0C082F999F9",
  6142 => x"C0C0C0C082F999A4",
  6143 => x"C0C0C0C082F999B0",
  6144 => x"C0C0C0C082F99999",
  6145 => x"C0C0C0C082F99992",
  6146 => x"C0C0C0C082F99982",
  6147 => x"C0C0C0C082F999F8",
  6148 => x"C0C0C0C082F99980",
  6149 => x"C0C0C0C082F99990",
  6150 => x"C0C0C0C082F992C0",
  6151 => x"C0C0C0C082F992F9",
  6152 => x"C0C0C0C082F992A4",
  6153 => x"C0C0C0C082F992B0",
  6154 => x"C0C0C0C082F99299",
  6155 => x"C0C0C0C082F99292",
  6156 => x"C0C0C0C082F99282",
  6157 => x"C0C0C0C082F992F8",
  6158 => x"C0C0C0C082F99280",
  6159 => x"C0C0C0C082F99290",
  6160 => x"C0C0C0C082F982C0",
  6161 => x"C0C0C0C082F982F9",
  6162 => x"C0C0C0C082F982A4",
  6163 => x"C0C0C0C082F982B0",
  6164 => x"C0C0C0C082F98299",
  6165 => x"C0C0C0C082F98292",
  6166 => x"C0C0C0C082F98282",
  6167 => x"C0C0C0C082F982F8",
  6168 => x"C0C0C0C082F98280",
  6169 => x"C0C0C0C082F98290",
  6170 => x"C0C0C0C082F9F8C0",
  6171 => x"C0C0C0C082F9F8F9",
  6172 => x"C0C0C0C082F9F8A4",
  6173 => x"C0C0C0C082F9F8B0",
  6174 => x"C0C0C0C082F9F899",
  6175 => x"C0C0C0C082F9F892",
  6176 => x"C0C0C0C082F9F882",
  6177 => x"C0C0C0C082F9F8F8",
  6178 => x"C0C0C0C082F9F880",
  6179 => x"C0C0C0C082F9F890",
  6180 => x"C0C0C0C082F980C0",
  6181 => x"C0C0C0C082F980F9",
  6182 => x"C0C0C0C082F980A4",
  6183 => x"C0C0C0C082F980B0",
  6184 => x"C0C0C0C082F98099",
  6185 => x"C0C0C0C082F98092",
  6186 => x"C0C0C0C082F98082",
  6187 => x"C0C0C0C082F980F8",
  6188 => x"C0C0C0C082F98080",
  6189 => x"C0C0C0C082F98090",
  6190 => x"C0C0C0C082F990C0",
  6191 => x"C0C0C0C082F990F9",
  6192 => x"C0C0C0C082F990A4",
  6193 => x"C0C0C0C082F990B0",
  6194 => x"C0C0C0C082F99099",
  6195 => x"C0C0C0C082F99092",
  6196 => x"C0C0C0C082F99082",
  6197 => x"C0C0C0C082F990F8",
  6198 => x"C0C0C0C082F99080",
  6199 => x"C0C0C0C082F99090",
  6200 => x"C0C0C0C082A4C0C0",
  6201 => x"C0C0C0C082A4C0F9",
  6202 => x"C0C0C0C082A4C0A4",
  6203 => x"C0C0C0C082A4C0B0",
  6204 => x"C0C0C0C082A4C099",
  6205 => x"C0C0C0C082A4C092",
  6206 => x"C0C0C0C082A4C082",
  6207 => x"C0C0C0C082A4C0F8",
  6208 => x"C0C0C0C082A4C080",
  6209 => x"C0C0C0C082A4C090",
  6210 => x"C0C0C0C082A4F9C0",
  6211 => x"C0C0C0C082A4F9F9",
  6212 => x"C0C0C0C082A4F9A4",
  6213 => x"C0C0C0C082A4F9B0",
  6214 => x"C0C0C0C082A4F999",
  6215 => x"C0C0C0C082A4F992",
  6216 => x"C0C0C0C082A4F982",
  6217 => x"C0C0C0C082A4F9F8",
  6218 => x"C0C0C0C082A4F980",
  6219 => x"C0C0C0C082A4F990",
  6220 => x"C0C0C0C082A4A4C0",
  6221 => x"C0C0C0C082A4A4F9",
  6222 => x"C0C0C0C082A4A4A4",
  6223 => x"C0C0C0C082A4A4B0",
  6224 => x"C0C0C0C082A4A499",
  6225 => x"C0C0C0C082A4A492",
  6226 => x"C0C0C0C082A4A482",
  6227 => x"C0C0C0C082A4A4F8",
  6228 => x"C0C0C0C082A4A480",
  6229 => x"C0C0C0C082A4A490",
  6230 => x"C0C0C0C082A4B0C0",
  6231 => x"C0C0C0C082A4B0F9",
  6232 => x"C0C0C0C082A4B0A4",
  6233 => x"C0C0C0C082A4B0B0",
  6234 => x"C0C0C0C082A4B099",
  6235 => x"C0C0C0C082A4B092",
  6236 => x"C0C0C0C082A4B082",
  6237 => x"C0C0C0C082A4B0F8",
  6238 => x"C0C0C0C082A4B080",
  6239 => x"C0C0C0C082A4B090",
  6240 => x"C0C0C0C082A499C0",
  6241 => x"C0C0C0C082A499F9",
  6242 => x"C0C0C0C082A499A4",
  6243 => x"C0C0C0C082A499B0",
  6244 => x"C0C0C0C082A49999",
  6245 => x"C0C0C0C082A49992",
  6246 => x"C0C0C0C082A49982",
  6247 => x"C0C0C0C082A499F8",
  6248 => x"C0C0C0C082A49980",
  6249 => x"C0C0C0C082A49990",
  6250 => x"C0C0C0C082A492C0",
  6251 => x"C0C0C0C082A492F9",
  6252 => x"C0C0C0C082A492A4",
  6253 => x"C0C0C0C082A492B0",
  6254 => x"C0C0C0C082A49299",
  6255 => x"C0C0C0C082A49292",
  6256 => x"C0C0C0C082A49282",
  6257 => x"C0C0C0C082A492F8",
  6258 => x"C0C0C0C082A49280",
  6259 => x"C0C0C0C082A49290",
  6260 => x"C0C0C0C082A482C0",
  6261 => x"C0C0C0C082A482F9",
  6262 => x"C0C0C0C082A482A4",
  6263 => x"C0C0C0C082A482B0",
  6264 => x"C0C0C0C082A48299",
  6265 => x"C0C0C0C082A48292",
  6266 => x"C0C0C0C082A48282",
  6267 => x"C0C0C0C082A482F8",
  6268 => x"C0C0C0C082A48280",
  6269 => x"C0C0C0C082A48290",
  6270 => x"C0C0C0C082A4F8C0",
  6271 => x"C0C0C0C082A4F8F9",
  6272 => x"C0C0C0C082A4F8A4",
  6273 => x"C0C0C0C082A4F8B0",
  6274 => x"C0C0C0C082A4F899",
  6275 => x"C0C0C0C082A4F892",
  6276 => x"C0C0C0C082A4F882",
  6277 => x"C0C0C0C082A4F8F8",
  6278 => x"C0C0C0C082A4F880",
  6279 => x"C0C0C0C082A4F890",
  6280 => x"C0C0C0C082A480C0",
  6281 => x"C0C0C0C082A480F9",
  6282 => x"C0C0C0C082A480A4",
  6283 => x"C0C0C0C082A480B0",
  6284 => x"C0C0C0C082A48099",
  6285 => x"C0C0C0C082A48092",
  6286 => x"C0C0C0C082A48082",
  6287 => x"C0C0C0C082A480F8",
  6288 => x"C0C0C0C082A48080",
  6289 => x"C0C0C0C082A48090",
  6290 => x"C0C0C0C082A490C0",
  6291 => x"C0C0C0C082A490F9",
  6292 => x"C0C0C0C082A490A4",
  6293 => x"C0C0C0C082A490B0",
  6294 => x"C0C0C0C082A49099",
  6295 => x"C0C0C0C082A49092",
  6296 => x"C0C0C0C082A49082",
  6297 => x"C0C0C0C082A490F8",
  6298 => x"C0C0C0C082A49080",
  6299 => x"C0C0C0C082A49090",
  6300 => x"C0C0C0C082B0C0C0",
  6301 => x"C0C0C0C082B0C0F9",
  6302 => x"C0C0C0C082B0C0A4",
  6303 => x"C0C0C0C082B0C0B0",
  6304 => x"C0C0C0C082B0C099",
  6305 => x"C0C0C0C082B0C092",
  6306 => x"C0C0C0C082B0C082",
  6307 => x"C0C0C0C082B0C0F8",
  6308 => x"C0C0C0C082B0C080",
  6309 => x"C0C0C0C082B0C090",
  6310 => x"C0C0C0C082B0F9C0",
  6311 => x"C0C0C0C082B0F9F9",
  6312 => x"C0C0C0C082B0F9A4",
  6313 => x"C0C0C0C082B0F9B0",
  6314 => x"C0C0C0C082B0F999",
  6315 => x"C0C0C0C082B0F992",
  6316 => x"C0C0C0C082B0F982",
  6317 => x"C0C0C0C082B0F9F8",
  6318 => x"C0C0C0C082B0F980",
  6319 => x"C0C0C0C082B0F990",
  6320 => x"C0C0C0C082B0A4C0",
  6321 => x"C0C0C0C082B0A4F9",
  6322 => x"C0C0C0C082B0A4A4",
  6323 => x"C0C0C0C082B0A4B0",
  6324 => x"C0C0C0C082B0A499",
  6325 => x"C0C0C0C082B0A492",
  6326 => x"C0C0C0C082B0A482",
  6327 => x"C0C0C0C082B0A4F8",
  6328 => x"C0C0C0C082B0A480",
  6329 => x"C0C0C0C082B0A490",
  6330 => x"C0C0C0C082B0B0C0",
  6331 => x"C0C0C0C082B0B0F9",
  6332 => x"C0C0C0C082B0B0A4",
  6333 => x"C0C0C0C082B0B0B0",
  6334 => x"C0C0C0C082B0B099",
  6335 => x"C0C0C0C082B0B092",
  6336 => x"C0C0C0C082B0B082",
  6337 => x"C0C0C0C082B0B0F8",
  6338 => x"C0C0C0C082B0B080",
  6339 => x"C0C0C0C082B0B090",
  6340 => x"C0C0C0C082B099C0",
  6341 => x"C0C0C0C082B099F9",
  6342 => x"C0C0C0C082B099A4",
  6343 => x"C0C0C0C082B099B0",
  6344 => x"C0C0C0C082B09999",
  6345 => x"C0C0C0C082B09992",
  6346 => x"C0C0C0C082B09982",
  6347 => x"C0C0C0C082B099F8",
  6348 => x"C0C0C0C082B09980",
  6349 => x"C0C0C0C082B09990",
  6350 => x"C0C0C0C082B092C0",
  6351 => x"C0C0C0C082B092F9",
  6352 => x"C0C0C0C082B092A4",
  6353 => x"C0C0C0C082B092B0",
  6354 => x"C0C0C0C082B09299",
  6355 => x"C0C0C0C082B09292",
  6356 => x"C0C0C0C082B09282",
  6357 => x"C0C0C0C082B092F8",
  6358 => x"C0C0C0C082B09280",
  6359 => x"C0C0C0C082B09290",
  6360 => x"C0C0C0C082B082C0",
  6361 => x"C0C0C0C082B082F9",
  6362 => x"C0C0C0C082B082A4",
  6363 => x"C0C0C0C082B082B0",
  6364 => x"C0C0C0C082B08299",
  6365 => x"C0C0C0C082B08292",
  6366 => x"C0C0C0C082B08282",
  6367 => x"C0C0C0C082B082F8",
  6368 => x"C0C0C0C082B08280",
  6369 => x"C0C0C0C082B08290",
  6370 => x"C0C0C0C082B0F8C0",
  6371 => x"C0C0C0C082B0F8F9",
  6372 => x"C0C0C0C082B0F8A4",
  6373 => x"C0C0C0C082B0F8B0",
  6374 => x"C0C0C0C082B0F899",
  6375 => x"C0C0C0C082B0F892",
  6376 => x"C0C0C0C082B0F882",
  6377 => x"C0C0C0C082B0F8F8",
  6378 => x"C0C0C0C082B0F880",
  6379 => x"C0C0C0C082B0F890",
  6380 => x"C0C0C0C082B080C0",
  6381 => x"C0C0C0C082B080F9",
  6382 => x"C0C0C0C082B080A4",
  6383 => x"C0C0C0C082B080B0",
  6384 => x"C0C0C0C082B08099",
  6385 => x"C0C0C0C082B08092",
  6386 => x"C0C0C0C082B08082",
  6387 => x"C0C0C0C082B080F8",
  6388 => x"C0C0C0C082B08080",
  6389 => x"C0C0C0C082B08090",
  6390 => x"C0C0C0C082B090C0",
  6391 => x"C0C0C0C082B090F9",
  6392 => x"C0C0C0C082B090A4",
  6393 => x"C0C0C0C082B090B0",
  6394 => x"C0C0C0C082B09099",
  6395 => x"C0C0C0C082B09092",
  6396 => x"C0C0C0C082B09082",
  6397 => x"C0C0C0C082B090F8",
  6398 => x"C0C0C0C082B09080",
  6399 => x"C0C0C0C082B09090",
  6400 => x"C0C0C0C08299C0C0",
  6401 => x"C0C0C0C08299C0F9",
  6402 => x"C0C0C0C08299C0A4",
  6403 => x"C0C0C0C08299C0B0",
  6404 => x"C0C0C0C08299C099",
  6405 => x"C0C0C0C08299C092",
  6406 => x"C0C0C0C08299C082",
  6407 => x"C0C0C0C08299C0F8",
  6408 => x"C0C0C0C08299C080",
  6409 => x"C0C0C0C08299C090",
  6410 => x"C0C0C0C08299F9C0",
  6411 => x"C0C0C0C08299F9F9",
  6412 => x"C0C0C0C08299F9A4",
  6413 => x"C0C0C0C08299F9B0",
  6414 => x"C0C0C0C08299F999",
  6415 => x"C0C0C0C08299F992",
  6416 => x"C0C0C0C08299F982",
  6417 => x"C0C0C0C08299F9F8",
  6418 => x"C0C0C0C08299F980",
  6419 => x"C0C0C0C08299F990",
  6420 => x"C0C0C0C08299A4C0",
  6421 => x"C0C0C0C08299A4F9",
  6422 => x"C0C0C0C08299A4A4",
  6423 => x"C0C0C0C08299A4B0",
  6424 => x"C0C0C0C08299A499",
  6425 => x"C0C0C0C08299A492",
  6426 => x"C0C0C0C08299A482",
  6427 => x"C0C0C0C08299A4F8",
  6428 => x"C0C0C0C08299A480",
  6429 => x"C0C0C0C08299A490",
  6430 => x"C0C0C0C08299B0C0",
  6431 => x"C0C0C0C08299B0F9",
  6432 => x"C0C0C0C08299B0A4",
  6433 => x"C0C0C0C08299B0B0",
  6434 => x"C0C0C0C08299B099",
  6435 => x"C0C0C0C08299B092",
  6436 => x"C0C0C0C08299B082",
  6437 => x"C0C0C0C08299B0F8",
  6438 => x"C0C0C0C08299B080",
  6439 => x"C0C0C0C08299B090",
  6440 => x"C0C0C0C0829999C0",
  6441 => x"C0C0C0C0829999F9",
  6442 => x"C0C0C0C0829999A4",
  6443 => x"C0C0C0C0829999B0",
  6444 => x"C0C0C0C082999999",
  6445 => x"C0C0C0C082999992",
  6446 => x"C0C0C0C082999982",
  6447 => x"C0C0C0C0829999F8",
  6448 => x"C0C0C0C082999980",
  6449 => x"C0C0C0C082999990",
  6450 => x"C0C0C0C0829992C0",
  6451 => x"C0C0C0C0829992F9",
  6452 => x"C0C0C0C0829992A4",
  6453 => x"C0C0C0C0829992B0",
  6454 => x"C0C0C0C082999299",
  6455 => x"C0C0C0C082999292",
  6456 => x"C0C0C0C082999282",
  6457 => x"C0C0C0C0829992F8",
  6458 => x"C0C0C0C082999280",
  6459 => x"C0C0C0C082999290",
  6460 => x"C0C0C0C0829982C0",
  6461 => x"C0C0C0C0829982F9",
  6462 => x"C0C0C0C0829982A4",
  6463 => x"C0C0C0C0829982B0",
  6464 => x"C0C0C0C082998299",
  6465 => x"C0C0C0C082998292",
  6466 => x"C0C0C0C082998282",
  6467 => x"C0C0C0C0829982F8",
  6468 => x"C0C0C0C082998280",
  6469 => x"C0C0C0C082998290",
  6470 => x"C0C0C0C08299F8C0",
  6471 => x"C0C0C0C08299F8F9",
  6472 => x"C0C0C0C08299F8A4",
  6473 => x"C0C0C0C08299F8B0",
  6474 => x"C0C0C0C08299F899",
  6475 => x"C0C0C0C08299F892",
  6476 => x"C0C0C0C08299F882",
  6477 => x"C0C0C0C08299F8F8",
  6478 => x"C0C0C0C08299F880",
  6479 => x"C0C0C0C08299F890",
  6480 => x"C0C0C0C0829980C0",
  6481 => x"C0C0C0C0829980F9",
  6482 => x"C0C0C0C0829980A4",
  6483 => x"C0C0C0C0829980B0",
  6484 => x"C0C0C0C082998099",
  6485 => x"C0C0C0C082998092",
  6486 => x"C0C0C0C082998082",
  6487 => x"C0C0C0C0829980F8",
  6488 => x"C0C0C0C082998080",
  6489 => x"C0C0C0C082998090",
  6490 => x"C0C0C0C0829990C0",
  6491 => x"C0C0C0C0829990F9",
  6492 => x"C0C0C0C0829990A4",
  6493 => x"C0C0C0C0829990B0",
  6494 => x"C0C0C0C082999099",
  6495 => x"C0C0C0C082999092",
  6496 => x"C0C0C0C082999082",
  6497 => x"C0C0C0C0829990F8",
  6498 => x"C0C0C0C082999080",
  6499 => x"C0C0C0C082999090",
  6500 => x"C0C0C0C08292C0C0",
  6501 => x"C0C0C0C08292C0F9",
  6502 => x"C0C0C0C08292C0A4",
  6503 => x"C0C0C0C08292C0B0",
  6504 => x"C0C0C0C08292C099",
  6505 => x"C0C0C0C08292C092",
  6506 => x"C0C0C0C08292C082",
  6507 => x"C0C0C0C08292C0F8",
  6508 => x"C0C0C0C08292C080",
  6509 => x"C0C0C0C08292C090",
  6510 => x"C0C0C0C08292F9C0",
  6511 => x"C0C0C0C08292F9F9",
  6512 => x"C0C0C0C08292F9A4",
  6513 => x"C0C0C0C08292F9B0",
  6514 => x"C0C0C0C08292F999",
  6515 => x"C0C0C0C08292F992",
  6516 => x"C0C0C0C08292F982",
  6517 => x"C0C0C0C08292F9F8",
  6518 => x"C0C0C0C08292F980",
  6519 => x"C0C0C0C08292F990",
  6520 => x"C0C0C0C08292A4C0",
  6521 => x"C0C0C0C08292A4F9",
  6522 => x"C0C0C0C08292A4A4",
  6523 => x"C0C0C0C08292A4B0",
  6524 => x"C0C0C0C08292A499",
  6525 => x"C0C0C0C08292A492",
  6526 => x"C0C0C0C08292A482",
  6527 => x"C0C0C0C08292A4F8",
  6528 => x"C0C0C0C08292A480",
  6529 => x"C0C0C0C08292A490",
  6530 => x"C0C0C0C08292B0C0",
  6531 => x"C0C0C0C08292B0F9",
  6532 => x"C0C0C0C08292B0A4",
  6533 => x"C0C0C0C08292B0B0",
  6534 => x"C0C0C0C08292B099",
  6535 => x"C0C0C0C08292B092",
  6536 => x"C0C0C0C08292B082",
  6537 => x"C0C0C0C08292B0F8",
  6538 => x"C0C0C0C08292B080",
  6539 => x"C0C0C0C08292B090",
  6540 => x"C0C0C0C0829299C0",
  6541 => x"C0C0C0C0829299F9",
  6542 => x"C0C0C0C0829299A4",
  6543 => x"C0C0C0C0829299B0",
  6544 => x"C0C0C0C082929999",
  6545 => x"C0C0C0C082929992",
  6546 => x"C0C0C0C082929982",
  6547 => x"C0C0C0C0829299F8",
  6548 => x"C0C0C0C082929980",
  6549 => x"C0C0C0C082929990",
  6550 => x"C0C0C0C0829292C0",
  6551 => x"C0C0C0C0829292F9",
  6552 => x"C0C0C0C0829292A4",
  6553 => x"C0C0C0C0829292B0",
  6554 => x"C0C0C0C082929299",
  6555 => x"C0C0C0C082929292",
  6556 => x"C0C0C0C082929282",
  6557 => x"C0C0C0C0829292F8",
  6558 => x"C0C0C0C082929280",
  6559 => x"C0C0C0C082929290",
  6560 => x"C0C0C0C0829282C0",
  6561 => x"C0C0C0C0829282F9",
  6562 => x"C0C0C0C0829282A4",
  6563 => x"C0C0C0C0829282B0",
  6564 => x"C0C0C0C082928299",
  6565 => x"C0C0C0C082928292",
  6566 => x"C0C0C0C082928282",
  6567 => x"C0C0C0C0829282F8",
  6568 => x"C0C0C0C082928280",
  6569 => x"C0C0C0C082928290",
  6570 => x"C0C0C0C08292F8C0",
  6571 => x"C0C0C0C08292F8F9",
  6572 => x"C0C0C0C08292F8A4",
  6573 => x"C0C0C0C08292F8B0",
  6574 => x"C0C0C0C08292F899",
  6575 => x"C0C0C0C08292F892",
  6576 => x"C0C0C0C08292F882",
  6577 => x"C0C0C0C08292F8F8",
  6578 => x"C0C0C0C08292F880",
  6579 => x"C0C0C0C08292F890",
  6580 => x"C0C0C0C0829280C0",
  6581 => x"C0C0C0C0829280F9",
  6582 => x"C0C0C0C0829280A4",
  6583 => x"C0C0C0C0829280B0",
  6584 => x"C0C0C0C082928099",
  6585 => x"C0C0C0C082928092",
  6586 => x"C0C0C0C082928082",
  6587 => x"C0C0C0C0829280F8",
  6588 => x"C0C0C0C082928080",
  6589 => x"C0C0C0C082928090",
  6590 => x"C0C0C0C0829290C0",
  6591 => x"C0C0C0C0829290F9",
  6592 => x"C0C0C0C0829290A4",
  6593 => x"C0C0C0C0829290B0",
  6594 => x"C0C0C0C082929099",
  6595 => x"C0C0C0C082929092",
  6596 => x"C0C0C0C082929082",
  6597 => x"C0C0C0C0829290F8",
  6598 => x"C0C0C0C082929080",
  6599 => x"C0C0C0C082929090",
  6600 => x"C0C0C0C08282C0C0",
  6601 => x"C0C0C0C08282C0F9",
  6602 => x"C0C0C0C08282C0A4",
  6603 => x"C0C0C0C08282C0B0",
  6604 => x"C0C0C0C08282C099",
  6605 => x"C0C0C0C08282C092",
  6606 => x"C0C0C0C08282C082",
  6607 => x"C0C0C0C08282C0F8",
  6608 => x"C0C0C0C08282C080",
  6609 => x"C0C0C0C08282C090",
  6610 => x"C0C0C0C08282F9C0",
  6611 => x"C0C0C0C08282F9F9",
  6612 => x"C0C0C0C08282F9A4",
  6613 => x"C0C0C0C08282F9B0",
  6614 => x"C0C0C0C08282F999",
  6615 => x"C0C0C0C08282F992",
  6616 => x"C0C0C0C08282F982",
  6617 => x"C0C0C0C08282F9F8",
  6618 => x"C0C0C0C08282F980",
  6619 => x"C0C0C0C08282F990",
  6620 => x"C0C0C0C08282A4C0",
  6621 => x"C0C0C0C08282A4F9",
  6622 => x"C0C0C0C08282A4A4",
  6623 => x"C0C0C0C08282A4B0",
  6624 => x"C0C0C0C08282A499",
  6625 => x"C0C0C0C08282A492",
  6626 => x"C0C0C0C08282A482",
  6627 => x"C0C0C0C08282A4F8",
  6628 => x"C0C0C0C08282A480",
  6629 => x"C0C0C0C08282A490",
  6630 => x"C0C0C0C08282B0C0",
  6631 => x"C0C0C0C08282B0F9",
  6632 => x"C0C0C0C08282B0A4",
  6633 => x"C0C0C0C08282B0B0",
  6634 => x"C0C0C0C08282B099",
  6635 => x"C0C0C0C08282B092",
  6636 => x"C0C0C0C08282B082",
  6637 => x"C0C0C0C08282B0F8",
  6638 => x"C0C0C0C08282B080",
  6639 => x"C0C0C0C08282B090",
  6640 => x"C0C0C0C0828299C0",
  6641 => x"C0C0C0C0828299F9",
  6642 => x"C0C0C0C0828299A4",
  6643 => x"C0C0C0C0828299B0",
  6644 => x"C0C0C0C082829999",
  6645 => x"C0C0C0C082829992",
  6646 => x"C0C0C0C082829982",
  6647 => x"C0C0C0C0828299F8",
  6648 => x"C0C0C0C082829980",
  6649 => x"C0C0C0C082829990",
  6650 => x"C0C0C0C0828292C0",
  6651 => x"C0C0C0C0828292F9",
  6652 => x"C0C0C0C0828292A4",
  6653 => x"C0C0C0C0828292B0",
  6654 => x"C0C0C0C082829299",
  6655 => x"C0C0C0C082829292",
  6656 => x"C0C0C0C082829282",
  6657 => x"C0C0C0C0828292F8",
  6658 => x"C0C0C0C082829280",
  6659 => x"C0C0C0C082829290",
  6660 => x"C0C0C0C0828282C0",
  6661 => x"C0C0C0C0828282F9",
  6662 => x"C0C0C0C0828282A4",
  6663 => x"C0C0C0C0828282B0",
  6664 => x"C0C0C0C082828299",
  6665 => x"C0C0C0C082828292",
  6666 => x"C0C0C0C082828282",
  6667 => x"C0C0C0C0828282F8",
  6668 => x"C0C0C0C082828280",
  6669 => x"C0C0C0C082828290",
  6670 => x"C0C0C0C08282F8C0",
  6671 => x"C0C0C0C08282F8F9",
  6672 => x"C0C0C0C08282F8A4",
  6673 => x"C0C0C0C08282F8B0",
  6674 => x"C0C0C0C08282F899",
  6675 => x"C0C0C0C08282F892",
  6676 => x"C0C0C0C08282F882",
  6677 => x"C0C0C0C08282F8F8",
  6678 => x"C0C0C0C08282F880",
  6679 => x"C0C0C0C08282F890",
  6680 => x"C0C0C0C0828280C0",
  6681 => x"C0C0C0C0828280F9",
  6682 => x"C0C0C0C0828280A4",
  6683 => x"C0C0C0C0828280B0",
  6684 => x"C0C0C0C082828099",
  6685 => x"C0C0C0C082828092",
  6686 => x"C0C0C0C082828082",
  6687 => x"C0C0C0C0828280F8",
  6688 => x"C0C0C0C082828080",
  6689 => x"C0C0C0C082828090",
  6690 => x"C0C0C0C0828290C0",
  6691 => x"C0C0C0C0828290F9",
  6692 => x"C0C0C0C0828290A4",
  6693 => x"C0C0C0C0828290B0",
  6694 => x"C0C0C0C082829099",
  6695 => x"C0C0C0C082829092",
  6696 => x"C0C0C0C082829082",
  6697 => x"C0C0C0C0828290F8",
  6698 => x"C0C0C0C082829080",
  6699 => x"C0C0C0C082829090",
  6700 => x"C0C0C0C082F8C0C0",
  6701 => x"C0C0C0C082F8C0F9",
  6702 => x"C0C0C0C082F8C0A4",
  6703 => x"C0C0C0C082F8C0B0",
  6704 => x"C0C0C0C082F8C099",
  6705 => x"C0C0C0C082F8C092",
  6706 => x"C0C0C0C082F8C082",
  6707 => x"C0C0C0C082F8C0F8",
  6708 => x"C0C0C0C082F8C080",
  6709 => x"C0C0C0C082F8C090",
  6710 => x"C0C0C0C082F8F9C0",
  6711 => x"C0C0C0C082F8F9F9",
  6712 => x"C0C0C0C082F8F9A4",
  6713 => x"C0C0C0C082F8F9B0",
  6714 => x"C0C0C0C082F8F999",
  6715 => x"C0C0C0C082F8F992",
  6716 => x"C0C0C0C082F8F982",
  6717 => x"C0C0C0C082F8F9F8",
  6718 => x"C0C0C0C082F8F980",
  6719 => x"C0C0C0C082F8F990",
  6720 => x"C0C0C0C082F8A4C0",
  6721 => x"C0C0C0C082F8A4F9",
  6722 => x"C0C0C0C082F8A4A4",
  6723 => x"C0C0C0C082F8A4B0",
  6724 => x"C0C0C0C082F8A499",
  6725 => x"C0C0C0C082F8A492",
  6726 => x"C0C0C0C082F8A482",
  6727 => x"C0C0C0C082F8A4F8",
  6728 => x"C0C0C0C082F8A480",
  6729 => x"C0C0C0C082F8A490",
  6730 => x"C0C0C0C082F8B0C0",
  6731 => x"C0C0C0C082F8B0F9",
  6732 => x"C0C0C0C082F8B0A4",
  6733 => x"C0C0C0C082F8B0B0",
  6734 => x"C0C0C0C082F8B099",
  6735 => x"C0C0C0C082F8B092",
  6736 => x"C0C0C0C082F8B082",
  6737 => x"C0C0C0C082F8B0F8",
  6738 => x"C0C0C0C082F8B080",
  6739 => x"C0C0C0C082F8B090",
  6740 => x"C0C0C0C082F899C0",
  6741 => x"C0C0C0C082F899F9",
  6742 => x"C0C0C0C082F899A4",
  6743 => x"C0C0C0C082F899B0",
  6744 => x"C0C0C0C082F89999",
  6745 => x"C0C0C0C082F89992",
  6746 => x"C0C0C0C082F89982",
  6747 => x"C0C0C0C082F899F8",
  6748 => x"C0C0C0C082F89980",
  6749 => x"C0C0C0C082F89990",
  6750 => x"C0C0C0C082F892C0",
  6751 => x"C0C0C0C082F892F9",
  6752 => x"C0C0C0C082F892A4",
  6753 => x"C0C0C0C082F892B0",
  6754 => x"C0C0C0C082F89299",
  6755 => x"C0C0C0C082F89292",
  6756 => x"C0C0C0C082F89282",
  6757 => x"C0C0C0C082F892F8",
  6758 => x"C0C0C0C082F89280",
  6759 => x"C0C0C0C082F89290",
  6760 => x"C0C0C0C082F882C0",
  6761 => x"C0C0C0C082F882F9",
  6762 => x"C0C0C0C082F882A4",
  6763 => x"C0C0C0C082F882B0",
  6764 => x"C0C0C0C082F88299",
  6765 => x"C0C0C0C082F88292",
  6766 => x"C0C0C0C082F88282",
  6767 => x"C0C0C0C082F882F8",
  6768 => x"C0C0C0C082F88280",
  6769 => x"C0C0C0C082F88290",
  6770 => x"C0C0C0C082F8F8C0",
  6771 => x"C0C0C0C082F8F8F9",
  6772 => x"C0C0C0C082F8F8A4",
  6773 => x"C0C0C0C082F8F8B0",
  6774 => x"C0C0C0C082F8F899",
  6775 => x"C0C0C0C082F8F892",
  6776 => x"C0C0C0C082F8F882",
  6777 => x"C0C0C0C082F8F8F8",
  6778 => x"C0C0C0C082F8F880",
  6779 => x"C0C0C0C082F8F890",
  6780 => x"C0C0C0C082F880C0",
  6781 => x"C0C0C0C082F880F9",
  6782 => x"C0C0C0C082F880A4",
  6783 => x"C0C0C0C082F880B0",
  6784 => x"C0C0C0C082F88099",
  6785 => x"C0C0C0C082F88092",
  6786 => x"C0C0C0C082F88082",
  6787 => x"C0C0C0C082F880F8",
  6788 => x"C0C0C0C082F88080",
  6789 => x"C0C0C0C082F88090",
  6790 => x"C0C0C0C082F890C0",
  6791 => x"C0C0C0C082F890F9",
  6792 => x"C0C0C0C082F890A4",
  6793 => x"C0C0C0C082F890B0",
  6794 => x"C0C0C0C082F89099",
  6795 => x"C0C0C0C082F89092",
  6796 => x"C0C0C0C082F89082",
  6797 => x"C0C0C0C082F890F8",
  6798 => x"C0C0C0C082F89080",
  6799 => x"C0C0C0C082F89090",
  6800 => x"C0C0C0C08280C0C0",
  6801 => x"C0C0C0C08280C0F9",
  6802 => x"C0C0C0C08280C0A4",
  6803 => x"C0C0C0C08280C0B0",
  6804 => x"C0C0C0C08280C099",
  6805 => x"C0C0C0C08280C092",
  6806 => x"C0C0C0C08280C082",
  6807 => x"C0C0C0C08280C0F8",
  6808 => x"C0C0C0C08280C080",
  6809 => x"C0C0C0C08280C090",
  6810 => x"C0C0C0C08280F9C0",
  6811 => x"C0C0C0C08280F9F9",
  6812 => x"C0C0C0C08280F9A4",
  6813 => x"C0C0C0C08280F9B0",
  6814 => x"C0C0C0C08280F999",
  6815 => x"C0C0C0C08280F992",
  6816 => x"C0C0C0C08280F982",
  6817 => x"C0C0C0C08280F9F8",
  6818 => x"C0C0C0C08280F980",
  6819 => x"C0C0C0C08280F990",
  6820 => x"C0C0C0C08280A4C0",
  6821 => x"C0C0C0C08280A4F9",
  6822 => x"C0C0C0C08280A4A4",
  6823 => x"C0C0C0C08280A4B0",
  6824 => x"C0C0C0C08280A499",
  6825 => x"C0C0C0C08280A492",
  6826 => x"C0C0C0C08280A482",
  6827 => x"C0C0C0C08280A4F8",
  6828 => x"C0C0C0C08280A480",
  6829 => x"C0C0C0C08280A490",
  6830 => x"C0C0C0C08280B0C0",
  6831 => x"C0C0C0C08280B0F9",
  6832 => x"C0C0C0C08280B0A4",
  6833 => x"C0C0C0C08280B0B0",
  6834 => x"C0C0C0C08280B099",
  6835 => x"C0C0C0C08280B092",
  6836 => x"C0C0C0C08280B082",
  6837 => x"C0C0C0C08280B0F8",
  6838 => x"C0C0C0C08280B080",
  6839 => x"C0C0C0C08280B090",
  6840 => x"C0C0C0C0828099C0",
  6841 => x"C0C0C0C0828099F9",
  6842 => x"C0C0C0C0828099A4",
  6843 => x"C0C0C0C0828099B0",
  6844 => x"C0C0C0C082809999",
  6845 => x"C0C0C0C082809992",
  6846 => x"C0C0C0C082809982",
  6847 => x"C0C0C0C0828099F8",
  6848 => x"C0C0C0C082809980",
  6849 => x"C0C0C0C082809990",
  6850 => x"C0C0C0C0828092C0",
  6851 => x"C0C0C0C0828092F9",
  6852 => x"C0C0C0C0828092A4",
  6853 => x"C0C0C0C0828092B0",
  6854 => x"C0C0C0C082809299",
  6855 => x"C0C0C0C082809292",
  6856 => x"C0C0C0C082809282",
  6857 => x"C0C0C0C0828092F8",
  6858 => x"C0C0C0C082809280",
  6859 => x"C0C0C0C082809290",
  6860 => x"C0C0C0C0828082C0",
  6861 => x"C0C0C0C0828082F9",
  6862 => x"C0C0C0C0828082A4",
  6863 => x"C0C0C0C0828082B0",
  6864 => x"C0C0C0C082808299",
  6865 => x"C0C0C0C082808292",
  6866 => x"C0C0C0C082808282",
  6867 => x"C0C0C0C0828082F8",
  6868 => x"C0C0C0C082808280",
  6869 => x"C0C0C0C082808290",
  6870 => x"C0C0C0C08280F8C0",
  6871 => x"C0C0C0C08280F8F9",
  6872 => x"C0C0C0C08280F8A4",
  6873 => x"C0C0C0C08280F8B0",
  6874 => x"C0C0C0C08280F899",
  6875 => x"C0C0C0C08280F892",
  6876 => x"C0C0C0C08280F882",
  6877 => x"C0C0C0C08280F8F8",
  6878 => x"C0C0C0C08280F880",
  6879 => x"C0C0C0C08280F890",
  6880 => x"C0C0C0C0828080C0",
  6881 => x"C0C0C0C0828080F9",
  6882 => x"C0C0C0C0828080A4",
  6883 => x"C0C0C0C0828080B0",
  6884 => x"C0C0C0C082808099",
  6885 => x"C0C0C0C082808092",
  6886 => x"C0C0C0C082808082",
  6887 => x"C0C0C0C0828080F8",
  6888 => x"C0C0C0C082808080",
  6889 => x"C0C0C0C082808090",
  6890 => x"C0C0C0C0828090C0",
  6891 => x"C0C0C0C0828090F9",
  6892 => x"C0C0C0C0828090A4",
  6893 => x"C0C0C0C0828090B0",
  6894 => x"C0C0C0C082809099",
  6895 => x"C0C0C0C082809092",
  6896 => x"C0C0C0C082809082",
  6897 => x"C0C0C0C0828090F8",
  6898 => x"C0C0C0C082809080",
  6899 => x"C0C0C0C082809090",
  6900 => x"C0C0C0C08290C0C0",
  6901 => x"C0C0C0C08290C0F9",
  6902 => x"C0C0C0C08290C0A4",
  6903 => x"C0C0C0C08290C0B0",
  6904 => x"C0C0C0C08290C099",
  6905 => x"C0C0C0C08290C092",
  6906 => x"C0C0C0C08290C082",
  6907 => x"C0C0C0C08290C0F8",
  6908 => x"C0C0C0C08290C080",
  6909 => x"C0C0C0C08290C090",
  6910 => x"C0C0C0C08290F9C0",
  6911 => x"C0C0C0C08290F9F9",
  6912 => x"C0C0C0C08290F9A4",
  6913 => x"C0C0C0C08290F9B0",
  6914 => x"C0C0C0C08290F999",
  6915 => x"C0C0C0C08290F992",
  6916 => x"C0C0C0C08290F982",
  6917 => x"C0C0C0C08290F9F8",
  6918 => x"C0C0C0C08290F980",
  6919 => x"C0C0C0C08290F990",
  6920 => x"C0C0C0C08290A4C0",
  6921 => x"C0C0C0C08290A4F9",
  6922 => x"C0C0C0C08290A4A4",
  6923 => x"C0C0C0C08290A4B0",
  6924 => x"C0C0C0C08290A499",
  6925 => x"C0C0C0C08290A492",
  6926 => x"C0C0C0C08290A482",
  6927 => x"C0C0C0C08290A4F8",
  6928 => x"C0C0C0C08290A480",
  6929 => x"C0C0C0C08290A490",
  6930 => x"C0C0C0C08290B0C0",
  6931 => x"C0C0C0C08290B0F9",
  6932 => x"C0C0C0C08290B0A4",
  6933 => x"C0C0C0C08290B0B0",
  6934 => x"C0C0C0C08290B099",
  6935 => x"C0C0C0C08290B092",
  6936 => x"C0C0C0C08290B082",
  6937 => x"C0C0C0C08290B0F8",
  6938 => x"C0C0C0C08290B080",
  6939 => x"C0C0C0C08290B090",
  6940 => x"C0C0C0C0829099C0",
  6941 => x"C0C0C0C0829099F9",
  6942 => x"C0C0C0C0829099A4",
  6943 => x"C0C0C0C0829099B0",
  6944 => x"C0C0C0C082909999",
  6945 => x"C0C0C0C082909992",
  6946 => x"C0C0C0C082909982",
  6947 => x"C0C0C0C0829099F8",
  6948 => x"C0C0C0C082909980",
  6949 => x"C0C0C0C082909990",
  6950 => x"C0C0C0C0829092C0",
  6951 => x"C0C0C0C0829092F9",
  6952 => x"C0C0C0C0829092A4",
  6953 => x"C0C0C0C0829092B0",
  6954 => x"C0C0C0C082909299",
  6955 => x"C0C0C0C082909292",
  6956 => x"C0C0C0C082909282",
  6957 => x"C0C0C0C0829092F8",
  6958 => x"C0C0C0C082909280",
  6959 => x"C0C0C0C082909290",
  6960 => x"C0C0C0C0829082C0",
  6961 => x"C0C0C0C0829082F9",
  6962 => x"C0C0C0C0829082A4",
  6963 => x"C0C0C0C0829082B0",
  6964 => x"C0C0C0C082908299",
  6965 => x"C0C0C0C082908292",
  6966 => x"C0C0C0C082908282",
  6967 => x"C0C0C0C0829082F8",
  6968 => x"C0C0C0C082908280",
  6969 => x"C0C0C0C082908290",
  6970 => x"C0C0C0C08290F8C0",
  6971 => x"C0C0C0C08290F8F9",
  6972 => x"C0C0C0C08290F8A4",
  6973 => x"C0C0C0C08290F8B0",
  6974 => x"C0C0C0C08290F899",
  6975 => x"C0C0C0C08290F892",
  6976 => x"C0C0C0C08290F882",
  6977 => x"C0C0C0C08290F8F8",
  6978 => x"C0C0C0C08290F880",
  6979 => x"C0C0C0C08290F890",
  6980 => x"C0C0C0C0829080C0",
  6981 => x"C0C0C0C0829080F9",
  6982 => x"C0C0C0C0829080A4",
  6983 => x"C0C0C0C0829080B0",
  6984 => x"C0C0C0C082908099",
  6985 => x"C0C0C0C082908092",
  6986 => x"C0C0C0C082908082",
  6987 => x"C0C0C0C0829080F8",
  6988 => x"C0C0C0C082908080",
  6989 => x"C0C0C0C082908090",
  6990 => x"C0C0C0C0829090C0",
  6991 => x"C0C0C0C0829090F9",
  6992 => x"C0C0C0C0829090A4",
  6993 => x"C0C0C0C0829090B0",
  6994 => x"C0C0C0C082909099",
  6995 => x"C0C0C0C082909092",
  6996 => x"C0C0C0C082909082",
  6997 => x"C0C0C0C0829090F8",
  6998 => x"C0C0C0C082909080",
  6999 => x"C0C0C0C082909090",
  7000 => x"C0C0C0C0F8C0C0C0",
  7001 => x"C0C0C0C0F8C0C0F9",
  7002 => x"C0C0C0C0F8C0C0A4",
  7003 => x"C0C0C0C0F8C0C0B0",
  7004 => x"C0C0C0C0F8C0C099",
  7005 => x"C0C0C0C0F8C0C092",
  7006 => x"C0C0C0C0F8C0C082",
  7007 => x"C0C0C0C0F8C0C0F8",
  7008 => x"C0C0C0C0F8C0C080",
  7009 => x"C0C0C0C0F8C0C090",
  7010 => x"C0C0C0C0F8C0F9C0",
  7011 => x"C0C0C0C0F8C0F9F9",
  7012 => x"C0C0C0C0F8C0F9A4",
  7013 => x"C0C0C0C0F8C0F9B0",
  7014 => x"C0C0C0C0F8C0F999",
  7015 => x"C0C0C0C0F8C0F992",
  7016 => x"C0C0C0C0F8C0F982",
  7017 => x"C0C0C0C0F8C0F9F8",
  7018 => x"C0C0C0C0F8C0F980",
  7019 => x"C0C0C0C0F8C0F990",
  7020 => x"C0C0C0C0F8C0A4C0",
  7021 => x"C0C0C0C0F8C0A4F9",
  7022 => x"C0C0C0C0F8C0A4A4",
  7023 => x"C0C0C0C0F8C0A4B0",
  7024 => x"C0C0C0C0F8C0A499",
  7025 => x"C0C0C0C0F8C0A492",
  7026 => x"C0C0C0C0F8C0A482",
  7027 => x"C0C0C0C0F8C0A4F8",
  7028 => x"C0C0C0C0F8C0A480",
  7029 => x"C0C0C0C0F8C0A490",
  7030 => x"C0C0C0C0F8C0B0C0",
  7031 => x"C0C0C0C0F8C0B0F9",
  7032 => x"C0C0C0C0F8C0B0A4",
  7033 => x"C0C0C0C0F8C0B0B0",
  7034 => x"C0C0C0C0F8C0B099",
  7035 => x"C0C0C0C0F8C0B092",
  7036 => x"C0C0C0C0F8C0B082",
  7037 => x"C0C0C0C0F8C0B0F8",
  7038 => x"C0C0C0C0F8C0B080",
  7039 => x"C0C0C0C0F8C0B090",
  7040 => x"C0C0C0C0F8C099C0",
  7041 => x"C0C0C0C0F8C099F9",
  7042 => x"C0C0C0C0F8C099A4",
  7043 => x"C0C0C0C0F8C099B0",
  7044 => x"C0C0C0C0F8C09999",
  7045 => x"C0C0C0C0F8C09992",
  7046 => x"C0C0C0C0F8C09982",
  7047 => x"C0C0C0C0F8C099F8",
  7048 => x"C0C0C0C0F8C09980",
  7049 => x"C0C0C0C0F8C09990",
  7050 => x"C0C0C0C0F8C092C0",
  7051 => x"C0C0C0C0F8C092F9",
  7052 => x"C0C0C0C0F8C092A4",
  7053 => x"C0C0C0C0F8C092B0",
  7054 => x"C0C0C0C0F8C09299",
  7055 => x"C0C0C0C0F8C09292",
  7056 => x"C0C0C0C0F8C09282",
  7057 => x"C0C0C0C0F8C092F8",
  7058 => x"C0C0C0C0F8C09280",
  7059 => x"C0C0C0C0F8C09290",
  7060 => x"C0C0C0C0F8C082C0",
  7061 => x"C0C0C0C0F8C082F9",
  7062 => x"C0C0C0C0F8C082A4",
  7063 => x"C0C0C0C0F8C082B0",
  7064 => x"C0C0C0C0F8C08299",
  7065 => x"C0C0C0C0F8C08292",
  7066 => x"C0C0C0C0F8C08282",
  7067 => x"C0C0C0C0F8C082F8",
  7068 => x"C0C0C0C0F8C08280",
  7069 => x"C0C0C0C0F8C08290",
  7070 => x"C0C0C0C0F8C0F8C0",
  7071 => x"C0C0C0C0F8C0F8F9",
  7072 => x"C0C0C0C0F8C0F8A4",
  7073 => x"C0C0C0C0F8C0F8B0",
  7074 => x"C0C0C0C0F8C0F899",
  7075 => x"C0C0C0C0F8C0F892",
  7076 => x"C0C0C0C0F8C0F882",
  7077 => x"C0C0C0C0F8C0F8F8",
  7078 => x"C0C0C0C0F8C0F880",
  7079 => x"C0C0C0C0F8C0F890",
  7080 => x"C0C0C0C0F8C080C0",
  7081 => x"C0C0C0C0F8C080F9",
  7082 => x"C0C0C0C0F8C080A4",
  7083 => x"C0C0C0C0F8C080B0",
  7084 => x"C0C0C0C0F8C08099",
  7085 => x"C0C0C0C0F8C08092",
  7086 => x"C0C0C0C0F8C08082",
  7087 => x"C0C0C0C0F8C080F8",
  7088 => x"C0C0C0C0F8C08080",
  7089 => x"C0C0C0C0F8C08090",
  7090 => x"C0C0C0C0F8C090C0",
  7091 => x"C0C0C0C0F8C090F9",
  7092 => x"C0C0C0C0F8C090A4",
  7093 => x"C0C0C0C0F8C090B0",
  7094 => x"C0C0C0C0F8C09099",
  7095 => x"C0C0C0C0F8C09092",
  7096 => x"C0C0C0C0F8C09082",
  7097 => x"C0C0C0C0F8C090F8",
  7098 => x"C0C0C0C0F8C09080",
  7099 => x"C0C0C0C0F8C09090",
  7100 => x"C0C0C0C0F8F9C0C0",
  7101 => x"C0C0C0C0F8F9C0F9",
  7102 => x"C0C0C0C0F8F9C0A4",
  7103 => x"C0C0C0C0F8F9C0B0",
  7104 => x"C0C0C0C0F8F9C099",
  7105 => x"C0C0C0C0F8F9C092",
  7106 => x"C0C0C0C0F8F9C082",
  7107 => x"C0C0C0C0F8F9C0F8",
  7108 => x"C0C0C0C0F8F9C080",
  7109 => x"C0C0C0C0F8F9C090",
  7110 => x"C0C0C0C0F8F9F9C0",
  7111 => x"C0C0C0C0F8F9F9F9",
  7112 => x"C0C0C0C0F8F9F9A4",
  7113 => x"C0C0C0C0F8F9F9B0",
  7114 => x"C0C0C0C0F8F9F999",
  7115 => x"C0C0C0C0F8F9F992",
  7116 => x"C0C0C0C0F8F9F982",
  7117 => x"C0C0C0C0F8F9F9F8",
  7118 => x"C0C0C0C0F8F9F980",
  7119 => x"C0C0C0C0F8F9F990",
  7120 => x"C0C0C0C0F8F9A4C0",
  7121 => x"C0C0C0C0F8F9A4F9",
  7122 => x"C0C0C0C0F8F9A4A4",
  7123 => x"C0C0C0C0F8F9A4B0",
  7124 => x"C0C0C0C0F8F9A499",
  7125 => x"C0C0C0C0F8F9A492",
  7126 => x"C0C0C0C0F8F9A482",
  7127 => x"C0C0C0C0F8F9A4F8",
  7128 => x"C0C0C0C0F8F9A480",
  7129 => x"C0C0C0C0F8F9A490",
  7130 => x"C0C0C0C0F8F9B0C0",
  7131 => x"C0C0C0C0F8F9B0F9",
  7132 => x"C0C0C0C0F8F9B0A4",
  7133 => x"C0C0C0C0F8F9B0B0",
  7134 => x"C0C0C0C0F8F9B099",
  7135 => x"C0C0C0C0F8F9B092",
  7136 => x"C0C0C0C0F8F9B082",
  7137 => x"C0C0C0C0F8F9B0F8",
  7138 => x"C0C0C0C0F8F9B080",
  7139 => x"C0C0C0C0F8F9B090",
  7140 => x"C0C0C0C0F8F999C0",
  7141 => x"C0C0C0C0F8F999F9",
  7142 => x"C0C0C0C0F8F999A4",
  7143 => x"C0C0C0C0F8F999B0",
  7144 => x"C0C0C0C0F8F99999",
  7145 => x"C0C0C0C0F8F99992",
  7146 => x"C0C0C0C0F8F99982",
  7147 => x"C0C0C0C0F8F999F8",
  7148 => x"C0C0C0C0F8F99980",
  7149 => x"C0C0C0C0F8F99990",
  7150 => x"C0C0C0C0F8F992C0",
  7151 => x"C0C0C0C0F8F992F9",
  7152 => x"C0C0C0C0F8F992A4",
  7153 => x"C0C0C0C0F8F992B0",
  7154 => x"C0C0C0C0F8F99299",
  7155 => x"C0C0C0C0F8F99292",
  7156 => x"C0C0C0C0F8F99282",
  7157 => x"C0C0C0C0F8F992F8",
  7158 => x"C0C0C0C0F8F99280",
  7159 => x"C0C0C0C0F8F99290",
  7160 => x"C0C0C0C0F8F982C0",
  7161 => x"C0C0C0C0F8F982F9",
  7162 => x"C0C0C0C0F8F982A4",
  7163 => x"C0C0C0C0F8F982B0",
  7164 => x"C0C0C0C0F8F98299",
  7165 => x"C0C0C0C0F8F98292",
  7166 => x"C0C0C0C0F8F98282",
  7167 => x"C0C0C0C0F8F982F8",
  7168 => x"C0C0C0C0F8F98280",
  7169 => x"C0C0C0C0F8F98290",
  7170 => x"C0C0C0C0F8F9F8C0",
  7171 => x"C0C0C0C0F8F9F8F9",
  7172 => x"C0C0C0C0F8F9F8A4",
  7173 => x"C0C0C0C0F8F9F8B0",
  7174 => x"C0C0C0C0F8F9F899",
  7175 => x"C0C0C0C0F8F9F892",
  7176 => x"C0C0C0C0F8F9F882",
  7177 => x"C0C0C0C0F8F9F8F8",
  7178 => x"C0C0C0C0F8F9F880",
  7179 => x"C0C0C0C0F8F9F890",
  7180 => x"C0C0C0C0F8F980C0",
  7181 => x"C0C0C0C0F8F980F9",
  7182 => x"C0C0C0C0F8F980A4",
  7183 => x"C0C0C0C0F8F980B0",
  7184 => x"C0C0C0C0F8F98099",
  7185 => x"C0C0C0C0F8F98092",
  7186 => x"C0C0C0C0F8F98082",
  7187 => x"C0C0C0C0F8F980F8",
  7188 => x"C0C0C0C0F8F98080",
  7189 => x"C0C0C0C0F8F98090",
  7190 => x"C0C0C0C0F8F990C0",
  7191 => x"C0C0C0C0F8F990F9",
  7192 => x"C0C0C0C0F8F990A4",
  7193 => x"C0C0C0C0F8F990B0",
  7194 => x"C0C0C0C0F8F99099",
  7195 => x"C0C0C0C0F8F99092",
  7196 => x"C0C0C0C0F8F99082",
  7197 => x"C0C0C0C0F8F990F8",
  7198 => x"C0C0C0C0F8F99080",
  7199 => x"C0C0C0C0F8F99090",
  7200 => x"C0C0C0C0F8A4C0C0",
  7201 => x"C0C0C0C0F8A4C0F9",
  7202 => x"C0C0C0C0F8A4C0A4",
  7203 => x"C0C0C0C0F8A4C0B0",
  7204 => x"C0C0C0C0F8A4C099",
  7205 => x"C0C0C0C0F8A4C092",
  7206 => x"C0C0C0C0F8A4C082",
  7207 => x"C0C0C0C0F8A4C0F8",
  7208 => x"C0C0C0C0F8A4C080",
  7209 => x"C0C0C0C0F8A4C090",
  7210 => x"C0C0C0C0F8A4F9C0",
  7211 => x"C0C0C0C0F8A4F9F9",
  7212 => x"C0C0C0C0F8A4F9A4",
  7213 => x"C0C0C0C0F8A4F9B0",
  7214 => x"C0C0C0C0F8A4F999",
  7215 => x"C0C0C0C0F8A4F992",
  7216 => x"C0C0C0C0F8A4F982",
  7217 => x"C0C0C0C0F8A4F9F8",
  7218 => x"C0C0C0C0F8A4F980",
  7219 => x"C0C0C0C0F8A4F990",
  7220 => x"C0C0C0C0F8A4A4C0",
  7221 => x"C0C0C0C0F8A4A4F9",
  7222 => x"C0C0C0C0F8A4A4A4",
  7223 => x"C0C0C0C0F8A4A4B0",
  7224 => x"C0C0C0C0F8A4A499",
  7225 => x"C0C0C0C0F8A4A492",
  7226 => x"C0C0C0C0F8A4A482",
  7227 => x"C0C0C0C0F8A4A4F8",
  7228 => x"C0C0C0C0F8A4A480",
  7229 => x"C0C0C0C0F8A4A490",
  7230 => x"C0C0C0C0F8A4B0C0",
  7231 => x"C0C0C0C0F8A4B0F9",
  7232 => x"C0C0C0C0F8A4B0A4",
  7233 => x"C0C0C0C0F8A4B0B0",
  7234 => x"C0C0C0C0F8A4B099",
  7235 => x"C0C0C0C0F8A4B092",
  7236 => x"C0C0C0C0F8A4B082",
  7237 => x"C0C0C0C0F8A4B0F8",
  7238 => x"C0C0C0C0F8A4B080",
  7239 => x"C0C0C0C0F8A4B090",
  7240 => x"C0C0C0C0F8A499C0",
  7241 => x"C0C0C0C0F8A499F9",
  7242 => x"C0C0C0C0F8A499A4",
  7243 => x"C0C0C0C0F8A499B0",
  7244 => x"C0C0C0C0F8A49999",
  7245 => x"C0C0C0C0F8A49992",
  7246 => x"C0C0C0C0F8A49982",
  7247 => x"C0C0C0C0F8A499F8",
  7248 => x"C0C0C0C0F8A49980",
  7249 => x"C0C0C0C0F8A49990",
  7250 => x"C0C0C0C0F8A492C0",
  7251 => x"C0C0C0C0F8A492F9",
  7252 => x"C0C0C0C0F8A492A4",
  7253 => x"C0C0C0C0F8A492B0",
  7254 => x"C0C0C0C0F8A49299",
  7255 => x"C0C0C0C0F8A49292",
  7256 => x"C0C0C0C0F8A49282",
  7257 => x"C0C0C0C0F8A492F8",
  7258 => x"C0C0C0C0F8A49280",
  7259 => x"C0C0C0C0F8A49290",
  7260 => x"C0C0C0C0F8A482C0",
  7261 => x"C0C0C0C0F8A482F9",
  7262 => x"C0C0C0C0F8A482A4",
  7263 => x"C0C0C0C0F8A482B0",
  7264 => x"C0C0C0C0F8A48299",
  7265 => x"C0C0C0C0F8A48292",
  7266 => x"C0C0C0C0F8A48282",
  7267 => x"C0C0C0C0F8A482F8",
  7268 => x"C0C0C0C0F8A48280",
  7269 => x"C0C0C0C0F8A48290",
  7270 => x"C0C0C0C0F8A4F8C0",
  7271 => x"C0C0C0C0F8A4F8F9",
  7272 => x"C0C0C0C0F8A4F8A4",
  7273 => x"C0C0C0C0F8A4F8B0",
  7274 => x"C0C0C0C0F8A4F899",
  7275 => x"C0C0C0C0F8A4F892",
  7276 => x"C0C0C0C0F8A4F882",
  7277 => x"C0C0C0C0F8A4F8F8",
  7278 => x"C0C0C0C0F8A4F880",
  7279 => x"C0C0C0C0F8A4F890",
  7280 => x"C0C0C0C0F8A480C0",
  7281 => x"C0C0C0C0F8A480F9",
  7282 => x"C0C0C0C0F8A480A4",
  7283 => x"C0C0C0C0F8A480B0",
  7284 => x"C0C0C0C0F8A48099",
  7285 => x"C0C0C0C0F8A48092",
  7286 => x"C0C0C0C0F8A48082",
  7287 => x"C0C0C0C0F8A480F8",
  7288 => x"C0C0C0C0F8A48080",
  7289 => x"C0C0C0C0F8A48090",
  7290 => x"C0C0C0C0F8A490C0",
  7291 => x"C0C0C0C0F8A490F9",
  7292 => x"C0C0C0C0F8A490A4",
  7293 => x"C0C0C0C0F8A490B0",
  7294 => x"C0C0C0C0F8A49099",
  7295 => x"C0C0C0C0F8A49092",
  7296 => x"C0C0C0C0F8A49082",
  7297 => x"C0C0C0C0F8A490F8",
  7298 => x"C0C0C0C0F8A49080",
  7299 => x"C0C0C0C0F8A49090",
  7300 => x"C0C0C0C0F8B0C0C0",
  7301 => x"C0C0C0C0F8B0C0F9",
  7302 => x"C0C0C0C0F8B0C0A4",
  7303 => x"C0C0C0C0F8B0C0B0",
  7304 => x"C0C0C0C0F8B0C099",
  7305 => x"C0C0C0C0F8B0C092",
  7306 => x"C0C0C0C0F8B0C082",
  7307 => x"C0C0C0C0F8B0C0F8",
  7308 => x"C0C0C0C0F8B0C080",
  7309 => x"C0C0C0C0F8B0C090",
  7310 => x"C0C0C0C0F8B0F9C0",
  7311 => x"C0C0C0C0F8B0F9F9",
  7312 => x"C0C0C0C0F8B0F9A4",
  7313 => x"C0C0C0C0F8B0F9B0",
  7314 => x"C0C0C0C0F8B0F999",
  7315 => x"C0C0C0C0F8B0F992",
  7316 => x"C0C0C0C0F8B0F982",
  7317 => x"C0C0C0C0F8B0F9F8",
  7318 => x"C0C0C0C0F8B0F980",
  7319 => x"C0C0C0C0F8B0F990",
  7320 => x"C0C0C0C0F8B0A4C0",
  7321 => x"C0C0C0C0F8B0A4F9",
  7322 => x"C0C0C0C0F8B0A4A4",
  7323 => x"C0C0C0C0F8B0A4B0",
  7324 => x"C0C0C0C0F8B0A499",
  7325 => x"C0C0C0C0F8B0A492",
  7326 => x"C0C0C0C0F8B0A482",
  7327 => x"C0C0C0C0F8B0A4F8",
  7328 => x"C0C0C0C0F8B0A480",
  7329 => x"C0C0C0C0F8B0A490",
  7330 => x"C0C0C0C0F8B0B0C0",
  7331 => x"C0C0C0C0F8B0B0F9",
  7332 => x"C0C0C0C0F8B0B0A4",
  7333 => x"C0C0C0C0F8B0B0B0",
  7334 => x"C0C0C0C0F8B0B099",
  7335 => x"C0C0C0C0F8B0B092",
  7336 => x"C0C0C0C0F8B0B082",
  7337 => x"C0C0C0C0F8B0B0F8",
  7338 => x"C0C0C0C0F8B0B080",
  7339 => x"C0C0C0C0F8B0B090",
  7340 => x"C0C0C0C0F8B099C0",
  7341 => x"C0C0C0C0F8B099F9",
  7342 => x"C0C0C0C0F8B099A4",
  7343 => x"C0C0C0C0F8B099B0",
  7344 => x"C0C0C0C0F8B09999",
  7345 => x"C0C0C0C0F8B09992",
  7346 => x"C0C0C0C0F8B09982",
  7347 => x"C0C0C0C0F8B099F8",
  7348 => x"C0C0C0C0F8B09980",
  7349 => x"C0C0C0C0F8B09990",
  7350 => x"C0C0C0C0F8B092C0",
  7351 => x"C0C0C0C0F8B092F9",
  7352 => x"C0C0C0C0F8B092A4",
  7353 => x"C0C0C0C0F8B092B0",
  7354 => x"C0C0C0C0F8B09299",
  7355 => x"C0C0C0C0F8B09292",
  7356 => x"C0C0C0C0F8B09282",
  7357 => x"C0C0C0C0F8B092F8",
  7358 => x"C0C0C0C0F8B09280",
  7359 => x"C0C0C0C0F8B09290",
  7360 => x"C0C0C0C0F8B082C0",
  7361 => x"C0C0C0C0F8B082F9",
  7362 => x"C0C0C0C0F8B082A4",
  7363 => x"C0C0C0C0F8B082B0",
  7364 => x"C0C0C0C0F8B08299",
  7365 => x"C0C0C0C0F8B08292",
  7366 => x"C0C0C0C0F8B08282",
  7367 => x"C0C0C0C0F8B082F8",
  7368 => x"C0C0C0C0F8B08280",
  7369 => x"C0C0C0C0F8B08290",
  7370 => x"C0C0C0C0F8B0F8C0",
  7371 => x"C0C0C0C0F8B0F8F9",
  7372 => x"C0C0C0C0F8B0F8A4",
  7373 => x"C0C0C0C0F8B0F8B0",
  7374 => x"C0C0C0C0F8B0F899",
  7375 => x"C0C0C0C0F8B0F892",
  7376 => x"C0C0C0C0F8B0F882",
  7377 => x"C0C0C0C0F8B0F8F8",
  7378 => x"C0C0C0C0F8B0F880",
  7379 => x"C0C0C0C0F8B0F890",
  7380 => x"C0C0C0C0F8B080C0",
  7381 => x"C0C0C0C0F8B080F9",
  7382 => x"C0C0C0C0F8B080A4",
  7383 => x"C0C0C0C0F8B080B0",
  7384 => x"C0C0C0C0F8B08099",
  7385 => x"C0C0C0C0F8B08092",
  7386 => x"C0C0C0C0F8B08082",
  7387 => x"C0C0C0C0F8B080F8",
  7388 => x"C0C0C0C0F8B08080",
  7389 => x"C0C0C0C0F8B08090",
  7390 => x"C0C0C0C0F8B090C0",
  7391 => x"C0C0C0C0F8B090F9",
  7392 => x"C0C0C0C0F8B090A4",
  7393 => x"C0C0C0C0F8B090B0",
  7394 => x"C0C0C0C0F8B09099",
  7395 => x"C0C0C0C0F8B09092",
  7396 => x"C0C0C0C0F8B09082",
  7397 => x"C0C0C0C0F8B090F8",
  7398 => x"C0C0C0C0F8B09080",
  7399 => x"C0C0C0C0F8B09090",
  7400 => x"C0C0C0C0F899C0C0",
  7401 => x"C0C0C0C0F899C0F9",
  7402 => x"C0C0C0C0F899C0A4",
  7403 => x"C0C0C0C0F899C0B0",
  7404 => x"C0C0C0C0F899C099",
  7405 => x"C0C0C0C0F899C092",
  7406 => x"C0C0C0C0F899C082",
  7407 => x"C0C0C0C0F899C0F8",
  7408 => x"C0C0C0C0F899C080",
  7409 => x"C0C0C0C0F899C090",
  7410 => x"C0C0C0C0F899F9C0",
  7411 => x"C0C0C0C0F899F9F9",
  7412 => x"C0C0C0C0F899F9A4",
  7413 => x"C0C0C0C0F899F9B0",
  7414 => x"C0C0C0C0F899F999",
  7415 => x"C0C0C0C0F899F992",
  7416 => x"C0C0C0C0F899F982",
  7417 => x"C0C0C0C0F899F9F8",
  7418 => x"C0C0C0C0F899F980",
  7419 => x"C0C0C0C0F899F990",
  7420 => x"C0C0C0C0F899A4C0",
  7421 => x"C0C0C0C0F899A4F9",
  7422 => x"C0C0C0C0F899A4A4",
  7423 => x"C0C0C0C0F899A4B0",
  7424 => x"C0C0C0C0F899A499",
  7425 => x"C0C0C0C0F899A492",
  7426 => x"C0C0C0C0F899A482",
  7427 => x"C0C0C0C0F899A4F8",
  7428 => x"C0C0C0C0F899A480",
  7429 => x"C0C0C0C0F899A490",
  7430 => x"C0C0C0C0F899B0C0",
  7431 => x"C0C0C0C0F899B0F9",
  7432 => x"C0C0C0C0F899B0A4",
  7433 => x"C0C0C0C0F899B0B0",
  7434 => x"C0C0C0C0F899B099",
  7435 => x"C0C0C0C0F899B092",
  7436 => x"C0C0C0C0F899B082",
  7437 => x"C0C0C0C0F899B0F8",
  7438 => x"C0C0C0C0F899B080",
  7439 => x"C0C0C0C0F899B090",
  7440 => x"C0C0C0C0F89999C0",
  7441 => x"C0C0C0C0F89999F9",
  7442 => x"C0C0C0C0F89999A4",
  7443 => x"C0C0C0C0F89999B0",
  7444 => x"C0C0C0C0F8999999",
  7445 => x"C0C0C0C0F8999992",
  7446 => x"C0C0C0C0F8999982",
  7447 => x"C0C0C0C0F89999F8",
  7448 => x"C0C0C0C0F8999980",
  7449 => x"C0C0C0C0F8999990",
  7450 => x"C0C0C0C0F89992C0",
  7451 => x"C0C0C0C0F89992F9",
  7452 => x"C0C0C0C0F89992A4",
  7453 => x"C0C0C0C0F89992B0",
  7454 => x"C0C0C0C0F8999299",
  7455 => x"C0C0C0C0F8999292",
  7456 => x"C0C0C0C0F8999282",
  7457 => x"C0C0C0C0F89992F8",
  7458 => x"C0C0C0C0F8999280",
  7459 => x"C0C0C0C0F8999290",
  7460 => x"C0C0C0C0F89982C0",
  7461 => x"C0C0C0C0F89982F9",
  7462 => x"C0C0C0C0F89982A4",
  7463 => x"C0C0C0C0F89982B0",
  7464 => x"C0C0C0C0F8998299",
  7465 => x"C0C0C0C0F8998292",
  7466 => x"C0C0C0C0F8998282",
  7467 => x"C0C0C0C0F89982F8",
  7468 => x"C0C0C0C0F8998280",
  7469 => x"C0C0C0C0F8998290",
  7470 => x"C0C0C0C0F899F8C0",
  7471 => x"C0C0C0C0F899F8F9",
  7472 => x"C0C0C0C0F899F8A4",
  7473 => x"C0C0C0C0F899F8B0",
  7474 => x"C0C0C0C0F899F899",
  7475 => x"C0C0C0C0F899F892",
  7476 => x"C0C0C0C0F899F882",
  7477 => x"C0C0C0C0F899F8F8",
  7478 => x"C0C0C0C0F899F880",
  7479 => x"C0C0C0C0F899F890",
  7480 => x"C0C0C0C0F89980C0",
  7481 => x"C0C0C0C0F89980F9",
  7482 => x"C0C0C0C0F89980A4",
  7483 => x"C0C0C0C0F89980B0",
  7484 => x"C0C0C0C0F8998099",
  7485 => x"C0C0C0C0F8998092",
  7486 => x"C0C0C0C0F8998082",
  7487 => x"C0C0C0C0F89980F8",
  7488 => x"C0C0C0C0F8998080",
  7489 => x"C0C0C0C0F8998090",
  7490 => x"C0C0C0C0F89990C0",
  7491 => x"C0C0C0C0F89990F9",
  7492 => x"C0C0C0C0F89990A4",
  7493 => x"C0C0C0C0F89990B0",
  7494 => x"C0C0C0C0F8999099",
  7495 => x"C0C0C0C0F8999092",
  7496 => x"C0C0C0C0F8999082",
  7497 => x"C0C0C0C0F89990F8",
  7498 => x"C0C0C0C0F8999080",
  7499 => x"C0C0C0C0F8999090",
  7500 => x"C0C0C0C0F892C0C0",
  7501 => x"C0C0C0C0F892C0F9",
  7502 => x"C0C0C0C0F892C0A4",
  7503 => x"C0C0C0C0F892C0B0",
  7504 => x"C0C0C0C0F892C099",
  7505 => x"C0C0C0C0F892C092",
  7506 => x"C0C0C0C0F892C082",
  7507 => x"C0C0C0C0F892C0F8",
  7508 => x"C0C0C0C0F892C080",
  7509 => x"C0C0C0C0F892C090",
  7510 => x"C0C0C0C0F892F9C0",
  7511 => x"C0C0C0C0F892F9F9",
  7512 => x"C0C0C0C0F892F9A4",
  7513 => x"C0C0C0C0F892F9B0",
  7514 => x"C0C0C0C0F892F999",
  7515 => x"C0C0C0C0F892F992",
  7516 => x"C0C0C0C0F892F982",
  7517 => x"C0C0C0C0F892F9F8",
  7518 => x"C0C0C0C0F892F980",
  7519 => x"C0C0C0C0F892F990",
  7520 => x"C0C0C0C0F892A4C0",
  7521 => x"C0C0C0C0F892A4F9",
  7522 => x"C0C0C0C0F892A4A4",
  7523 => x"C0C0C0C0F892A4B0",
  7524 => x"C0C0C0C0F892A499",
  7525 => x"C0C0C0C0F892A492",
  7526 => x"C0C0C0C0F892A482",
  7527 => x"C0C0C0C0F892A4F8",
  7528 => x"C0C0C0C0F892A480",
  7529 => x"C0C0C0C0F892A490",
  7530 => x"C0C0C0C0F892B0C0",
  7531 => x"C0C0C0C0F892B0F9",
  7532 => x"C0C0C0C0F892B0A4",
  7533 => x"C0C0C0C0F892B0B0",
  7534 => x"C0C0C0C0F892B099",
  7535 => x"C0C0C0C0F892B092",
  7536 => x"C0C0C0C0F892B082",
  7537 => x"C0C0C0C0F892B0F8",
  7538 => x"C0C0C0C0F892B080",
  7539 => x"C0C0C0C0F892B090",
  7540 => x"C0C0C0C0F89299C0",
  7541 => x"C0C0C0C0F89299F9",
  7542 => x"C0C0C0C0F89299A4",
  7543 => x"C0C0C0C0F89299B0",
  7544 => x"C0C0C0C0F8929999",
  7545 => x"C0C0C0C0F8929992",
  7546 => x"C0C0C0C0F8929982",
  7547 => x"C0C0C0C0F89299F8",
  7548 => x"C0C0C0C0F8929980",
  7549 => x"C0C0C0C0F8929990",
  7550 => x"C0C0C0C0F89292C0",
  7551 => x"C0C0C0C0F89292F9",
  7552 => x"C0C0C0C0F89292A4",
  7553 => x"C0C0C0C0F89292B0",
  7554 => x"C0C0C0C0F8929299",
  7555 => x"C0C0C0C0F8929292",
  7556 => x"C0C0C0C0F8929282",
  7557 => x"C0C0C0C0F89292F8",
  7558 => x"C0C0C0C0F8929280",
  7559 => x"C0C0C0C0F8929290",
  7560 => x"C0C0C0C0F89282C0",
  7561 => x"C0C0C0C0F89282F9",
  7562 => x"C0C0C0C0F89282A4",
  7563 => x"C0C0C0C0F89282B0",
  7564 => x"C0C0C0C0F8928299",
  7565 => x"C0C0C0C0F8928292",
  7566 => x"C0C0C0C0F8928282",
  7567 => x"C0C0C0C0F89282F8",
  7568 => x"C0C0C0C0F8928280",
  7569 => x"C0C0C0C0F8928290",
  7570 => x"C0C0C0C0F892F8C0",
  7571 => x"C0C0C0C0F892F8F9",
  7572 => x"C0C0C0C0F892F8A4",
  7573 => x"C0C0C0C0F892F8B0",
  7574 => x"C0C0C0C0F892F899",
  7575 => x"C0C0C0C0F892F892",
  7576 => x"C0C0C0C0F892F882",
  7577 => x"C0C0C0C0F892F8F8",
  7578 => x"C0C0C0C0F892F880",
  7579 => x"C0C0C0C0F892F890",
  7580 => x"C0C0C0C0F89280C0",
  7581 => x"C0C0C0C0F89280F9",
  7582 => x"C0C0C0C0F89280A4",
  7583 => x"C0C0C0C0F89280B0",
  7584 => x"C0C0C0C0F8928099",
  7585 => x"C0C0C0C0F8928092",
  7586 => x"C0C0C0C0F8928082",
  7587 => x"C0C0C0C0F89280F8",
  7588 => x"C0C0C0C0F8928080",
  7589 => x"C0C0C0C0F8928090",
  7590 => x"C0C0C0C0F89290C0",
  7591 => x"C0C0C0C0F89290F9",
  7592 => x"C0C0C0C0F89290A4",
  7593 => x"C0C0C0C0F89290B0",
  7594 => x"C0C0C0C0F8929099",
  7595 => x"C0C0C0C0F8929092",
  7596 => x"C0C0C0C0F8929082",
  7597 => x"C0C0C0C0F89290F8",
  7598 => x"C0C0C0C0F8929080",
  7599 => x"C0C0C0C0F8929090",
  7600 => x"C0C0C0C0F882C0C0",
  7601 => x"C0C0C0C0F882C0F9",
  7602 => x"C0C0C0C0F882C0A4",
  7603 => x"C0C0C0C0F882C0B0",
  7604 => x"C0C0C0C0F882C099",
  7605 => x"C0C0C0C0F882C092",
  7606 => x"C0C0C0C0F882C082",
  7607 => x"C0C0C0C0F882C0F8",
  7608 => x"C0C0C0C0F882C080",
  7609 => x"C0C0C0C0F882C090",
  7610 => x"C0C0C0C0F882F9C0",
  7611 => x"C0C0C0C0F882F9F9",
  7612 => x"C0C0C0C0F882F9A4",
  7613 => x"C0C0C0C0F882F9B0",
  7614 => x"C0C0C0C0F882F999",
  7615 => x"C0C0C0C0F882F992",
  7616 => x"C0C0C0C0F882F982",
  7617 => x"C0C0C0C0F882F9F8",
  7618 => x"C0C0C0C0F882F980",
  7619 => x"C0C0C0C0F882F990",
  7620 => x"C0C0C0C0F882A4C0",
  7621 => x"C0C0C0C0F882A4F9",
  7622 => x"C0C0C0C0F882A4A4",
  7623 => x"C0C0C0C0F882A4B0",
  7624 => x"C0C0C0C0F882A499",
  7625 => x"C0C0C0C0F882A492",
  7626 => x"C0C0C0C0F882A482",
  7627 => x"C0C0C0C0F882A4F8",
  7628 => x"C0C0C0C0F882A480",
  7629 => x"C0C0C0C0F882A490",
  7630 => x"C0C0C0C0F882B0C0",
  7631 => x"C0C0C0C0F882B0F9",
  7632 => x"C0C0C0C0F882B0A4",
  7633 => x"C0C0C0C0F882B0B0",
  7634 => x"C0C0C0C0F882B099",
  7635 => x"C0C0C0C0F882B092",
  7636 => x"C0C0C0C0F882B082",
  7637 => x"C0C0C0C0F882B0F8",
  7638 => x"C0C0C0C0F882B080",
  7639 => x"C0C0C0C0F882B090",
  7640 => x"C0C0C0C0F88299C0",
  7641 => x"C0C0C0C0F88299F9",
  7642 => x"C0C0C0C0F88299A4",
  7643 => x"C0C0C0C0F88299B0",
  7644 => x"C0C0C0C0F8829999",
  7645 => x"C0C0C0C0F8829992",
  7646 => x"C0C0C0C0F8829982",
  7647 => x"C0C0C0C0F88299F8",
  7648 => x"C0C0C0C0F8829980",
  7649 => x"C0C0C0C0F8829990",
  7650 => x"C0C0C0C0F88292C0",
  7651 => x"C0C0C0C0F88292F9",
  7652 => x"C0C0C0C0F88292A4",
  7653 => x"C0C0C0C0F88292B0",
  7654 => x"C0C0C0C0F8829299",
  7655 => x"C0C0C0C0F8829292",
  7656 => x"C0C0C0C0F8829282",
  7657 => x"C0C0C0C0F88292F8",
  7658 => x"C0C0C0C0F8829280",
  7659 => x"C0C0C0C0F8829290",
  7660 => x"C0C0C0C0F88282C0",
  7661 => x"C0C0C0C0F88282F9",
  7662 => x"C0C0C0C0F88282A4",
  7663 => x"C0C0C0C0F88282B0",
  7664 => x"C0C0C0C0F8828299",
  7665 => x"C0C0C0C0F8828292",
  7666 => x"C0C0C0C0F8828282",
  7667 => x"C0C0C0C0F88282F8",
  7668 => x"C0C0C0C0F8828280",
  7669 => x"C0C0C0C0F8828290",
  7670 => x"C0C0C0C0F882F8C0",
  7671 => x"C0C0C0C0F882F8F9",
  7672 => x"C0C0C0C0F882F8A4",
  7673 => x"C0C0C0C0F882F8B0",
  7674 => x"C0C0C0C0F882F899",
  7675 => x"C0C0C0C0F882F892",
  7676 => x"C0C0C0C0F882F882",
  7677 => x"C0C0C0C0F882F8F8",
  7678 => x"C0C0C0C0F882F880",
  7679 => x"C0C0C0C0F882F890",
  7680 => x"C0C0C0C0F88280C0",
  7681 => x"C0C0C0C0F88280F9",
  7682 => x"C0C0C0C0F88280A4",
  7683 => x"C0C0C0C0F88280B0",
  7684 => x"C0C0C0C0F8828099",
  7685 => x"C0C0C0C0F8828092",
  7686 => x"C0C0C0C0F8828082",
  7687 => x"C0C0C0C0F88280F8",
  7688 => x"C0C0C0C0F8828080",
  7689 => x"C0C0C0C0F8828090",
  7690 => x"C0C0C0C0F88290C0",
  7691 => x"C0C0C0C0F88290F9",
  7692 => x"C0C0C0C0F88290A4",
  7693 => x"C0C0C0C0F88290B0",
  7694 => x"C0C0C0C0F8829099",
  7695 => x"C0C0C0C0F8829092",
  7696 => x"C0C0C0C0F8829082",
  7697 => x"C0C0C0C0F88290F8",
  7698 => x"C0C0C0C0F8829080",
  7699 => x"C0C0C0C0F8829090",
  7700 => x"C0C0C0C0F8F8C0C0",
  7701 => x"C0C0C0C0F8F8C0F9",
  7702 => x"C0C0C0C0F8F8C0A4",
  7703 => x"C0C0C0C0F8F8C0B0",
  7704 => x"C0C0C0C0F8F8C099",
  7705 => x"C0C0C0C0F8F8C092",
  7706 => x"C0C0C0C0F8F8C082",
  7707 => x"C0C0C0C0F8F8C0F8",
  7708 => x"C0C0C0C0F8F8C080",
  7709 => x"C0C0C0C0F8F8C090",
  7710 => x"C0C0C0C0F8F8F9C0",
  7711 => x"C0C0C0C0F8F8F9F9",
  7712 => x"C0C0C0C0F8F8F9A4",
  7713 => x"C0C0C0C0F8F8F9B0",
  7714 => x"C0C0C0C0F8F8F999",
  7715 => x"C0C0C0C0F8F8F992",
  7716 => x"C0C0C0C0F8F8F982",
  7717 => x"C0C0C0C0F8F8F9F8",
  7718 => x"C0C0C0C0F8F8F980",
  7719 => x"C0C0C0C0F8F8F990",
  7720 => x"C0C0C0C0F8F8A4C0",
  7721 => x"C0C0C0C0F8F8A4F9",
  7722 => x"C0C0C0C0F8F8A4A4",
  7723 => x"C0C0C0C0F8F8A4B0",
  7724 => x"C0C0C0C0F8F8A499",
  7725 => x"C0C0C0C0F8F8A492",
  7726 => x"C0C0C0C0F8F8A482",
  7727 => x"C0C0C0C0F8F8A4F8",
  7728 => x"C0C0C0C0F8F8A480",
  7729 => x"C0C0C0C0F8F8A490",
  7730 => x"C0C0C0C0F8F8B0C0",
  7731 => x"C0C0C0C0F8F8B0F9",
  7732 => x"C0C0C0C0F8F8B0A4",
  7733 => x"C0C0C0C0F8F8B0B0",
  7734 => x"C0C0C0C0F8F8B099",
  7735 => x"C0C0C0C0F8F8B092",
  7736 => x"C0C0C0C0F8F8B082",
  7737 => x"C0C0C0C0F8F8B0F8",
  7738 => x"C0C0C0C0F8F8B080",
  7739 => x"C0C0C0C0F8F8B090",
  7740 => x"C0C0C0C0F8F899C0",
  7741 => x"C0C0C0C0F8F899F9",
  7742 => x"C0C0C0C0F8F899A4",
  7743 => x"C0C0C0C0F8F899B0",
  7744 => x"C0C0C0C0F8F89999",
  7745 => x"C0C0C0C0F8F89992",
  7746 => x"C0C0C0C0F8F89982",
  7747 => x"C0C0C0C0F8F899F8",
  7748 => x"C0C0C0C0F8F89980",
  7749 => x"C0C0C0C0F8F89990",
  7750 => x"C0C0C0C0F8F892C0",
  7751 => x"C0C0C0C0F8F892F9",
  7752 => x"C0C0C0C0F8F892A4",
  7753 => x"C0C0C0C0F8F892B0",
  7754 => x"C0C0C0C0F8F89299",
  7755 => x"C0C0C0C0F8F89292",
  7756 => x"C0C0C0C0F8F89282",
  7757 => x"C0C0C0C0F8F892F8",
  7758 => x"C0C0C0C0F8F89280",
  7759 => x"C0C0C0C0F8F89290",
  7760 => x"C0C0C0C0F8F882C0",
  7761 => x"C0C0C0C0F8F882F9",
  7762 => x"C0C0C0C0F8F882A4",
  7763 => x"C0C0C0C0F8F882B0",
  7764 => x"C0C0C0C0F8F88299",
  7765 => x"C0C0C0C0F8F88292",
  7766 => x"C0C0C0C0F8F88282",
  7767 => x"C0C0C0C0F8F882F8",
  7768 => x"C0C0C0C0F8F88280",
  7769 => x"C0C0C0C0F8F88290",
  7770 => x"C0C0C0C0F8F8F8C0",
  7771 => x"C0C0C0C0F8F8F8F9",
  7772 => x"C0C0C0C0F8F8F8A4",
  7773 => x"C0C0C0C0F8F8F8B0",
  7774 => x"C0C0C0C0F8F8F899",
  7775 => x"C0C0C0C0F8F8F892",
  7776 => x"C0C0C0C0F8F8F882",
  7777 => x"C0C0C0C0F8F8F8F8",
  7778 => x"C0C0C0C0F8F8F880",
  7779 => x"C0C0C0C0F8F8F890",
  7780 => x"C0C0C0C0F8F880C0",
  7781 => x"C0C0C0C0F8F880F9",
  7782 => x"C0C0C0C0F8F880A4",
  7783 => x"C0C0C0C0F8F880B0",
  7784 => x"C0C0C0C0F8F88099",
  7785 => x"C0C0C0C0F8F88092",
  7786 => x"C0C0C0C0F8F88082",
  7787 => x"C0C0C0C0F8F880F8",
  7788 => x"C0C0C0C0F8F88080",
  7789 => x"C0C0C0C0F8F88090",
  7790 => x"C0C0C0C0F8F890C0",
  7791 => x"C0C0C0C0F8F890F9",
  7792 => x"C0C0C0C0F8F890A4",
  7793 => x"C0C0C0C0F8F890B0",
  7794 => x"C0C0C0C0F8F89099",
  7795 => x"C0C0C0C0F8F89092",
  7796 => x"C0C0C0C0F8F89082",
  7797 => x"C0C0C0C0F8F890F8",
  7798 => x"C0C0C0C0F8F89080",
  7799 => x"C0C0C0C0F8F89090",
  7800 => x"C0C0C0C0F880C0C0",
  7801 => x"C0C0C0C0F880C0F9",
  7802 => x"C0C0C0C0F880C0A4",
  7803 => x"C0C0C0C0F880C0B0",
  7804 => x"C0C0C0C0F880C099",
  7805 => x"C0C0C0C0F880C092",
  7806 => x"C0C0C0C0F880C082",
  7807 => x"C0C0C0C0F880C0F8",
  7808 => x"C0C0C0C0F880C080",
  7809 => x"C0C0C0C0F880C090",
  7810 => x"C0C0C0C0F880F9C0",
  7811 => x"C0C0C0C0F880F9F9",
  7812 => x"C0C0C0C0F880F9A4",
  7813 => x"C0C0C0C0F880F9B0",
  7814 => x"C0C0C0C0F880F999",
  7815 => x"C0C0C0C0F880F992",
  7816 => x"C0C0C0C0F880F982",
  7817 => x"C0C0C0C0F880F9F8",
  7818 => x"C0C0C0C0F880F980",
  7819 => x"C0C0C0C0F880F990",
  7820 => x"C0C0C0C0F880A4C0",
  7821 => x"C0C0C0C0F880A4F9",
  7822 => x"C0C0C0C0F880A4A4",
  7823 => x"C0C0C0C0F880A4B0",
  7824 => x"C0C0C0C0F880A499",
  7825 => x"C0C0C0C0F880A492",
  7826 => x"C0C0C0C0F880A482",
  7827 => x"C0C0C0C0F880A4F8",
  7828 => x"C0C0C0C0F880A480",
  7829 => x"C0C0C0C0F880A490",
  7830 => x"C0C0C0C0F880B0C0",
  7831 => x"C0C0C0C0F880B0F9",
  7832 => x"C0C0C0C0F880B0A4",
  7833 => x"C0C0C0C0F880B0B0",
  7834 => x"C0C0C0C0F880B099",
  7835 => x"C0C0C0C0F880B092",
  7836 => x"C0C0C0C0F880B082",
  7837 => x"C0C0C0C0F880B0F8",
  7838 => x"C0C0C0C0F880B080",
  7839 => x"C0C0C0C0F880B090",
  7840 => x"C0C0C0C0F88099C0",
  7841 => x"C0C0C0C0F88099F9",
  7842 => x"C0C0C0C0F88099A4",
  7843 => x"C0C0C0C0F88099B0",
  7844 => x"C0C0C0C0F8809999",
  7845 => x"C0C0C0C0F8809992",
  7846 => x"C0C0C0C0F8809982",
  7847 => x"C0C0C0C0F88099F8",
  7848 => x"C0C0C0C0F8809980",
  7849 => x"C0C0C0C0F8809990",
  7850 => x"C0C0C0C0F88092C0",
  7851 => x"C0C0C0C0F88092F9",
  7852 => x"C0C0C0C0F88092A4",
  7853 => x"C0C0C0C0F88092B0",
  7854 => x"C0C0C0C0F8809299",
  7855 => x"C0C0C0C0F8809292",
  7856 => x"C0C0C0C0F8809282",
  7857 => x"C0C0C0C0F88092F8",
  7858 => x"C0C0C0C0F8809280",
  7859 => x"C0C0C0C0F8809290",
  7860 => x"C0C0C0C0F88082C0",
  7861 => x"C0C0C0C0F88082F9",
  7862 => x"C0C0C0C0F88082A4",
  7863 => x"C0C0C0C0F88082B0",
  7864 => x"C0C0C0C0F8808299",
  7865 => x"C0C0C0C0F8808292",
  7866 => x"C0C0C0C0F8808282",
  7867 => x"C0C0C0C0F88082F8",
  7868 => x"C0C0C0C0F8808280",
  7869 => x"C0C0C0C0F8808290",
  7870 => x"C0C0C0C0F880F8C0",
  7871 => x"C0C0C0C0F880F8F9",
  7872 => x"C0C0C0C0F880F8A4",
  7873 => x"C0C0C0C0F880F8B0",
  7874 => x"C0C0C0C0F880F899",
  7875 => x"C0C0C0C0F880F892",
  7876 => x"C0C0C0C0F880F882",
  7877 => x"C0C0C0C0F880F8F8",
  7878 => x"C0C0C0C0F880F880",
  7879 => x"C0C0C0C0F880F890",
  7880 => x"C0C0C0C0F88080C0",
  7881 => x"C0C0C0C0F88080F9",
  7882 => x"C0C0C0C0F88080A4",
  7883 => x"C0C0C0C0F88080B0",
  7884 => x"C0C0C0C0F8808099",
  7885 => x"C0C0C0C0F8808092",
  7886 => x"C0C0C0C0F8808082",
  7887 => x"C0C0C0C0F88080F8",
  7888 => x"C0C0C0C0F8808080",
  7889 => x"C0C0C0C0F8808090",
  7890 => x"C0C0C0C0F88090C0",
  7891 => x"C0C0C0C0F88090F9",
  7892 => x"C0C0C0C0F88090A4",
  7893 => x"C0C0C0C0F88090B0",
  7894 => x"C0C0C0C0F8809099",
  7895 => x"C0C0C0C0F8809092",
  7896 => x"C0C0C0C0F8809082",
  7897 => x"C0C0C0C0F88090F8",
  7898 => x"C0C0C0C0F8809080",
  7899 => x"C0C0C0C0F8809090",
  7900 => x"C0C0C0C0F890C0C0",
  7901 => x"C0C0C0C0F890C0F9",
  7902 => x"C0C0C0C0F890C0A4",
  7903 => x"C0C0C0C0F890C0B0",
  7904 => x"C0C0C0C0F890C099",
  7905 => x"C0C0C0C0F890C092",
  7906 => x"C0C0C0C0F890C082",
  7907 => x"C0C0C0C0F890C0F8",
  7908 => x"C0C0C0C0F890C080",
  7909 => x"C0C0C0C0F890C090",
  7910 => x"C0C0C0C0F890F9C0",
  7911 => x"C0C0C0C0F890F9F9",
  7912 => x"C0C0C0C0F890F9A4",
  7913 => x"C0C0C0C0F890F9B0",
  7914 => x"C0C0C0C0F890F999",
  7915 => x"C0C0C0C0F890F992",
  7916 => x"C0C0C0C0F890F982",
  7917 => x"C0C0C0C0F890F9F8",
  7918 => x"C0C0C0C0F890F980",
  7919 => x"C0C0C0C0F890F990",
  7920 => x"C0C0C0C0F890A4C0",
  7921 => x"C0C0C0C0F890A4F9",
  7922 => x"C0C0C0C0F890A4A4",
  7923 => x"C0C0C0C0F890A4B0",
  7924 => x"C0C0C0C0F890A499",
  7925 => x"C0C0C0C0F890A492",
  7926 => x"C0C0C0C0F890A482",
  7927 => x"C0C0C0C0F890A4F8",
  7928 => x"C0C0C0C0F890A480",
  7929 => x"C0C0C0C0F890A490",
  7930 => x"C0C0C0C0F890B0C0",
  7931 => x"C0C0C0C0F890B0F9",
  7932 => x"C0C0C0C0F890B0A4",
  7933 => x"C0C0C0C0F890B0B0",
  7934 => x"C0C0C0C0F890B099",
  7935 => x"C0C0C0C0F890B092",
  7936 => x"C0C0C0C0F890B082",
  7937 => x"C0C0C0C0F890B0F8",
  7938 => x"C0C0C0C0F890B080",
  7939 => x"C0C0C0C0F890B090",
  7940 => x"C0C0C0C0F89099C0",
  7941 => x"C0C0C0C0F89099F9",
  7942 => x"C0C0C0C0F89099A4",
  7943 => x"C0C0C0C0F89099B0",
  7944 => x"C0C0C0C0F8909999",
  7945 => x"C0C0C0C0F8909992",
  7946 => x"C0C0C0C0F8909982",
  7947 => x"C0C0C0C0F89099F8",
  7948 => x"C0C0C0C0F8909980",
  7949 => x"C0C0C0C0F8909990",
  7950 => x"C0C0C0C0F89092C0",
  7951 => x"C0C0C0C0F89092F9",
  7952 => x"C0C0C0C0F89092A4",
  7953 => x"C0C0C0C0F89092B0",
  7954 => x"C0C0C0C0F8909299",
  7955 => x"C0C0C0C0F8909292",
  7956 => x"C0C0C0C0F8909282",
  7957 => x"C0C0C0C0F89092F8",
  7958 => x"C0C0C0C0F8909280",
  7959 => x"C0C0C0C0F8909290",
  7960 => x"C0C0C0C0F89082C0",
  7961 => x"C0C0C0C0F89082F9",
  7962 => x"C0C0C0C0F89082A4",
  7963 => x"C0C0C0C0F89082B0",
  7964 => x"C0C0C0C0F8908299",
  7965 => x"C0C0C0C0F8908292",
  7966 => x"C0C0C0C0F8908282",
  7967 => x"C0C0C0C0F89082F8",
  7968 => x"C0C0C0C0F8908280",
  7969 => x"C0C0C0C0F8908290",
  7970 => x"C0C0C0C0F890F8C0",
  7971 => x"C0C0C0C0F890F8F9",
  7972 => x"C0C0C0C0F890F8A4",
  7973 => x"C0C0C0C0F890F8B0",
  7974 => x"C0C0C0C0F890F899",
  7975 => x"C0C0C0C0F890F892",
  7976 => x"C0C0C0C0F890F882",
  7977 => x"C0C0C0C0F890F8F8",
  7978 => x"C0C0C0C0F890F880",
  7979 => x"C0C0C0C0F890F890",
  7980 => x"C0C0C0C0F89080C0",
  7981 => x"C0C0C0C0F89080F9",
  7982 => x"C0C0C0C0F89080A4",
  7983 => x"C0C0C0C0F89080B0",
  7984 => x"C0C0C0C0F8908099",
  7985 => x"C0C0C0C0F8908092",
  7986 => x"C0C0C0C0F8908082",
  7987 => x"C0C0C0C0F89080F8",
  7988 => x"C0C0C0C0F8908080",
  7989 => x"C0C0C0C0F8908090",
  7990 => x"C0C0C0C0F89090C0",
  7991 => x"C0C0C0C0F89090F9",
  7992 => x"C0C0C0C0F89090A4",
  7993 => x"C0C0C0C0F89090B0",
  7994 => x"C0C0C0C0F8909099",
  7995 => x"C0C0C0C0F8909092",
  7996 => x"C0C0C0C0F8909082",
  7997 => x"C0C0C0C0F89090F8",
  7998 => x"C0C0C0C0F8909080",
  7999 => x"C0C0C0C0F8909090",
  8000 => x"C0C0C0C080C0C0C0",
  8001 => x"C0C0C0C080C0C0F9",
  8002 => x"C0C0C0C080C0C0A4",
  8003 => x"C0C0C0C080C0C0B0",
  8004 => x"C0C0C0C080C0C099",
  8005 => x"C0C0C0C080C0C092",
  8006 => x"C0C0C0C080C0C082",
  8007 => x"C0C0C0C080C0C0F8",
  8008 => x"C0C0C0C080C0C080",
  8009 => x"C0C0C0C080C0C090",
  8010 => x"C0C0C0C080C0F9C0",
  8011 => x"C0C0C0C080C0F9F9",
  8012 => x"C0C0C0C080C0F9A4",
  8013 => x"C0C0C0C080C0F9B0",
  8014 => x"C0C0C0C080C0F999",
  8015 => x"C0C0C0C080C0F992",
  8016 => x"C0C0C0C080C0F982",
  8017 => x"C0C0C0C080C0F9F8",
  8018 => x"C0C0C0C080C0F980",
  8019 => x"C0C0C0C080C0F990",
  8020 => x"C0C0C0C080C0A4C0",
  8021 => x"C0C0C0C080C0A4F9",
  8022 => x"C0C0C0C080C0A4A4",
  8023 => x"C0C0C0C080C0A4B0",
  8024 => x"C0C0C0C080C0A499",
  8025 => x"C0C0C0C080C0A492",
  8026 => x"C0C0C0C080C0A482",
  8027 => x"C0C0C0C080C0A4F8",
  8028 => x"C0C0C0C080C0A480",
  8029 => x"C0C0C0C080C0A490",
  8030 => x"C0C0C0C080C0B0C0",
  8031 => x"C0C0C0C080C0B0F9",
  8032 => x"C0C0C0C080C0B0A4",
  8033 => x"C0C0C0C080C0B0B0",
  8034 => x"C0C0C0C080C0B099",
  8035 => x"C0C0C0C080C0B092",
  8036 => x"C0C0C0C080C0B082",
  8037 => x"C0C0C0C080C0B0F8",
  8038 => x"C0C0C0C080C0B080",
  8039 => x"C0C0C0C080C0B090",
  8040 => x"C0C0C0C080C099C0",
  8041 => x"C0C0C0C080C099F9",
  8042 => x"C0C0C0C080C099A4",
  8043 => x"C0C0C0C080C099B0",
  8044 => x"C0C0C0C080C09999",
  8045 => x"C0C0C0C080C09992",
  8046 => x"C0C0C0C080C09982",
  8047 => x"C0C0C0C080C099F8",
  8048 => x"C0C0C0C080C09980",
  8049 => x"C0C0C0C080C09990",
  8050 => x"C0C0C0C080C092C0",
  8051 => x"C0C0C0C080C092F9",
  8052 => x"C0C0C0C080C092A4",
  8053 => x"C0C0C0C080C092B0",
  8054 => x"C0C0C0C080C09299",
  8055 => x"C0C0C0C080C09292",
  8056 => x"C0C0C0C080C09282",
  8057 => x"C0C0C0C080C092F8",
  8058 => x"C0C0C0C080C09280",
  8059 => x"C0C0C0C080C09290",
  8060 => x"C0C0C0C080C082C0",
  8061 => x"C0C0C0C080C082F9",
  8062 => x"C0C0C0C080C082A4",
  8063 => x"C0C0C0C080C082B0",
  8064 => x"C0C0C0C080C08299",
  8065 => x"C0C0C0C080C08292",
  8066 => x"C0C0C0C080C08282",
  8067 => x"C0C0C0C080C082F8",
  8068 => x"C0C0C0C080C08280",
  8069 => x"C0C0C0C080C08290",
  8070 => x"C0C0C0C080C0F8C0",
  8071 => x"C0C0C0C080C0F8F9",
  8072 => x"C0C0C0C080C0F8A4",
  8073 => x"C0C0C0C080C0F8B0",
  8074 => x"C0C0C0C080C0F899",
  8075 => x"C0C0C0C080C0F892",
  8076 => x"C0C0C0C080C0F882",
  8077 => x"C0C0C0C080C0F8F8",
  8078 => x"C0C0C0C080C0F880",
  8079 => x"C0C0C0C080C0F890",
  8080 => x"C0C0C0C080C080C0",
  8081 => x"C0C0C0C080C080F9",
  8082 => x"C0C0C0C080C080A4",
  8083 => x"C0C0C0C080C080B0",
  8084 => x"C0C0C0C080C08099",
  8085 => x"C0C0C0C080C08092",
  8086 => x"C0C0C0C080C08082",
  8087 => x"C0C0C0C080C080F8",
  8088 => x"C0C0C0C080C08080",
  8089 => x"C0C0C0C080C08090",
  8090 => x"C0C0C0C080C090C0",
  8091 => x"C0C0C0C080C090F9",
  8092 => x"C0C0C0C080C090A4",
  8093 => x"C0C0C0C080C090B0",
  8094 => x"C0C0C0C080C09099",
  8095 => x"C0C0C0C080C09092",
  8096 => x"C0C0C0C080C09082",
  8097 => x"C0C0C0C080C090F8",
  8098 => x"C0C0C0C080C09080",
  8099 => x"C0C0C0C080C09090",
  8100 => x"C0C0C0C080F9C0C0",
  8101 => x"C0C0C0C080F9C0F9",
  8102 => x"C0C0C0C080F9C0A4",
  8103 => x"C0C0C0C080F9C0B0",
  8104 => x"C0C0C0C080F9C099",
  8105 => x"C0C0C0C080F9C092",
  8106 => x"C0C0C0C080F9C082",
  8107 => x"C0C0C0C080F9C0F8",
  8108 => x"C0C0C0C080F9C080",
  8109 => x"C0C0C0C080F9C090",
  8110 => x"C0C0C0C080F9F9C0",
  8111 => x"C0C0C0C080F9F9F9",
  8112 => x"C0C0C0C080F9F9A4",
  8113 => x"C0C0C0C080F9F9B0",
  8114 => x"C0C0C0C080F9F999",
  8115 => x"C0C0C0C080F9F992",
  8116 => x"C0C0C0C080F9F982",
  8117 => x"C0C0C0C080F9F9F8",
  8118 => x"C0C0C0C080F9F980",
  8119 => x"C0C0C0C080F9F990",
  8120 => x"C0C0C0C080F9A4C0",
  8121 => x"C0C0C0C080F9A4F9",
  8122 => x"C0C0C0C080F9A4A4",
  8123 => x"C0C0C0C080F9A4B0",
  8124 => x"C0C0C0C080F9A499",
  8125 => x"C0C0C0C080F9A492",
  8126 => x"C0C0C0C080F9A482",
  8127 => x"C0C0C0C080F9A4F8",
  8128 => x"C0C0C0C080F9A480",
  8129 => x"C0C0C0C080F9A490",
  8130 => x"C0C0C0C080F9B0C0",
  8131 => x"C0C0C0C080F9B0F9",
  8132 => x"C0C0C0C080F9B0A4",
  8133 => x"C0C0C0C080F9B0B0",
  8134 => x"C0C0C0C080F9B099",
  8135 => x"C0C0C0C080F9B092",
  8136 => x"C0C0C0C080F9B082",
  8137 => x"C0C0C0C080F9B0F8",
  8138 => x"C0C0C0C080F9B080",
  8139 => x"C0C0C0C080F9B090",
  8140 => x"C0C0C0C080F999C0",
  8141 => x"C0C0C0C080F999F9",
  8142 => x"C0C0C0C080F999A4",
  8143 => x"C0C0C0C080F999B0",
  8144 => x"C0C0C0C080F99999",
  8145 => x"C0C0C0C080F99992",
  8146 => x"C0C0C0C080F99982",
  8147 => x"C0C0C0C080F999F8",
  8148 => x"C0C0C0C080F99980",
  8149 => x"C0C0C0C080F99990",
  8150 => x"C0C0C0C080F992C0",
  8151 => x"C0C0C0C080F992F9",
  8152 => x"C0C0C0C080F992A4",
  8153 => x"C0C0C0C080F992B0",
  8154 => x"C0C0C0C080F99299",
  8155 => x"C0C0C0C080F99292",
  8156 => x"C0C0C0C080F99282",
  8157 => x"C0C0C0C080F992F8",
  8158 => x"C0C0C0C080F99280",
  8159 => x"C0C0C0C080F99290",
  8160 => x"C0C0C0C080F982C0",
  8161 => x"C0C0C0C080F982F9",
  8162 => x"C0C0C0C080F982A4",
  8163 => x"C0C0C0C080F982B0",
  8164 => x"C0C0C0C080F98299",
  8165 => x"C0C0C0C080F98292",
  8166 => x"C0C0C0C080F98282",
  8167 => x"C0C0C0C080F982F8",
  8168 => x"C0C0C0C080F98280",
  8169 => x"C0C0C0C080F98290",
  8170 => x"C0C0C0C080F9F8C0",
  8171 => x"C0C0C0C080F9F8F9",
  8172 => x"C0C0C0C080F9F8A4",
  8173 => x"C0C0C0C080F9F8B0",
  8174 => x"C0C0C0C080F9F899",
  8175 => x"C0C0C0C080F9F892",
  8176 => x"C0C0C0C080F9F882",
  8177 => x"C0C0C0C080F9F8F8",
  8178 => x"C0C0C0C080F9F880",
  8179 => x"C0C0C0C080F9F890",
  8180 => x"C0C0C0C080F980C0",
  8181 => x"C0C0C0C080F980F9",
  8182 => x"C0C0C0C080F980A4",
  8183 => x"C0C0C0C080F980B0",
  8184 => x"C0C0C0C080F98099",
  8185 => x"C0C0C0C080F98092",
  8186 => x"C0C0C0C080F98082",
  8187 => x"C0C0C0C080F980F8",
  8188 => x"C0C0C0C080F98080",
  8189 => x"C0C0C0C080F98090",
  8190 => x"C0C0C0C080F990C0",
  8191 => x"C0C0C0C080F990F9",
  8192 => x"C0C0C0C080F990A4",
  8193 => x"C0C0C0C080F990B0",
  8194 => x"C0C0C0C080F99099",
  8195 => x"C0C0C0C080F99092",
  8196 => x"C0C0C0C080F99082",
  8197 => x"C0C0C0C080F990F8",
  8198 => x"C0C0C0C080F99080",
  8199 => x"C0C0C0C080F99090",
  8200 => x"C0C0C0C080A4C0C0",
  8201 => x"C0C0C0C080A4C0F9",
  8202 => x"C0C0C0C080A4C0A4",
  8203 => x"C0C0C0C080A4C0B0",
  8204 => x"C0C0C0C080A4C099",
  8205 => x"C0C0C0C080A4C092",
  8206 => x"C0C0C0C080A4C082",
  8207 => x"C0C0C0C080A4C0F8",
  8208 => x"C0C0C0C080A4C080",
  8209 => x"C0C0C0C080A4C090",
  8210 => x"C0C0C0C080A4F9C0",
  8211 => x"C0C0C0C080A4F9F9",
  8212 => x"C0C0C0C080A4F9A4",
  8213 => x"C0C0C0C080A4F9B0",
  8214 => x"C0C0C0C080A4F999",
  8215 => x"C0C0C0C080A4F992",
  8216 => x"C0C0C0C080A4F982",
  8217 => x"C0C0C0C080A4F9F8",
  8218 => x"C0C0C0C080A4F980",
  8219 => x"C0C0C0C080A4F990",
  8220 => x"C0C0C0C080A4A4C0",
  8221 => x"C0C0C0C080A4A4F9",
  8222 => x"C0C0C0C080A4A4A4",
  8223 => x"C0C0C0C080A4A4B0",
  8224 => x"C0C0C0C080A4A499",
  8225 => x"C0C0C0C080A4A492",
  8226 => x"C0C0C0C080A4A482",
  8227 => x"C0C0C0C080A4A4F8",
  8228 => x"C0C0C0C080A4A480",
  8229 => x"C0C0C0C080A4A490",
  8230 => x"C0C0C0C080A4B0C0",
  8231 => x"C0C0C0C080A4B0F9",
  8232 => x"C0C0C0C080A4B0A4",
  8233 => x"C0C0C0C080A4B0B0",
  8234 => x"C0C0C0C080A4B099",
  8235 => x"C0C0C0C080A4B092",
  8236 => x"C0C0C0C080A4B082",
  8237 => x"C0C0C0C080A4B0F8",
  8238 => x"C0C0C0C080A4B080",
  8239 => x"C0C0C0C080A4B090",
  8240 => x"C0C0C0C080A499C0",
  8241 => x"C0C0C0C080A499F9",
  8242 => x"C0C0C0C080A499A4",
  8243 => x"C0C0C0C080A499B0",
  8244 => x"C0C0C0C080A49999",
  8245 => x"C0C0C0C080A49992",
  8246 => x"C0C0C0C080A49982",
  8247 => x"C0C0C0C080A499F8",
  8248 => x"C0C0C0C080A49980",
  8249 => x"C0C0C0C080A49990",
  8250 => x"C0C0C0C080A492C0",
  8251 => x"C0C0C0C080A492F9",
  8252 => x"C0C0C0C080A492A4",
  8253 => x"C0C0C0C080A492B0",
  8254 => x"C0C0C0C080A49299",
  8255 => x"C0C0C0C080A49292",
  8256 => x"C0C0C0C080A49282",
  8257 => x"C0C0C0C080A492F8",
  8258 => x"C0C0C0C080A49280",
  8259 => x"C0C0C0C080A49290",
  8260 => x"C0C0C0C080A482C0",
  8261 => x"C0C0C0C080A482F9",
  8262 => x"C0C0C0C080A482A4",
  8263 => x"C0C0C0C080A482B0",
  8264 => x"C0C0C0C080A48299",
  8265 => x"C0C0C0C080A48292",
  8266 => x"C0C0C0C080A48282",
  8267 => x"C0C0C0C080A482F8",
  8268 => x"C0C0C0C080A48280",
  8269 => x"C0C0C0C080A48290",
  8270 => x"C0C0C0C080A4F8C0",
  8271 => x"C0C0C0C080A4F8F9",
  8272 => x"C0C0C0C080A4F8A4",
  8273 => x"C0C0C0C080A4F8B0",
  8274 => x"C0C0C0C080A4F899",
  8275 => x"C0C0C0C080A4F892",
  8276 => x"C0C0C0C080A4F882",
  8277 => x"C0C0C0C080A4F8F8",
  8278 => x"C0C0C0C080A4F880",
  8279 => x"C0C0C0C080A4F890",
  8280 => x"C0C0C0C080A480C0",
  8281 => x"C0C0C0C080A480F9",
  8282 => x"C0C0C0C080A480A4",
  8283 => x"C0C0C0C080A480B0",
  8284 => x"C0C0C0C080A48099",
  8285 => x"C0C0C0C080A48092",
  8286 => x"C0C0C0C080A48082",
  8287 => x"C0C0C0C080A480F8",
  8288 => x"C0C0C0C080A48080",
  8289 => x"C0C0C0C080A48090",
  8290 => x"C0C0C0C080A490C0",
  8291 => x"C0C0C0C080A490F9",
  8292 => x"C0C0C0C080A490A4",
  8293 => x"C0C0C0C080A490B0",
  8294 => x"C0C0C0C080A49099",
  8295 => x"C0C0C0C080A49092",
  8296 => x"C0C0C0C080A49082",
  8297 => x"C0C0C0C080A490F8",
  8298 => x"C0C0C0C080A49080",
  8299 => x"C0C0C0C080A49090",
  8300 => x"C0C0C0C080B0C0C0",
  8301 => x"C0C0C0C080B0C0F9",
  8302 => x"C0C0C0C080B0C0A4",
  8303 => x"C0C0C0C080B0C0B0",
  8304 => x"C0C0C0C080B0C099",
  8305 => x"C0C0C0C080B0C092",
  8306 => x"C0C0C0C080B0C082",
  8307 => x"C0C0C0C080B0C0F8",
  8308 => x"C0C0C0C080B0C080",
  8309 => x"C0C0C0C080B0C090",
  8310 => x"C0C0C0C080B0F9C0",
  8311 => x"C0C0C0C080B0F9F9",
  8312 => x"C0C0C0C080B0F9A4",
  8313 => x"C0C0C0C080B0F9B0",
  8314 => x"C0C0C0C080B0F999",
  8315 => x"C0C0C0C080B0F992",
  8316 => x"C0C0C0C080B0F982",
  8317 => x"C0C0C0C080B0F9F8",
  8318 => x"C0C0C0C080B0F980",
  8319 => x"C0C0C0C080B0F990",
  8320 => x"C0C0C0C080B0A4C0",
  8321 => x"C0C0C0C080B0A4F9",
  8322 => x"C0C0C0C080B0A4A4",
  8323 => x"C0C0C0C080B0A4B0",
  8324 => x"C0C0C0C080B0A499",
  8325 => x"C0C0C0C080B0A492",
  8326 => x"C0C0C0C080B0A482",
  8327 => x"C0C0C0C080B0A4F8",
  8328 => x"C0C0C0C080B0A480",
  8329 => x"C0C0C0C080B0A490",
  8330 => x"C0C0C0C080B0B0C0",
  8331 => x"C0C0C0C080B0B0F9",
  8332 => x"C0C0C0C080B0B0A4",
  8333 => x"C0C0C0C080B0B0B0",
  8334 => x"C0C0C0C080B0B099",
  8335 => x"C0C0C0C080B0B092",
  8336 => x"C0C0C0C080B0B082",
  8337 => x"C0C0C0C080B0B0F8",
  8338 => x"C0C0C0C080B0B080",
  8339 => x"C0C0C0C080B0B090",
  8340 => x"C0C0C0C080B099C0",
  8341 => x"C0C0C0C080B099F9",
  8342 => x"C0C0C0C080B099A4",
  8343 => x"C0C0C0C080B099B0",
  8344 => x"C0C0C0C080B09999",
  8345 => x"C0C0C0C080B09992",
  8346 => x"C0C0C0C080B09982",
  8347 => x"C0C0C0C080B099F8",
  8348 => x"C0C0C0C080B09980",
  8349 => x"C0C0C0C080B09990",
  8350 => x"C0C0C0C080B092C0",
  8351 => x"C0C0C0C080B092F9",
  8352 => x"C0C0C0C080B092A4",
  8353 => x"C0C0C0C080B092B0",
  8354 => x"C0C0C0C080B09299",
  8355 => x"C0C0C0C080B09292",
  8356 => x"C0C0C0C080B09282",
  8357 => x"C0C0C0C080B092F8",
  8358 => x"C0C0C0C080B09280",
  8359 => x"C0C0C0C080B09290",
  8360 => x"C0C0C0C080B082C0",
  8361 => x"C0C0C0C080B082F9",
  8362 => x"C0C0C0C080B082A4",
  8363 => x"C0C0C0C080B082B0",
  8364 => x"C0C0C0C080B08299",
  8365 => x"C0C0C0C080B08292",
  8366 => x"C0C0C0C080B08282",
  8367 => x"C0C0C0C080B082F8",
  8368 => x"C0C0C0C080B08280",
  8369 => x"C0C0C0C080B08290",
  8370 => x"C0C0C0C080B0F8C0",
  8371 => x"C0C0C0C080B0F8F9",
  8372 => x"C0C0C0C080B0F8A4",
  8373 => x"C0C0C0C080B0F8B0",
  8374 => x"C0C0C0C080B0F899",
  8375 => x"C0C0C0C080B0F892",
  8376 => x"C0C0C0C080B0F882",
  8377 => x"C0C0C0C080B0F8F8",
  8378 => x"C0C0C0C080B0F880",
  8379 => x"C0C0C0C080B0F890",
  8380 => x"C0C0C0C080B080C0",
  8381 => x"C0C0C0C080B080F9",
  8382 => x"C0C0C0C080B080A4",
  8383 => x"C0C0C0C080B080B0",
  8384 => x"C0C0C0C080B08099",
  8385 => x"C0C0C0C080B08092",
  8386 => x"C0C0C0C080B08082",
  8387 => x"C0C0C0C080B080F8",
  8388 => x"C0C0C0C080B08080",
  8389 => x"C0C0C0C080B08090",
  8390 => x"C0C0C0C080B090C0",
  8391 => x"C0C0C0C080B090F9",
  8392 => x"C0C0C0C080B090A4",
  8393 => x"C0C0C0C080B090B0",
  8394 => x"C0C0C0C080B09099",
  8395 => x"C0C0C0C080B09092",
  8396 => x"C0C0C0C080B09082",
  8397 => x"C0C0C0C080B090F8",
  8398 => x"C0C0C0C080B09080",
  8399 => x"C0C0C0C080B09090",
  8400 => x"C0C0C0C08099C0C0",
  8401 => x"C0C0C0C08099C0F9",
  8402 => x"C0C0C0C08099C0A4",
  8403 => x"C0C0C0C08099C0B0",
  8404 => x"C0C0C0C08099C099",
  8405 => x"C0C0C0C08099C092",
  8406 => x"C0C0C0C08099C082",
  8407 => x"C0C0C0C08099C0F8",
  8408 => x"C0C0C0C08099C080",
  8409 => x"C0C0C0C08099C090",
  8410 => x"C0C0C0C08099F9C0",
  8411 => x"C0C0C0C08099F9F9",
  8412 => x"C0C0C0C08099F9A4",
  8413 => x"C0C0C0C08099F9B0",
  8414 => x"C0C0C0C08099F999",
  8415 => x"C0C0C0C08099F992",
  8416 => x"C0C0C0C08099F982",
  8417 => x"C0C0C0C08099F9F8",
  8418 => x"C0C0C0C08099F980",
  8419 => x"C0C0C0C08099F990",
  8420 => x"C0C0C0C08099A4C0",
  8421 => x"C0C0C0C08099A4F9",
  8422 => x"C0C0C0C08099A4A4",
  8423 => x"C0C0C0C08099A4B0",
  8424 => x"C0C0C0C08099A499",
  8425 => x"C0C0C0C08099A492",
  8426 => x"C0C0C0C08099A482",
  8427 => x"C0C0C0C08099A4F8",
  8428 => x"C0C0C0C08099A480",
  8429 => x"C0C0C0C08099A490",
  8430 => x"C0C0C0C08099B0C0",
  8431 => x"C0C0C0C08099B0F9",
  8432 => x"C0C0C0C08099B0A4",
  8433 => x"C0C0C0C08099B0B0",
  8434 => x"C0C0C0C08099B099",
  8435 => x"C0C0C0C08099B092",
  8436 => x"C0C0C0C08099B082",
  8437 => x"C0C0C0C08099B0F8",
  8438 => x"C0C0C0C08099B080",
  8439 => x"C0C0C0C08099B090",
  8440 => x"C0C0C0C0809999C0",
  8441 => x"C0C0C0C0809999F9",
  8442 => x"C0C0C0C0809999A4",
  8443 => x"C0C0C0C0809999B0",
  8444 => x"C0C0C0C080999999",
  8445 => x"C0C0C0C080999992",
  8446 => x"C0C0C0C080999982",
  8447 => x"C0C0C0C0809999F8",
  8448 => x"C0C0C0C080999980",
  8449 => x"C0C0C0C080999990",
  8450 => x"C0C0C0C0809992C0",
  8451 => x"C0C0C0C0809992F9",
  8452 => x"C0C0C0C0809992A4",
  8453 => x"C0C0C0C0809992B0",
  8454 => x"C0C0C0C080999299",
  8455 => x"C0C0C0C080999292",
  8456 => x"C0C0C0C080999282",
  8457 => x"C0C0C0C0809992F8",
  8458 => x"C0C0C0C080999280",
  8459 => x"C0C0C0C080999290",
  8460 => x"C0C0C0C0809982C0",
  8461 => x"C0C0C0C0809982F9",
  8462 => x"C0C0C0C0809982A4",
  8463 => x"C0C0C0C0809982B0",
  8464 => x"C0C0C0C080998299",
  8465 => x"C0C0C0C080998292",
  8466 => x"C0C0C0C080998282",
  8467 => x"C0C0C0C0809982F8",
  8468 => x"C0C0C0C080998280",
  8469 => x"C0C0C0C080998290",
  8470 => x"C0C0C0C08099F8C0",
  8471 => x"C0C0C0C08099F8F9",
  8472 => x"C0C0C0C08099F8A4",
  8473 => x"C0C0C0C08099F8B0",
  8474 => x"C0C0C0C08099F899",
  8475 => x"C0C0C0C08099F892",
  8476 => x"C0C0C0C08099F882",
  8477 => x"C0C0C0C08099F8F8",
  8478 => x"C0C0C0C08099F880",
  8479 => x"C0C0C0C08099F890",
  8480 => x"C0C0C0C0809980C0",
  8481 => x"C0C0C0C0809980F9",
  8482 => x"C0C0C0C0809980A4",
  8483 => x"C0C0C0C0809980B0",
  8484 => x"C0C0C0C080998099",
  8485 => x"C0C0C0C080998092",
  8486 => x"C0C0C0C080998082",
  8487 => x"C0C0C0C0809980F8",
  8488 => x"C0C0C0C080998080",
  8489 => x"C0C0C0C080998090",
  8490 => x"C0C0C0C0809990C0",
  8491 => x"C0C0C0C0809990F9",
  8492 => x"C0C0C0C0809990A4",
  8493 => x"C0C0C0C0809990B0",
  8494 => x"C0C0C0C080999099",
  8495 => x"C0C0C0C080999092",
  8496 => x"C0C0C0C080999082",
  8497 => x"C0C0C0C0809990F8",
  8498 => x"C0C0C0C080999080",
  8499 => x"C0C0C0C080999090",
  8500 => x"C0C0C0C08092C0C0",
  8501 => x"C0C0C0C08092C0F9",
  8502 => x"C0C0C0C08092C0A4",
  8503 => x"C0C0C0C08092C0B0",
  8504 => x"C0C0C0C08092C099",
  8505 => x"C0C0C0C08092C092",
  8506 => x"C0C0C0C08092C082",
  8507 => x"C0C0C0C08092C0F8",
  8508 => x"C0C0C0C08092C080",
  8509 => x"C0C0C0C08092C090",
  8510 => x"C0C0C0C08092F9C0",
  8511 => x"C0C0C0C08092F9F9",
  8512 => x"C0C0C0C08092F9A4",
  8513 => x"C0C0C0C08092F9B0",
  8514 => x"C0C0C0C08092F999",
  8515 => x"C0C0C0C08092F992",
  8516 => x"C0C0C0C08092F982",
  8517 => x"C0C0C0C08092F9F8",
  8518 => x"C0C0C0C08092F980",
  8519 => x"C0C0C0C08092F990",
  8520 => x"C0C0C0C08092A4C0",
  8521 => x"C0C0C0C08092A4F9",
  8522 => x"C0C0C0C08092A4A4",
  8523 => x"C0C0C0C08092A4B0",
  8524 => x"C0C0C0C08092A499",
  8525 => x"C0C0C0C08092A492",
  8526 => x"C0C0C0C08092A482",
  8527 => x"C0C0C0C08092A4F8",
  8528 => x"C0C0C0C08092A480",
  8529 => x"C0C0C0C08092A490",
  8530 => x"C0C0C0C08092B0C0",
  8531 => x"C0C0C0C08092B0F9",
  8532 => x"C0C0C0C08092B0A4",
  8533 => x"C0C0C0C08092B0B0",
  8534 => x"C0C0C0C08092B099",
  8535 => x"C0C0C0C08092B092",
  8536 => x"C0C0C0C08092B082",
  8537 => x"C0C0C0C08092B0F8",
  8538 => x"C0C0C0C08092B080",
  8539 => x"C0C0C0C08092B090",
  8540 => x"C0C0C0C0809299C0",
  8541 => x"C0C0C0C0809299F9",
  8542 => x"C0C0C0C0809299A4",
  8543 => x"C0C0C0C0809299B0",
  8544 => x"C0C0C0C080929999",
  8545 => x"C0C0C0C080929992",
  8546 => x"C0C0C0C080929982",
  8547 => x"C0C0C0C0809299F8",
  8548 => x"C0C0C0C080929980",
  8549 => x"C0C0C0C080929990",
  8550 => x"C0C0C0C0809292C0",
  8551 => x"C0C0C0C0809292F9",
  8552 => x"C0C0C0C0809292A4",
  8553 => x"C0C0C0C0809292B0",
  8554 => x"C0C0C0C080929299",
  8555 => x"C0C0C0C080929292",
  8556 => x"C0C0C0C080929282",
  8557 => x"C0C0C0C0809292F8",
  8558 => x"C0C0C0C080929280",
  8559 => x"C0C0C0C080929290",
  8560 => x"C0C0C0C0809282C0",
  8561 => x"C0C0C0C0809282F9",
  8562 => x"C0C0C0C0809282A4",
  8563 => x"C0C0C0C0809282B0",
  8564 => x"C0C0C0C080928299",
  8565 => x"C0C0C0C080928292",
  8566 => x"C0C0C0C080928282",
  8567 => x"C0C0C0C0809282F8",
  8568 => x"C0C0C0C080928280",
  8569 => x"C0C0C0C080928290",
  8570 => x"C0C0C0C08092F8C0",
  8571 => x"C0C0C0C08092F8F9",
  8572 => x"C0C0C0C08092F8A4",
  8573 => x"C0C0C0C08092F8B0",
  8574 => x"C0C0C0C08092F899",
  8575 => x"C0C0C0C08092F892",
  8576 => x"C0C0C0C08092F882",
  8577 => x"C0C0C0C08092F8F8",
  8578 => x"C0C0C0C08092F880",
  8579 => x"C0C0C0C08092F890",
  8580 => x"C0C0C0C0809280C0",
  8581 => x"C0C0C0C0809280F9",
  8582 => x"C0C0C0C0809280A4",
  8583 => x"C0C0C0C0809280B0",
  8584 => x"C0C0C0C080928099",
  8585 => x"C0C0C0C080928092",
  8586 => x"C0C0C0C080928082",
  8587 => x"C0C0C0C0809280F8",
  8588 => x"C0C0C0C080928080",
  8589 => x"C0C0C0C080928090",
  8590 => x"C0C0C0C0809290C0",
  8591 => x"C0C0C0C0809290F9",
  8592 => x"C0C0C0C0809290A4",
  8593 => x"C0C0C0C0809290B0",
  8594 => x"C0C0C0C080929099",
  8595 => x"C0C0C0C080929092",
  8596 => x"C0C0C0C080929082",
  8597 => x"C0C0C0C0809290F8",
  8598 => x"C0C0C0C080929080",
  8599 => x"C0C0C0C080929090",
  8600 => x"C0C0C0C08082C0C0",
  8601 => x"C0C0C0C08082C0F9",
  8602 => x"C0C0C0C08082C0A4",
  8603 => x"C0C0C0C08082C0B0",
  8604 => x"C0C0C0C08082C099",
  8605 => x"C0C0C0C08082C092",
  8606 => x"C0C0C0C08082C082",
  8607 => x"C0C0C0C08082C0F8",
  8608 => x"C0C0C0C08082C080",
  8609 => x"C0C0C0C08082C090",
  8610 => x"C0C0C0C08082F9C0",
  8611 => x"C0C0C0C08082F9F9",
  8612 => x"C0C0C0C08082F9A4",
  8613 => x"C0C0C0C08082F9B0",
  8614 => x"C0C0C0C08082F999",
  8615 => x"C0C0C0C08082F992",
  8616 => x"C0C0C0C08082F982",
  8617 => x"C0C0C0C08082F9F8",
  8618 => x"C0C0C0C08082F980",
  8619 => x"C0C0C0C08082F990",
  8620 => x"C0C0C0C08082A4C0",
  8621 => x"C0C0C0C08082A4F9",
  8622 => x"C0C0C0C08082A4A4",
  8623 => x"C0C0C0C08082A4B0",
  8624 => x"C0C0C0C08082A499",
  8625 => x"C0C0C0C08082A492",
  8626 => x"C0C0C0C08082A482",
  8627 => x"C0C0C0C08082A4F8",
  8628 => x"C0C0C0C08082A480",
  8629 => x"C0C0C0C08082A490",
  8630 => x"C0C0C0C08082B0C0",
  8631 => x"C0C0C0C08082B0F9",
  8632 => x"C0C0C0C08082B0A4",
  8633 => x"C0C0C0C08082B0B0",
  8634 => x"C0C0C0C08082B099",
  8635 => x"C0C0C0C08082B092",
  8636 => x"C0C0C0C08082B082",
  8637 => x"C0C0C0C08082B0F8",
  8638 => x"C0C0C0C08082B080",
  8639 => x"C0C0C0C08082B090",
  8640 => x"C0C0C0C0808299C0",
  8641 => x"C0C0C0C0808299F9",
  8642 => x"C0C0C0C0808299A4",
  8643 => x"C0C0C0C0808299B0",
  8644 => x"C0C0C0C080829999",
  8645 => x"C0C0C0C080829992",
  8646 => x"C0C0C0C080829982",
  8647 => x"C0C0C0C0808299F8",
  8648 => x"C0C0C0C080829980",
  8649 => x"C0C0C0C080829990",
  8650 => x"C0C0C0C0808292C0",
  8651 => x"C0C0C0C0808292F9",
  8652 => x"C0C0C0C0808292A4",
  8653 => x"C0C0C0C0808292B0",
  8654 => x"C0C0C0C080829299",
  8655 => x"C0C0C0C080829292",
  8656 => x"C0C0C0C080829282",
  8657 => x"C0C0C0C0808292F8",
  8658 => x"C0C0C0C080829280",
  8659 => x"C0C0C0C080829290",
  8660 => x"C0C0C0C0808282C0",
  8661 => x"C0C0C0C0808282F9",
  8662 => x"C0C0C0C0808282A4",
  8663 => x"C0C0C0C0808282B0",
  8664 => x"C0C0C0C080828299",
  8665 => x"C0C0C0C080828292",
  8666 => x"C0C0C0C080828282",
  8667 => x"C0C0C0C0808282F8",
  8668 => x"C0C0C0C080828280",
  8669 => x"C0C0C0C080828290",
  8670 => x"C0C0C0C08082F8C0",
  8671 => x"C0C0C0C08082F8F9",
  8672 => x"C0C0C0C08082F8A4",
  8673 => x"C0C0C0C08082F8B0",
  8674 => x"C0C0C0C08082F899",
  8675 => x"C0C0C0C08082F892",
  8676 => x"C0C0C0C08082F882",
  8677 => x"C0C0C0C08082F8F8",
  8678 => x"C0C0C0C08082F880",
  8679 => x"C0C0C0C08082F890",
  8680 => x"C0C0C0C0808280C0",
  8681 => x"C0C0C0C0808280F9",
  8682 => x"C0C0C0C0808280A4",
  8683 => x"C0C0C0C0808280B0",
  8684 => x"C0C0C0C080828099",
  8685 => x"C0C0C0C080828092",
  8686 => x"C0C0C0C080828082",
  8687 => x"C0C0C0C0808280F8",
  8688 => x"C0C0C0C080828080",
  8689 => x"C0C0C0C080828090",
  8690 => x"C0C0C0C0808290C0",
  8691 => x"C0C0C0C0808290F9",
  8692 => x"C0C0C0C0808290A4",
  8693 => x"C0C0C0C0808290B0",
  8694 => x"C0C0C0C080829099",
  8695 => x"C0C0C0C080829092",
  8696 => x"C0C0C0C080829082",
  8697 => x"C0C0C0C0808290F8",
  8698 => x"C0C0C0C080829080",
  8699 => x"C0C0C0C080829090",
  8700 => x"C0C0C0C080F8C0C0",
  8701 => x"C0C0C0C080F8C0F9",
  8702 => x"C0C0C0C080F8C0A4",
  8703 => x"C0C0C0C080F8C0B0",
  8704 => x"C0C0C0C080F8C099",
  8705 => x"C0C0C0C080F8C092",
  8706 => x"C0C0C0C080F8C082",
  8707 => x"C0C0C0C080F8C0F8",
  8708 => x"C0C0C0C080F8C080",
  8709 => x"C0C0C0C080F8C090",
  8710 => x"C0C0C0C080F8F9C0",
  8711 => x"C0C0C0C080F8F9F9",
  8712 => x"C0C0C0C080F8F9A4",
  8713 => x"C0C0C0C080F8F9B0",
  8714 => x"C0C0C0C080F8F999",
  8715 => x"C0C0C0C080F8F992",
  8716 => x"C0C0C0C080F8F982",
  8717 => x"C0C0C0C080F8F9F8",
  8718 => x"C0C0C0C080F8F980",
  8719 => x"C0C0C0C080F8F990",
  8720 => x"C0C0C0C080F8A4C0",
  8721 => x"C0C0C0C080F8A4F9",
  8722 => x"C0C0C0C080F8A4A4",
  8723 => x"C0C0C0C080F8A4B0",
  8724 => x"C0C0C0C080F8A499",
  8725 => x"C0C0C0C080F8A492",
  8726 => x"C0C0C0C080F8A482",
  8727 => x"C0C0C0C080F8A4F8",
  8728 => x"C0C0C0C080F8A480",
  8729 => x"C0C0C0C080F8A490",
  8730 => x"C0C0C0C080F8B0C0",
  8731 => x"C0C0C0C080F8B0F9",
  8732 => x"C0C0C0C080F8B0A4",
  8733 => x"C0C0C0C080F8B0B0",
  8734 => x"C0C0C0C080F8B099",
  8735 => x"C0C0C0C080F8B092",
  8736 => x"C0C0C0C080F8B082",
  8737 => x"C0C0C0C080F8B0F8",
  8738 => x"C0C0C0C080F8B080",
  8739 => x"C0C0C0C080F8B090",
  8740 => x"C0C0C0C080F899C0",
  8741 => x"C0C0C0C080F899F9",
  8742 => x"C0C0C0C080F899A4",
  8743 => x"C0C0C0C080F899B0",
  8744 => x"C0C0C0C080F89999",
  8745 => x"C0C0C0C080F89992",
  8746 => x"C0C0C0C080F89982",
  8747 => x"C0C0C0C080F899F8",
  8748 => x"C0C0C0C080F89980",
  8749 => x"C0C0C0C080F89990",
  8750 => x"C0C0C0C080F892C0",
  8751 => x"C0C0C0C080F892F9",
  8752 => x"C0C0C0C080F892A4",
  8753 => x"C0C0C0C080F892B0",
  8754 => x"C0C0C0C080F89299",
  8755 => x"C0C0C0C080F89292",
  8756 => x"C0C0C0C080F89282",
  8757 => x"C0C0C0C080F892F8",
  8758 => x"C0C0C0C080F89280",
  8759 => x"C0C0C0C080F89290",
  8760 => x"C0C0C0C080F882C0",
  8761 => x"C0C0C0C080F882F9",
  8762 => x"C0C0C0C080F882A4",
  8763 => x"C0C0C0C080F882B0",
  8764 => x"C0C0C0C080F88299",
  8765 => x"C0C0C0C080F88292",
  8766 => x"C0C0C0C080F88282",
  8767 => x"C0C0C0C080F882F8",
  8768 => x"C0C0C0C080F88280",
  8769 => x"C0C0C0C080F88290",
  8770 => x"C0C0C0C080F8F8C0",
  8771 => x"C0C0C0C080F8F8F9",
  8772 => x"C0C0C0C080F8F8A4",
  8773 => x"C0C0C0C080F8F8B0",
  8774 => x"C0C0C0C080F8F899",
  8775 => x"C0C0C0C080F8F892",
  8776 => x"C0C0C0C080F8F882",
  8777 => x"C0C0C0C080F8F8F8",
  8778 => x"C0C0C0C080F8F880",
  8779 => x"C0C0C0C080F8F890",
  8780 => x"C0C0C0C080F880C0",
  8781 => x"C0C0C0C080F880F9",
  8782 => x"C0C0C0C080F880A4",
  8783 => x"C0C0C0C080F880B0",
  8784 => x"C0C0C0C080F88099",
  8785 => x"C0C0C0C080F88092",
  8786 => x"C0C0C0C080F88082",
  8787 => x"C0C0C0C080F880F8",
  8788 => x"C0C0C0C080F88080",
  8789 => x"C0C0C0C080F88090",
  8790 => x"C0C0C0C080F890C0",
  8791 => x"C0C0C0C080F890F9",
  8792 => x"C0C0C0C080F890A4",
  8793 => x"C0C0C0C080F890B0",
  8794 => x"C0C0C0C080F89099",
  8795 => x"C0C0C0C080F89092",
  8796 => x"C0C0C0C080F89082",
  8797 => x"C0C0C0C080F890F8",
  8798 => x"C0C0C0C080F89080",
  8799 => x"C0C0C0C080F89090",
  8800 => x"C0C0C0C08080C0C0",
  8801 => x"C0C0C0C08080C0F9",
  8802 => x"C0C0C0C08080C0A4",
  8803 => x"C0C0C0C08080C0B0",
  8804 => x"C0C0C0C08080C099",
  8805 => x"C0C0C0C08080C092",
  8806 => x"C0C0C0C08080C082",
  8807 => x"C0C0C0C08080C0F8",
  8808 => x"C0C0C0C08080C080",
  8809 => x"C0C0C0C08080C090",
  8810 => x"C0C0C0C08080F9C0",
  8811 => x"C0C0C0C08080F9F9",
  8812 => x"C0C0C0C08080F9A4",
  8813 => x"C0C0C0C08080F9B0",
  8814 => x"C0C0C0C08080F999",
  8815 => x"C0C0C0C08080F992",
  8816 => x"C0C0C0C08080F982",
  8817 => x"C0C0C0C08080F9F8",
  8818 => x"C0C0C0C08080F980",
  8819 => x"C0C0C0C08080F990",
  8820 => x"C0C0C0C08080A4C0",
  8821 => x"C0C0C0C08080A4F9",
  8822 => x"C0C0C0C08080A4A4",
  8823 => x"C0C0C0C08080A4B0",
  8824 => x"C0C0C0C08080A499",
  8825 => x"C0C0C0C08080A492",
  8826 => x"C0C0C0C08080A482",
  8827 => x"C0C0C0C08080A4F8",
  8828 => x"C0C0C0C08080A480",
  8829 => x"C0C0C0C08080A490",
  8830 => x"C0C0C0C08080B0C0",
  8831 => x"C0C0C0C08080B0F9",
  8832 => x"C0C0C0C08080B0A4",
  8833 => x"C0C0C0C08080B0B0",
  8834 => x"C0C0C0C08080B099",
  8835 => x"C0C0C0C08080B092",
  8836 => x"C0C0C0C08080B082",
  8837 => x"C0C0C0C08080B0F8",
  8838 => x"C0C0C0C08080B080",
  8839 => x"C0C0C0C08080B090",
  8840 => x"C0C0C0C0808099C0",
  8841 => x"C0C0C0C0808099F9",
  8842 => x"C0C0C0C0808099A4",
  8843 => x"C0C0C0C0808099B0",
  8844 => x"C0C0C0C080809999",
  8845 => x"C0C0C0C080809992",
  8846 => x"C0C0C0C080809982",
  8847 => x"C0C0C0C0808099F8",
  8848 => x"C0C0C0C080809980",
  8849 => x"C0C0C0C080809990",
  8850 => x"C0C0C0C0808092C0",
  8851 => x"C0C0C0C0808092F9",
  8852 => x"C0C0C0C0808092A4",
  8853 => x"C0C0C0C0808092B0",
  8854 => x"C0C0C0C080809299",
  8855 => x"C0C0C0C080809292",
  8856 => x"C0C0C0C080809282",
  8857 => x"C0C0C0C0808092F8",
  8858 => x"C0C0C0C080809280",
  8859 => x"C0C0C0C080809290",
  8860 => x"C0C0C0C0808082C0",
  8861 => x"C0C0C0C0808082F9",
  8862 => x"C0C0C0C0808082A4",
  8863 => x"C0C0C0C0808082B0",
  8864 => x"C0C0C0C080808299",
  8865 => x"C0C0C0C080808292",
  8866 => x"C0C0C0C080808282",
  8867 => x"C0C0C0C0808082F8",
  8868 => x"C0C0C0C080808280",
  8869 => x"C0C0C0C080808290",
  8870 => x"C0C0C0C08080F8C0",
  8871 => x"C0C0C0C08080F8F9",
  8872 => x"C0C0C0C08080F8A4",
  8873 => x"C0C0C0C08080F8B0",
  8874 => x"C0C0C0C08080F899",
  8875 => x"C0C0C0C08080F892",
  8876 => x"C0C0C0C08080F882",
  8877 => x"C0C0C0C08080F8F8",
  8878 => x"C0C0C0C08080F880",
  8879 => x"C0C0C0C08080F890",
  8880 => x"C0C0C0C0808080C0",
  8881 => x"C0C0C0C0808080F9",
  8882 => x"C0C0C0C0808080A4",
  8883 => x"C0C0C0C0808080B0",
  8884 => x"C0C0C0C080808099",
  8885 => x"C0C0C0C080808092",
  8886 => x"C0C0C0C080808082",
  8887 => x"C0C0C0C0808080F8",
  8888 => x"C0C0C0C080808080",
  8889 => x"C0C0C0C080808090",
  8890 => x"C0C0C0C0808090C0",
  8891 => x"C0C0C0C0808090F9",
  8892 => x"C0C0C0C0808090A4",
  8893 => x"C0C0C0C0808090B0",
  8894 => x"C0C0C0C080809099",
  8895 => x"C0C0C0C080809092",
  8896 => x"C0C0C0C080809082",
  8897 => x"C0C0C0C0808090F8",
  8898 => x"C0C0C0C080809080",
  8899 => x"C0C0C0C080809090",
  8900 => x"C0C0C0C08090C0C0",
  8901 => x"C0C0C0C08090C0F9",
  8902 => x"C0C0C0C08090C0A4",
  8903 => x"C0C0C0C08090C0B0",
  8904 => x"C0C0C0C08090C099",
  8905 => x"C0C0C0C08090C092",
  8906 => x"C0C0C0C08090C082",
  8907 => x"C0C0C0C08090C0F8",
  8908 => x"C0C0C0C08090C080",
  8909 => x"C0C0C0C08090C090",
  8910 => x"C0C0C0C08090F9C0",
  8911 => x"C0C0C0C08090F9F9",
  8912 => x"C0C0C0C08090F9A4",
  8913 => x"C0C0C0C08090F9B0",
  8914 => x"C0C0C0C08090F999",
  8915 => x"C0C0C0C08090F992",
  8916 => x"C0C0C0C08090F982",
  8917 => x"C0C0C0C08090F9F8",
  8918 => x"C0C0C0C08090F980",
  8919 => x"C0C0C0C08090F990",
  8920 => x"C0C0C0C08090A4C0",
  8921 => x"C0C0C0C08090A4F9",
  8922 => x"C0C0C0C08090A4A4",
  8923 => x"C0C0C0C08090A4B0",
  8924 => x"C0C0C0C08090A499",
  8925 => x"C0C0C0C08090A492",
  8926 => x"C0C0C0C08090A482",
  8927 => x"C0C0C0C08090A4F8",
  8928 => x"C0C0C0C08090A480",
  8929 => x"C0C0C0C08090A490",
  8930 => x"C0C0C0C08090B0C0",
  8931 => x"C0C0C0C08090B0F9",
  8932 => x"C0C0C0C08090B0A4",
  8933 => x"C0C0C0C08090B0B0",
  8934 => x"C0C0C0C08090B099",
  8935 => x"C0C0C0C08090B092",
  8936 => x"C0C0C0C08090B082",
  8937 => x"C0C0C0C08090B0F8",
  8938 => x"C0C0C0C08090B080",
  8939 => x"C0C0C0C08090B090",
  8940 => x"C0C0C0C0809099C0",
  8941 => x"C0C0C0C0809099F9",
  8942 => x"C0C0C0C0809099A4",
  8943 => x"C0C0C0C0809099B0",
  8944 => x"C0C0C0C080909999",
  8945 => x"C0C0C0C080909992",
  8946 => x"C0C0C0C080909982",
  8947 => x"C0C0C0C0809099F8",
  8948 => x"C0C0C0C080909980",
  8949 => x"C0C0C0C080909990",
  8950 => x"C0C0C0C0809092C0",
  8951 => x"C0C0C0C0809092F9",
  8952 => x"C0C0C0C0809092A4",
  8953 => x"C0C0C0C0809092B0",
  8954 => x"C0C0C0C080909299",
  8955 => x"C0C0C0C080909292",
  8956 => x"C0C0C0C080909282",
  8957 => x"C0C0C0C0809092F8",
  8958 => x"C0C0C0C080909280",
  8959 => x"C0C0C0C080909290",
  8960 => x"C0C0C0C0809082C0",
  8961 => x"C0C0C0C0809082F9",
  8962 => x"C0C0C0C0809082A4",
  8963 => x"C0C0C0C0809082B0",
  8964 => x"C0C0C0C080908299",
  8965 => x"C0C0C0C080908292",
  8966 => x"C0C0C0C080908282",
  8967 => x"C0C0C0C0809082F8",
  8968 => x"C0C0C0C080908280",
  8969 => x"C0C0C0C080908290",
  8970 => x"C0C0C0C08090F8C0",
  8971 => x"C0C0C0C08090F8F9",
  8972 => x"C0C0C0C08090F8A4",
  8973 => x"C0C0C0C08090F8B0",
  8974 => x"C0C0C0C08090F899",
  8975 => x"C0C0C0C08090F892",
  8976 => x"C0C0C0C08090F882",
  8977 => x"C0C0C0C08090F8F8",
  8978 => x"C0C0C0C08090F880",
  8979 => x"C0C0C0C08090F890",
  8980 => x"C0C0C0C0809080C0",
  8981 => x"C0C0C0C0809080F9",
  8982 => x"C0C0C0C0809080A4",
  8983 => x"C0C0C0C0809080B0",
  8984 => x"C0C0C0C080908099",
  8985 => x"C0C0C0C080908092",
  8986 => x"C0C0C0C080908082",
  8987 => x"C0C0C0C0809080F8",
  8988 => x"C0C0C0C080908080",
  8989 => x"C0C0C0C080908090",
  8990 => x"C0C0C0C0809090C0",
  8991 => x"C0C0C0C0809090F9",
  8992 => x"C0C0C0C0809090A4",
  8993 => x"C0C0C0C0809090B0",
  8994 => x"C0C0C0C080909099",
  8995 => x"C0C0C0C080909092",
  8996 => x"C0C0C0C080909082",
  8997 => x"C0C0C0C0809090F8",
  8998 => x"C0C0C0C080909080",
  8999 => x"C0C0C0C080909090",
  9000 => x"C0C0C0C090C0C0C0",
  9001 => x"C0C0C0C090C0C0F9",
  9002 => x"C0C0C0C090C0C0A4",
  9003 => x"C0C0C0C090C0C0B0",
  9004 => x"C0C0C0C090C0C099",
  9005 => x"C0C0C0C090C0C092",
  9006 => x"C0C0C0C090C0C082",
  9007 => x"C0C0C0C090C0C0F8",
  9008 => x"C0C0C0C090C0C080",
  9009 => x"C0C0C0C090C0C090",
  9010 => x"C0C0C0C090C0F9C0",
  9011 => x"C0C0C0C090C0F9F9",
  9012 => x"C0C0C0C090C0F9A4",
  9013 => x"C0C0C0C090C0F9B0",
  9014 => x"C0C0C0C090C0F999",
  9015 => x"C0C0C0C090C0F992",
  9016 => x"C0C0C0C090C0F982",
  9017 => x"C0C0C0C090C0F9F8",
  9018 => x"C0C0C0C090C0F980",
  9019 => x"C0C0C0C090C0F990",
  9020 => x"C0C0C0C090C0A4C0",
  9021 => x"C0C0C0C090C0A4F9",
  9022 => x"C0C0C0C090C0A4A4",
  9023 => x"C0C0C0C090C0A4B0",
  9024 => x"C0C0C0C090C0A499",
  9025 => x"C0C0C0C090C0A492",
  9026 => x"C0C0C0C090C0A482",
  9027 => x"C0C0C0C090C0A4F8",
  9028 => x"C0C0C0C090C0A480",
  9029 => x"C0C0C0C090C0A490",
  9030 => x"C0C0C0C090C0B0C0",
  9031 => x"C0C0C0C090C0B0F9",
  9032 => x"C0C0C0C090C0B0A4",
  9033 => x"C0C0C0C090C0B0B0",
  9034 => x"C0C0C0C090C0B099",
  9035 => x"C0C0C0C090C0B092",
  9036 => x"C0C0C0C090C0B082",
  9037 => x"C0C0C0C090C0B0F8",
  9038 => x"C0C0C0C090C0B080",
  9039 => x"C0C0C0C090C0B090",
  9040 => x"C0C0C0C090C099C0",
  9041 => x"C0C0C0C090C099F9",
  9042 => x"C0C0C0C090C099A4",
  9043 => x"C0C0C0C090C099B0",
  9044 => x"C0C0C0C090C09999",
  9045 => x"C0C0C0C090C09992",
  9046 => x"C0C0C0C090C09982",
  9047 => x"C0C0C0C090C099F8",
  9048 => x"C0C0C0C090C09980",
  9049 => x"C0C0C0C090C09990",
  9050 => x"C0C0C0C090C092C0",
  9051 => x"C0C0C0C090C092F9",
  9052 => x"C0C0C0C090C092A4",
  9053 => x"C0C0C0C090C092B0",
  9054 => x"C0C0C0C090C09299",
  9055 => x"C0C0C0C090C09292",
  9056 => x"C0C0C0C090C09282",
  9057 => x"C0C0C0C090C092F8",
  9058 => x"C0C0C0C090C09280",
  9059 => x"C0C0C0C090C09290",
  9060 => x"C0C0C0C090C082C0",
  9061 => x"C0C0C0C090C082F9",
  9062 => x"C0C0C0C090C082A4",
  9063 => x"C0C0C0C090C082B0",
  9064 => x"C0C0C0C090C08299",
  9065 => x"C0C0C0C090C08292",
  9066 => x"C0C0C0C090C08282",
  9067 => x"C0C0C0C090C082F8",
  9068 => x"C0C0C0C090C08280",
  9069 => x"C0C0C0C090C08290",
  9070 => x"C0C0C0C090C0F8C0",
  9071 => x"C0C0C0C090C0F8F9",
  9072 => x"C0C0C0C090C0F8A4",
  9073 => x"C0C0C0C090C0F8B0",
  9074 => x"C0C0C0C090C0F899",
  9075 => x"C0C0C0C090C0F892",
  9076 => x"C0C0C0C090C0F882",
  9077 => x"C0C0C0C090C0F8F8",
  9078 => x"C0C0C0C090C0F880",
  9079 => x"C0C0C0C090C0F890",
  9080 => x"C0C0C0C090C080C0",
  9081 => x"C0C0C0C090C080F9",
  9082 => x"C0C0C0C090C080A4",
  9083 => x"C0C0C0C090C080B0",
  9084 => x"C0C0C0C090C08099",
  9085 => x"C0C0C0C090C08092",
  9086 => x"C0C0C0C090C08082",
  9087 => x"C0C0C0C090C080F8",
  9088 => x"C0C0C0C090C08080",
  9089 => x"C0C0C0C090C08090",
  9090 => x"C0C0C0C090C090C0",
  9091 => x"C0C0C0C090C090F9",
  9092 => x"C0C0C0C090C090A4",
  9093 => x"C0C0C0C090C090B0",
  9094 => x"C0C0C0C090C09099",
  9095 => x"C0C0C0C090C09092",
  9096 => x"C0C0C0C090C09082",
  9097 => x"C0C0C0C090C090F8",
  9098 => x"C0C0C0C090C09080",
  9099 => x"C0C0C0C090C09090",
  9100 => x"C0C0C0C090F9C0C0",
  9101 => x"C0C0C0C090F9C0F9",
  9102 => x"C0C0C0C090F9C0A4",
  9103 => x"C0C0C0C090F9C0B0",
  9104 => x"C0C0C0C090F9C099",
  9105 => x"C0C0C0C090F9C092",
  9106 => x"C0C0C0C090F9C082",
  9107 => x"C0C0C0C090F9C0F8",
  9108 => x"C0C0C0C090F9C080",
  9109 => x"C0C0C0C090F9C090",
  9110 => x"C0C0C0C090F9F9C0",
  9111 => x"C0C0C0C090F9F9F9",
  9112 => x"C0C0C0C090F9F9A4",
  9113 => x"C0C0C0C090F9F9B0",
  9114 => x"C0C0C0C090F9F999",
  9115 => x"C0C0C0C090F9F992",
  9116 => x"C0C0C0C090F9F982",
  9117 => x"C0C0C0C090F9F9F8",
  9118 => x"C0C0C0C090F9F980",
  9119 => x"C0C0C0C090F9F990",
  9120 => x"C0C0C0C090F9A4C0",
  9121 => x"C0C0C0C090F9A4F9",
  9122 => x"C0C0C0C090F9A4A4",
  9123 => x"C0C0C0C090F9A4B0",
  9124 => x"C0C0C0C090F9A499",
  9125 => x"C0C0C0C090F9A492",
  9126 => x"C0C0C0C090F9A482",
  9127 => x"C0C0C0C090F9A4F8",
  9128 => x"C0C0C0C090F9A480",
  9129 => x"C0C0C0C090F9A490",
  9130 => x"C0C0C0C090F9B0C0",
  9131 => x"C0C0C0C090F9B0F9",
  9132 => x"C0C0C0C090F9B0A4",
  9133 => x"C0C0C0C090F9B0B0",
  9134 => x"C0C0C0C090F9B099",
  9135 => x"C0C0C0C090F9B092",
  9136 => x"C0C0C0C090F9B082",
  9137 => x"C0C0C0C090F9B0F8",
  9138 => x"C0C0C0C090F9B080",
  9139 => x"C0C0C0C090F9B090",
  9140 => x"C0C0C0C090F999C0",
  9141 => x"C0C0C0C090F999F9",
  9142 => x"C0C0C0C090F999A4",
  9143 => x"C0C0C0C090F999B0",
  9144 => x"C0C0C0C090F99999",
  9145 => x"C0C0C0C090F99992",
  9146 => x"C0C0C0C090F99982",
  9147 => x"C0C0C0C090F999F8",
  9148 => x"C0C0C0C090F99980",
  9149 => x"C0C0C0C090F99990",
  9150 => x"C0C0C0C090F992C0",
  9151 => x"C0C0C0C090F992F9",
  9152 => x"C0C0C0C090F992A4",
  9153 => x"C0C0C0C090F992B0",
  9154 => x"C0C0C0C090F99299",
  9155 => x"C0C0C0C090F99292",
  9156 => x"C0C0C0C090F99282",
  9157 => x"C0C0C0C090F992F8",
  9158 => x"C0C0C0C090F99280",
  9159 => x"C0C0C0C090F99290",
  9160 => x"C0C0C0C090F982C0",
  9161 => x"C0C0C0C090F982F9",
  9162 => x"C0C0C0C090F982A4",
  9163 => x"C0C0C0C090F982B0",
  9164 => x"C0C0C0C090F98299",
  9165 => x"C0C0C0C090F98292",
  9166 => x"C0C0C0C090F98282",
  9167 => x"C0C0C0C090F982F8",
  9168 => x"C0C0C0C090F98280",
  9169 => x"C0C0C0C090F98290",
  9170 => x"C0C0C0C090F9F8C0",
  9171 => x"C0C0C0C090F9F8F9",
  9172 => x"C0C0C0C090F9F8A4",
  9173 => x"C0C0C0C090F9F8B0",
  9174 => x"C0C0C0C090F9F899",
  9175 => x"C0C0C0C090F9F892",
  9176 => x"C0C0C0C090F9F882",
  9177 => x"C0C0C0C090F9F8F8",
  9178 => x"C0C0C0C090F9F880",
  9179 => x"C0C0C0C090F9F890",
  9180 => x"C0C0C0C090F980C0",
  9181 => x"C0C0C0C090F980F9",
  9182 => x"C0C0C0C090F980A4",
  9183 => x"C0C0C0C090F980B0",
  9184 => x"C0C0C0C090F98099",
  9185 => x"C0C0C0C090F98092",
  9186 => x"C0C0C0C090F98082",
  9187 => x"C0C0C0C090F980F8",
  9188 => x"C0C0C0C090F98080",
  9189 => x"C0C0C0C090F98090",
  9190 => x"C0C0C0C090F990C0",
  9191 => x"C0C0C0C090F990F9",
  9192 => x"C0C0C0C090F990A4",
  9193 => x"C0C0C0C090F990B0",
  9194 => x"C0C0C0C090F99099",
  9195 => x"C0C0C0C090F99092",
  9196 => x"C0C0C0C090F99082",
  9197 => x"C0C0C0C090F990F8",
  9198 => x"C0C0C0C090F99080",
  9199 => x"C0C0C0C090F99090",
  9200 => x"C0C0C0C090A4C0C0",
  9201 => x"C0C0C0C090A4C0F9",
  9202 => x"C0C0C0C090A4C0A4",
  9203 => x"C0C0C0C090A4C0B0",
  9204 => x"C0C0C0C090A4C099",
  9205 => x"C0C0C0C090A4C092",
  9206 => x"C0C0C0C090A4C082",
  9207 => x"C0C0C0C090A4C0F8",
  9208 => x"C0C0C0C090A4C080",
  9209 => x"C0C0C0C090A4C090",
  9210 => x"C0C0C0C090A4F9C0",
  9211 => x"C0C0C0C090A4F9F9",
  9212 => x"C0C0C0C090A4F9A4",
  9213 => x"C0C0C0C090A4F9B0",
  9214 => x"C0C0C0C090A4F999",
  9215 => x"C0C0C0C090A4F992",
  9216 => x"C0C0C0C090A4F982",
  9217 => x"C0C0C0C090A4F9F8",
  9218 => x"C0C0C0C090A4F980",
  9219 => x"C0C0C0C090A4F990",
  9220 => x"C0C0C0C090A4A4C0",
  9221 => x"C0C0C0C090A4A4F9",
  9222 => x"C0C0C0C090A4A4A4",
  9223 => x"C0C0C0C090A4A4B0",
  9224 => x"C0C0C0C090A4A499",
  9225 => x"C0C0C0C090A4A492",
  9226 => x"C0C0C0C090A4A482",
  9227 => x"C0C0C0C090A4A4F8",
  9228 => x"C0C0C0C090A4A480",
  9229 => x"C0C0C0C090A4A490",
  9230 => x"C0C0C0C090A4B0C0",
  9231 => x"C0C0C0C090A4B0F9",
  9232 => x"C0C0C0C090A4B0A4",
  9233 => x"C0C0C0C090A4B0B0",
  9234 => x"C0C0C0C090A4B099",
  9235 => x"C0C0C0C090A4B092",
  9236 => x"C0C0C0C090A4B082",
  9237 => x"C0C0C0C090A4B0F8",
  9238 => x"C0C0C0C090A4B080",
  9239 => x"C0C0C0C090A4B090",
  9240 => x"C0C0C0C090A499C0",
  9241 => x"C0C0C0C090A499F9",
  9242 => x"C0C0C0C090A499A4",
  9243 => x"C0C0C0C090A499B0",
  9244 => x"C0C0C0C090A49999",
  9245 => x"C0C0C0C090A49992",
  9246 => x"C0C0C0C090A49982",
  9247 => x"C0C0C0C090A499F8",
  9248 => x"C0C0C0C090A49980",
  9249 => x"C0C0C0C090A49990",
  9250 => x"C0C0C0C090A492C0",
  9251 => x"C0C0C0C090A492F9",
  9252 => x"C0C0C0C090A492A4",
  9253 => x"C0C0C0C090A492B0",
  9254 => x"C0C0C0C090A49299",
  9255 => x"C0C0C0C090A49292",
  9256 => x"C0C0C0C090A49282",
  9257 => x"C0C0C0C090A492F8",
  9258 => x"C0C0C0C090A49280",
  9259 => x"C0C0C0C090A49290",
  9260 => x"C0C0C0C090A482C0",
  9261 => x"C0C0C0C090A482F9",
  9262 => x"C0C0C0C090A482A4",
  9263 => x"C0C0C0C090A482B0",
  9264 => x"C0C0C0C090A48299",
  9265 => x"C0C0C0C090A48292",
  9266 => x"C0C0C0C090A48282",
  9267 => x"C0C0C0C090A482F8",
  9268 => x"C0C0C0C090A48280",
  9269 => x"C0C0C0C090A48290",
  9270 => x"C0C0C0C090A4F8C0",
  9271 => x"C0C0C0C090A4F8F9",
  9272 => x"C0C0C0C090A4F8A4",
  9273 => x"C0C0C0C090A4F8B0",
  9274 => x"C0C0C0C090A4F899",
  9275 => x"C0C0C0C090A4F892",
  9276 => x"C0C0C0C090A4F882",
  9277 => x"C0C0C0C090A4F8F8",
  9278 => x"C0C0C0C090A4F880",
  9279 => x"C0C0C0C090A4F890",
  9280 => x"C0C0C0C090A480C0",
  9281 => x"C0C0C0C090A480F9",
  9282 => x"C0C0C0C090A480A4",
  9283 => x"C0C0C0C090A480B0",
  9284 => x"C0C0C0C090A48099",
  9285 => x"C0C0C0C090A48092",
  9286 => x"C0C0C0C090A48082",
  9287 => x"C0C0C0C090A480F8",
  9288 => x"C0C0C0C090A48080",
  9289 => x"C0C0C0C090A48090",
  9290 => x"C0C0C0C090A490C0",
  9291 => x"C0C0C0C090A490F9",
  9292 => x"C0C0C0C090A490A4",
  9293 => x"C0C0C0C090A490B0",
  9294 => x"C0C0C0C090A49099",
  9295 => x"C0C0C0C090A49092",
  9296 => x"C0C0C0C090A49082",
  9297 => x"C0C0C0C090A490F8",
  9298 => x"C0C0C0C090A49080",
  9299 => x"C0C0C0C090A49090",
  9300 => x"C0C0C0C090B0C0C0",
  9301 => x"C0C0C0C090B0C0F9",
  9302 => x"C0C0C0C090B0C0A4",
  9303 => x"C0C0C0C090B0C0B0",
  9304 => x"C0C0C0C090B0C099",
  9305 => x"C0C0C0C090B0C092",
  9306 => x"C0C0C0C090B0C082",
  9307 => x"C0C0C0C090B0C0F8",
  9308 => x"C0C0C0C090B0C080",
  9309 => x"C0C0C0C090B0C090",
  9310 => x"C0C0C0C090B0F9C0",
  9311 => x"C0C0C0C090B0F9F9",
  9312 => x"C0C0C0C090B0F9A4",
  9313 => x"C0C0C0C090B0F9B0",
  9314 => x"C0C0C0C090B0F999",
  9315 => x"C0C0C0C090B0F992",
  9316 => x"C0C0C0C090B0F982",
  9317 => x"C0C0C0C090B0F9F8",
  9318 => x"C0C0C0C090B0F980",
  9319 => x"C0C0C0C090B0F990",
  9320 => x"C0C0C0C090B0A4C0",
  9321 => x"C0C0C0C090B0A4F9",
  9322 => x"C0C0C0C090B0A4A4",
  9323 => x"C0C0C0C090B0A4B0",
  9324 => x"C0C0C0C090B0A499",
  9325 => x"C0C0C0C090B0A492",
  9326 => x"C0C0C0C090B0A482",
  9327 => x"C0C0C0C090B0A4F8",
  9328 => x"C0C0C0C090B0A480",
  9329 => x"C0C0C0C090B0A490",
  9330 => x"C0C0C0C090B0B0C0",
  9331 => x"C0C0C0C090B0B0F9",
  9332 => x"C0C0C0C090B0B0A4",
  9333 => x"C0C0C0C090B0B0B0",
  9334 => x"C0C0C0C090B0B099",
  9335 => x"C0C0C0C090B0B092",
  9336 => x"C0C0C0C090B0B082",
  9337 => x"C0C0C0C090B0B0F8",
  9338 => x"C0C0C0C090B0B080",
  9339 => x"C0C0C0C090B0B090",
  9340 => x"C0C0C0C090B099C0",
  9341 => x"C0C0C0C090B099F9",
  9342 => x"C0C0C0C090B099A4",
  9343 => x"C0C0C0C090B099B0",
  9344 => x"C0C0C0C090B09999",
  9345 => x"C0C0C0C090B09992",
  9346 => x"C0C0C0C090B09982",
  9347 => x"C0C0C0C090B099F8",
  9348 => x"C0C0C0C090B09980",
  9349 => x"C0C0C0C090B09990",
  9350 => x"C0C0C0C090B092C0",
  9351 => x"C0C0C0C090B092F9",
  9352 => x"C0C0C0C090B092A4",
  9353 => x"C0C0C0C090B092B0",
  9354 => x"C0C0C0C090B09299",
  9355 => x"C0C0C0C090B09292",
  9356 => x"C0C0C0C090B09282",
  9357 => x"C0C0C0C090B092F8",
  9358 => x"C0C0C0C090B09280",
  9359 => x"C0C0C0C090B09290",
  9360 => x"C0C0C0C090B082C0",
  9361 => x"C0C0C0C090B082F9",
  9362 => x"C0C0C0C090B082A4",
  9363 => x"C0C0C0C090B082B0",
  9364 => x"C0C0C0C090B08299",
  9365 => x"C0C0C0C090B08292",
  9366 => x"C0C0C0C090B08282",
  9367 => x"C0C0C0C090B082F8",
  9368 => x"C0C0C0C090B08280",
  9369 => x"C0C0C0C090B08290",
  9370 => x"C0C0C0C090B0F8C0",
  9371 => x"C0C0C0C090B0F8F9",
  9372 => x"C0C0C0C090B0F8A4",
  9373 => x"C0C0C0C090B0F8B0",
  9374 => x"C0C0C0C090B0F899",
  9375 => x"C0C0C0C090B0F892",
  9376 => x"C0C0C0C090B0F882",
  9377 => x"C0C0C0C090B0F8F8",
  9378 => x"C0C0C0C090B0F880",
  9379 => x"C0C0C0C090B0F890",
  9380 => x"C0C0C0C090B080C0",
  9381 => x"C0C0C0C090B080F9",
  9382 => x"C0C0C0C090B080A4",
  9383 => x"C0C0C0C090B080B0",
  9384 => x"C0C0C0C090B08099",
  9385 => x"C0C0C0C090B08092",
  9386 => x"C0C0C0C090B08082",
  9387 => x"C0C0C0C090B080F8",
  9388 => x"C0C0C0C090B08080",
  9389 => x"C0C0C0C090B08090",
  9390 => x"C0C0C0C090B090C0",
  9391 => x"C0C0C0C090B090F9",
  9392 => x"C0C0C0C090B090A4",
  9393 => x"C0C0C0C090B090B0",
  9394 => x"C0C0C0C090B09099",
  9395 => x"C0C0C0C090B09092",
  9396 => x"C0C0C0C090B09082",
  9397 => x"C0C0C0C090B090F8",
  9398 => x"C0C0C0C090B09080",
  9399 => x"C0C0C0C090B09090",
  9400 => x"C0C0C0C09099C0C0",
  9401 => x"C0C0C0C09099C0F9",
  9402 => x"C0C0C0C09099C0A4",
  9403 => x"C0C0C0C09099C0B0",
  9404 => x"C0C0C0C09099C099",
  9405 => x"C0C0C0C09099C092",
  9406 => x"C0C0C0C09099C082",
  9407 => x"C0C0C0C09099C0F8",
  9408 => x"C0C0C0C09099C080",
  9409 => x"C0C0C0C09099C090",
  9410 => x"C0C0C0C09099F9C0",
  9411 => x"C0C0C0C09099F9F9",
  9412 => x"C0C0C0C09099F9A4",
  9413 => x"C0C0C0C09099F9B0",
  9414 => x"C0C0C0C09099F999",
  9415 => x"C0C0C0C09099F992",
  9416 => x"C0C0C0C09099F982",
  9417 => x"C0C0C0C09099F9F8",
  9418 => x"C0C0C0C09099F980",
  9419 => x"C0C0C0C09099F990",
  9420 => x"C0C0C0C09099A4C0",
  9421 => x"C0C0C0C09099A4F9",
  9422 => x"C0C0C0C09099A4A4",
  9423 => x"C0C0C0C09099A4B0",
  9424 => x"C0C0C0C09099A499",
  9425 => x"C0C0C0C09099A492",
  9426 => x"C0C0C0C09099A482",
  9427 => x"C0C0C0C09099A4F8",
  9428 => x"C0C0C0C09099A480",
  9429 => x"C0C0C0C09099A490",
  9430 => x"C0C0C0C09099B0C0",
  9431 => x"C0C0C0C09099B0F9",
  9432 => x"C0C0C0C09099B0A4",
  9433 => x"C0C0C0C09099B0B0",
  9434 => x"C0C0C0C09099B099",
  9435 => x"C0C0C0C09099B092",
  9436 => x"C0C0C0C09099B082",
  9437 => x"C0C0C0C09099B0F8",
  9438 => x"C0C0C0C09099B080",
  9439 => x"C0C0C0C09099B090",
  9440 => x"C0C0C0C0909999C0",
  9441 => x"C0C0C0C0909999F9",
  9442 => x"C0C0C0C0909999A4",
  9443 => x"C0C0C0C0909999B0",
  9444 => x"C0C0C0C090999999",
  9445 => x"C0C0C0C090999992",
  9446 => x"C0C0C0C090999982",
  9447 => x"C0C0C0C0909999F8",
  9448 => x"C0C0C0C090999980",
  9449 => x"C0C0C0C090999990",
  9450 => x"C0C0C0C0909992C0",
  9451 => x"C0C0C0C0909992F9",
  9452 => x"C0C0C0C0909992A4",
  9453 => x"C0C0C0C0909992B0",
  9454 => x"C0C0C0C090999299",
  9455 => x"C0C0C0C090999292",
  9456 => x"C0C0C0C090999282",
  9457 => x"C0C0C0C0909992F8",
  9458 => x"C0C0C0C090999280",
  9459 => x"C0C0C0C090999290",
  9460 => x"C0C0C0C0909982C0",
  9461 => x"C0C0C0C0909982F9",
  9462 => x"C0C0C0C0909982A4",
  9463 => x"C0C0C0C0909982B0",
  9464 => x"C0C0C0C090998299",
  9465 => x"C0C0C0C090998292",
  9466 => x"C0C0C0C090998282",
  9467 => x"C0C0C0C0909982F8",
  9468 => x"C0C0C0C090998280",
  9469 => x"C0C0C0C090998290",
  9470 => x"C0C0C0C09099F8C0",
  9471 => x"C0C0C0C09099F8F9",
  9472 => x"C0C0C0C09099F8A4",
  9473 => x"C0C0C0C09099F8B0",
  9474 => x"C0C0C0C09099F899",
  9475 => x"C0C0C0C09099F892",
  9476 => x"C0C0C0C09099F882",
  9477 => x"C0C0C0C09099F8F8",
  9478 => x"C0C0C0C09099F880",
  9479 => x"C0C0C0C09099F890",
  9480 => x"C0C0C0C0909980C0",
  9481 => x"C0C0C0C0909980F9",
  9482 => x"C0C0C0C0909980A4",
  9483 => x"C0C0C0C0909980B0",
  9484 => x"C0C0C0C090998099",
  9485 => x"C0C0C0C090998092",
  9486 => x"C0C0C0C090998082",
  9487 => x"C0C0C0C0909980F8",
  9488 => x"C0C0C0C090998080",
  9489 => x"C0C0C0C090998090",
  9490 => x"C0C0C0C0909990C0",
  9491 => x"C0C0C0C0909990F9",
  9492 => x"C0C0C0C0909990A4",
  9493 => x"C0C0C0C0909990B0",
  9494 => x"C0C0C0C090999099",
  9495 => x"C0C0C0C090999092",
  9496 => x"C0C0C0C090999082",
  9497 => x"C0C0C0C0909990F8",
  9498 => x"C0C0C0C090999080",
  9499 => x"C0C0C0C090999090",
  9500 => x"C0C0C0C09092C0C0",
  9501 => x"C0C0C0C09092C0F9",
  9502 => x"C0C0C0C09092C0A4",
  9503 => x"C0C0C0C09092C0B0",
  9504 => x"C0C0C0C09092C099",
  9505 => x"C0C0C0C09092C092",
  9506 => x"C0C0C0C09092C082",
  9507 => x"C0C0C0C09092C0F8",
  9508 => x"C0C0C0C09092C080",
  9509 => x"C0C0C0C09092C090",
  9510 => x"C0C0C0C09092F9C0",
  9511 => x"C0C0C0C09092F9F9",
  9512 => x"C0C0C0C09092F9A4",
  9513 => x"C0C0C0C09092F9B0",
  9514 => x"C0C0C0C09092F999",
  9515 => x"C0C0C0C09092F992",
  9516 => x"C0C0C0C09092F982",
  9517 => x"C0C0C0C09092F9F8",
  9518 => x"C0C0C0C09092F980",
  9519 => x"C0C0C0C09092F990",
  9520 => x"C0C0C0C09092A4C0",
  9521 => x"C0C0C0C09092A4F9",
  9522 => x"C0C0C0C09092A4A4",
  9523 => x"C0C0C0C09092A4B0",
  9524 => x"C0C0C0C09092A499",
  9525 => x"C0C0C0C09092A492",
  9526 => x"C0C0C0C09092A482",
  9527 => x"C0C0C0C09092A4F8",
  9528 => x"C0C0C0C09092A480",
  9529 => x"C0C0C0C09092A490",
  9530 => x"C0C0C0C09092B0C0",
  9531 => x"C0C0C0C09092B0F9",
  9532 => x"C0C0C0C09092B0A4",
  9533 => x"C0C0C0C09092B0B0",
  9534 => x"C0C0C0C09092B099",
  9535 => x"C0C0C0C09092B092",
  9536 => x"C0C0C0C09092B082",
  9537 => x"C0C0C0C09092B0F8",
  9538 => x"C0C0C0C09092B080",
  9539 => x"C0C0C0C09092B090",
  9540 => x"C0C0C0C0909299C0",
  9541 => x"C0C0C0C0909299F9",
  9542 => x"C0C0C0C0909299A4",
  9543 => x"C0C0C0C0909299B0",
  9544 => x"C0C0C0C090929999",
  9545 => x"C0C0C0C090929992",
  9546 => x"C0C0C0C090929982",
  9547 => x"C0C0C0C0909299F8",
  9548 => x"C0C0C0C090929980",
  9549 => x"C0C0C0C090929990",
  9550 => x"C0C0C0C0909292C0",
  9551 => x"C0C0C0C0909292F9",
  9552 => x"C0C0C0C0909292A4",
  9553 => x"C0C0C0C0909292B0",
  9554 => x"C0C0C0C090929299",
  9555 => x"C0C0C0C090929292",
  9556 => x"C0C0C0C090929282",
  9557 => x"C0C0C0C0909292F8",
  9558 => x"C0C0C0C090929280",
  9559 => x"C0C0C0C090929290",
  9560 => x"C0C0C0C0909282C0",
  9561 => x"C0C0C0C0909282F9",
  9562 => x"C0C0C0C0909282A4",
  9563 => x"C0C0C0C0909282B0",
  9564 => x"C0C0C0C090928299",
  9565 => x"C0C0C0C090928292",
  9566 => x"C0C0C0C090928282",
  9567 => x"C0C0C0C0909282F8",
  9568 => x"C0C0C0C090928280",
  9569 => x"C0C0C0C090928290",
  9570 => x"C0C0C0C09092F8C0",
  9571 => x"C0C0C0C09092F8F9",
  9572 => x"C0C0C0C09092F8A4",
  9573 => x"C0C0C0C09092F8B0",
  9574 => x"C0C0C0C09092F899",
  9575 => x"C0C0C0C09092F892",
  9576 => x"C0C0C0C09092F882",
  9577 => x"C0C0C0C09092F8F8",
  9578 => x"C0C0C0C09092F880",
  9579 => x"C0C0C0C09092F890",
  9580 => x"C0C0C0C0909280C0",
  9581 => x"C0C0C0C0909280F9",
  9582 => x"C0C0C0C0909280A4",
  9583 => x"C0C0C0C0909280B0",
  9584 => x"C0C0C0C090928099",
  9585 => x"C0C0C0C090928092",
  9586 => x"C0C0C0C090928082",
  9587 => x"C0C0C0C0909280F8",
  9588 => x"C0C0C0C090928080",
  9589 => x"C0C0C0C090928090",
  9590 => x"C0C0C0C0909290C0",
  9591 => x"C0C0C0C0909290F9",
  9592 => x"C0C0C0C0909290A4",
  9593 => x"C0C0C0C0909290B0",
  9594 => x"C0C0C0C090929099",
  9595 => x"C0C0C0C090929092",
  9596 => x"C0C0C0C090929082",
  9597 => x"C0C0C0C0909290F8",
  9598 => x"C0C0C0C090929080",
  9599 => x"C0C0C0C090929090",
  9600 => x"C0C0C0C09082C0C0",
  9601 => x"C0C0C0C09082C0F9",
  9602 => x"C0C0C0C09082C0A4",
  9603 => x"C0C0C0C09082C0B0",
  9604 => x"C0C0C0C09082C099",
  9605 => x"C0C0C0C09082C092",
  9606 => x"C0C0C0C09082C082",
  9607 => x"C0C0C0C09082C0F8",
  9608 => x"C0C0C0C09082C080",
  9609 => x"C0C0C0C09082C090",
  9610 => x"C0C0C0C09082F9C0",
  9611 => x"C0C0C0C09082F9F9",
  9612 => x"C0C0C0C09082F9A4",
  9613 => x"C0C0C0C09082F9B0",
  9614 => x"C0C0C0C09082F999",
  9615 => x"C0C0C0C09082F992",
  9616 => x"C0C0C0C09082F982",
  9617 => x"C0C0C0C09082F9F8",
  9618 => x"C0C0C0C09082F980",
  9619 => x"C0C0C0C09082F990",
  9620 => x"C0C0C0C09082A4C0",
  9621 => x"C0C0C0C09082A4F9",
  9622 => x"C0C0C0C09082A4A4",
  9623 => x"C0C0C0C09082A4B0",
  9624 => x"C0C0C0C09082A499",
  9625 => x"C0C0C0C09082A492",
  9626 => x"C0C0C0C09082A482",
  9627 => x"C0C0C0C09082A4F8",
  9628 => x"C0C0C0C09082A480",
  9629 => x"C0C0C0C09082A490",
  9630 => x"C0C0C0C09082B0C0",
  9631 => x"C0C0C0C09082B0F9",
  9632 => x"C0C0C0C09082B0A4",
  9633 => x"C0C0C0C09082B0B0",
  9634 => x"C0C0C0C09082B099",
  9635 => x"C0C0C0C09082B092",
  9636 => x"C0C0C0C09082B082",
  9637 => x"C0C0C0C09082B0F8",
  9638 => x"C0C0C0C09082B080",
  9639 => x"C0C0C0C09082B090",
  9640 => x"C0C0C0C0908299C0",
  9641 => x"C0C0C0C0908299F9",
  9642 => x"C0C0C0C0908299A4",
  9643 => x"C0C0C0C0908299B0",
  9644 => x"C0C0C0C090829999",
  9645 => x"C0C0C0C090829992",
  9646 => x"C0C0C0C090829982",
  9647 => x"C0C0C0C0908299F8",
  9648 => x"C0C0C0C090829980",
  9649 => x"C0C0C0C090829990",
  9650 => x"C0C0C0C0908292C0",
  9651 => x"C0C0C0C0908292F9",
  9652 => x"C0C0C0C0908292A4",
  9653 => x"C0C0C0C0908292B0",
  9654 => x"C0C0C0C090829299",
  9655 => x"C0C0C0C090829292",
  9656 => x"C0C0C0C090829282",
  9657 => x"C0C0C0C0908292F8",
  9658 => x"C0C0C0C090829280",
  9659 => x"C0C0C0C090829290",
  9660 => x"C0C0C0C0908282C0",
  9661 => x"C0C0C0C0908282F9",
  9662 => x"C0C0C0C0908282A4",
  9663 => x"C0C0C0C0908282B0",
  9664 => x"C0C0C0C090828299",
  9665 => x"C0C0C0C090828292",
  9666 => x"C0C0C0C090828282",
  9667 => x"C0C0C0C0908282F8",
  9668 => x"C0C0C0C090828280",
  9669 => x"C0C0C0C090828290",
  9670 => x"C0C0C0C09082F8C0",
  9671 => x"C0C0C0C09082F8F9",
  9672 => x"C0C0C0C09082F8A4",
  9673 => x"C0C0C0C09082F8B0",
  9674 => x"C0C0C0C09082F899",
  9675 => x"C0C0C0C09082F892",
  9676 => x"C0C0C0C09082F882",
  9677 => x"C0C0C0C09082F8F8",
  9678 => x"C0C0C0C09082F880",
  9679 => x"C0C0C0C09082F890",
  9680 => x"C0C0C0C0908280C0",
  9681 => x"C0C0C0C0908280F9",
  9682 => x"C0C0C0C0908280A4",
  9683 => x"C0C0C0C0908280B0",
  9684 => x"C0C0C0C090828099",
  9685 => x"C0C0C0C090828092",
  9686 => x"C0C0C0C090828082",
  9687 => x"C0C0C0C0908280F8",
  9688 => x"C0C0C0C090828080",
  9689 => x"C0C0C0C090828090",
  9690 => x"C0C0C0C0908290C0",
  9691 => x"C0C0C0C0908290F9",
  9692 => x"C0C0C0C0908290A4",
  9693 => x"C0C0C0C0908290B0",
  9694 => x"C0C0C0C090829099",
  9695 => x"C0C0C0C090829092",
  9696 => x"C0C0C0C090829082",
  9697 => x"C0C0C0C0908290F8",
  9698 => x"C0C0C0C090829080",
  9699 => x"C0C0C0C090829090",
  9700 => x"C0C0C0C090F8C0C0",
  9701 => x"C0C0C0C090F8C0F9",
  9702 => x"C0C0C0C090F8C0A4",
  9703 => x"C0C0C0C090F8C0B0",
  9704 => x"C0C0C0C090F8C099",
  9705 => x"C0C0C0C090F8C092",
  9706 => x"C0C0C0C090F8C082",
  9707 => x"C0C0C0C090F8C0F8",
  9708 => x"C0C0C0C090F8C080",
  9709 => x"C0C0C0C090F8C090",
  9710 => x"C0C0C0C090F8F9C0",
  9711 => x"C0C0C0C090F8F9F9",
  9712 => x"C0C0C0C090F8F9A4",
  9713 => x"C0C0C0C090F8F9B0",
  9714 => x"C0C0C0C090F8F999",
  9715 => x"C0C0C0C090F8F992",
  9716 => x"C0C0C0C090F8F982",
  9717 => x"C0C0C0C090F8F9F8",
  9718 => x"C0C0C0C090F8F980",
  9719 => x"C0C0C0C090F8F990",
  9720 => x"C0C0C0C090F8A4C0",
  9721 => x"C0C0C0C090F8A4F9",
  9722 => x"C0C0C0C090F8A4A4",
  9723 => x"C0C0C0C090F8A4B0",
  9724 => x"C0C0C0C090F8A499",
  9725 => x"C0C0C0C090F8A492",
  9726 => x"C0C0C0C090F8A482",
  9727 => x"C0C0C0C090F8A4F8",
  9728 => x"C0C0C0C090F8A480",
  9729 => x"C0C0C0C090F8A490",
  9730 => x"C0C0C0C090F8B0C0",
  9731 => x"C0C0C0C090F8B0F9",
  9732 => x"C0C0C0C090F8B0A4",
  9733 => x"C0C0C0C090F8B0B0",
  9734 => x"C0C0C0C090F8B099",
  9735 => x"C0C0C0C090F8B092",
  9736 => x"C0C0C0C090F8B082",
  9737 => x"C0C0C0C090F8B0F8",
  9738 => x"C0C0C0C090F8B080",
  9739 => x"C0C0C0C090F8B090",
  9740 => x"C0C0C0C090F899C0",
  9741 => x"C0C0C0C090F899F9",
  9742 => x"C0C0C0C090F899A4",
  9743 => x"C0C0C0C090F899B0",
  9744 => x"C0C0C0C090F89999",
  9745 => x"C0C0C0C090F89992",
  9746 => x"C0C0C0C090F89982",
  9747 => x"C0C0C0C090F899F8",
  9748 => x"C0C0C0C090F89980",
  9749 => x"C0C0C0C090F89990",
  9750 => x"C0C0C0C090F892C0",
  9751 => x"C0C0C0C090F892F9",
  9752 => x"C0C0C0C090F892A4",
  9753 => x"C0C0C0C090F892B0",
  9754 => x"C0C0C0C090F89299",
  9755 => x"C0C0C0C090F89292",
  9756 => x"C0C0C0C090F89282",
  9757 => x"C0C0C0C090F892F8",
  9758 => x"C0C0C0C090F89280",
  9759 => x"C0C0C0C090F89290",
  9760 => x"C0C0C0C090F882C0",
  9761 => x"C0C0C0C090F882F9",
  9762 => x"C0C0C0C090F882A4",
  9763 => x"C0C0C0C090F882B0",
  9764 => x"C0C0C0C090F88299",
  9765 => x"C0C0C0C090F88292",
  9766 => x"C0C0C0C090F88282",
  9767 => x"C0C0C0C090F882F8",
  9768 => x"C0C0C0C090F88280",
  9769 => x"C0C0C0C090F88290",
  9770 => x"C0C0C0C090F8F8C0",
  9771 => x"C0C0C0C090F8F8F9",
  9772 => x"C0C0C0C090F8F8A4",
  9773 => x"C0C0C0C090F8F8B0",
  9774 => x"C0C0C0C090F8F899",
  9775 => x"C0C0C0C090F8F892",
  9776 => x"C0C0C0C090F8F882",
  9777 => x"C0C0C0C090F8F8F8",
  9778 => x"C0C0C0C090F8F880",
  9779 => x"C0C0C0C090F8F890",
  9780 => x"C0C0C0C090F880C0",
  9781 => x"C0C0C0C090F880F9",
  9782 => x"C0C0C0C090F880A4",
  9783 => x"C0C0C0C090F880B0",
  9784 => x"C0C0C0C090F88099",
  9785 => x"C0C0C0C090F88092",
  9786 => x"C0C0C0C090F88082",
  9787 => x"C0C0C0C090F880F8",
  9788 => x"C0C0C0C090F88080",
  9789 => x"C0C0C0C090F88090",
  9790 => x"C0C0C0C090F890C0",
  9791 => x"C0C0C0C090F890F9",
  9792 => x"C0C0C0C090F890A4",
  9793 => x"C0C0C0C090F890B0",
  9794 => x"C0C0C0C090F89099",
  9795 => x"C0C0C0C090F89092",
  9796 => x"C0C0C0C090F89082",
  9797 => x"C0C0C0C090F890F8",
  9798 => x"C0C0C0C090F89080",
  9799 => x"C0C0C0C090F89090",
  9800 => x"C0C0C0C09080C0C0",
  9801 => x"C0C0C0C09080C0F9",
  9802 => x"C0C0C0C09080C0A4",
  9803 => x"C0C0C0C09080C0B0",
  9804 => x"C0C0C0C09080C099",
  9805 => x"C0C0C0C09080C092",
  9806 => x"C0C0C0C09080C082",
  9807 => x"C0C0C0C09080C0F8",
  9808 => x"C0C0C0C09080C080",
  9809 => x"C0C0C0C09080C090",
  9810 => x"C0C0C0C09080F9C0",
  9811 => x"C0C0C0C09080F9F9",
  9812 => x"C0C0C0C09080F9A4",
  9813 => x"C0C0C0C09080F9B0",
  9814 => x"C0C0C0C09080F999",
  9815 => x"C0C0C0C09080F992",
  9816 => x"C0C0C0C09080F982",
  9817 => x"C0C0C0C09080F9F8",
  9818 => x"C0C0C0C09080F980",
  9819 => x"C0C0C0C09080F990",
  9820 => x"C0C0C0C09080A4C0",
  9821 => x"C0C0C0C09080A4F9",
  9822 => x"C0C0C0C09080A4A4",
  9823 => x"C0C0C0C09080A4B0",
  9824 => x"C0C0C0C09080A499",
  9825 => x"C0C0C0C09080A492",
  9826 => x"C0C0C0C09080A482",
  9827 => x"C0C0C0C09080A4F8",
  9828 => x"C0C0C0C09080A480",
  9829 => x"C0C0C0C09080A490",
  9830 => x"C0C0C0C09080B0C0",
  9831 => x"C0C0C0C09080B0F9",
  9832 => x"C0C0C0C09080B0A4",
  9833 => x"C0C0C0C09080B0B0",
  9834 => x"C0C0C0C09080B099",
  9835 => x"C0C0C0C09080B092",
  9836 => x"C0C0C0C09080B082",
  9837 => x"C0C0C0C09080B0F8",
  9838 => x"C0C0C0C09080B080",
  9839 => x"C0C0C0C09080B090",
  9840 => x"C0C0C0C0908099C0",
  9841 => x"C0C0C0C0908099F9",
  9842 => x"C0C0C0C0908099A4",
  9843 => x"C0C0C0C0908099B0",
  9844 => x"C0C0C0C090809999",
  9845 => x"C0C0C0C090809992",
  9846 => x"C0C0C0C090809982",
  9847 => x"C0C0C0C0908099F8",
  9848 => x"C0C0C0C090809980",
  9849 => x"C0C0C0C090809990",
  9850 => x"C0C0C0C0908092C0",
  9851 => x"C0C0C0C0908092F9",
  9852 => x"C0C0C0C0908092A4",
  9853 => x"C0C0C0C0908092B0",
  9854 => x"C0C0C0C090809299",
  9855 => x"C0C0C0C090809292",
  9856 => x"C0C0C0C090809282",
  9857 => x"C0C0C0C0908092F8",
  9858 => x"C0C0C0C090809280",
  9859 => x"C0C0C0C090809290",
  9860 => x"C0C0C0C0908082C0",
  9861 => x"C0C0C0C0908082F9",
  9862 => x"C0C0C0C0908082A4",
  9863 => x"C0C0C0C0908082B0",
  9864 => x"C0C0C0C090808299",
  9865 => x"C0C0C0C090808292",
  9866 => x"C0C0C0C090808282",
  9867 => x"C0C0C0C0908082F8",
  9868 => x"C0C0C0C090808280",
  9869 => x"C0C0C0C090808290",
  9870 => x"C0C0C0C09080F8C0",
  9871 => x"C0C0C0C09080F8F9",
  9872 => x"C0C0C0C09080F8A4",
  9873 => x"C0C0C0C09080F8B0",
  9874 => x"C0C0C0C09080F899",
  9875 => x"C0C0C0C09080F892",
  9876 => x"C0C0C0C09080F882",
  9877 => x"C0C0C0C09080F8F8",
  9878 => x"C0C0C0C09080F880",
  9879 => x"C0C0C0C09080F890",
  9880 => x"C0C0C0C0908080C0",
  9881 => x"C0C0C0C0908080F9",
  9882 => x"C0C0C0C0908080A4",
  9883 => x"C0C0C0C0908080B0",
  9884 => x"C0C0C0C090808099",
  9885 => x"C0C0C0C090808092",
  9886 => x"C0C0C0C090808082",
  9887 => x"C0C0C0C0908080F8",
  9888 => x"C0C0C0C090808080",
  9889 => x"C0C0C0C090808090",
  9890 => x"C0C0C0C0908090C0",
  9891 => x"C0C0C0C0908090F9",
  9892 => x"C0C0C0C0908090A4",
  9893 => x"C0C0C0C0908090B0",
  9894 => x"C0C0C0C090809099",
  9895 => x"C0C0C0C090809092",
  9896 => x"C0C0C0C090809082",
  9897 => x"C0C0C0C0908090F8",
  9898 => x"C0C0C0C090809080",
  9899 => x"C0C0C0C090809090",
  9900 => x"C0C0C0C09090C0C0",
  9901 => x"C0C0C0C09090C0F9",
  9902 => x"C0C0C0C09090C0A4",
  9903 => x"C0C0C0C09090C0B0",
  9904 => x"C0C0C0C09090C099",
  9905 => x"C0C0C0C09090C092",
  9906 => x"C0C0C0C09090C082",
  9907 => x"C0C0C0C09090C0F8",
  9908 => x"C0C0C0C09090C080",
  9909 => x"C0C0C0C09090C090",
  9910 => x"C0C0C0C09090F9C0",
  9911 => x"C0C0C0C09090F9F9",
  9912 => x"C0C0C0C09090F9A4",
  9913 => x"C0C0C0C09090F9B0",
  9914 => x"C0C0C0C09090F999",
  9915 => x"C0C0C0C09090F992",
  9916 => x"C0C0C0C09090F982",
  9917 => x"C0C0C0C09090F9F8",
  9918 => x"C0C0C0C09090F980",
  9919 => x"C0C0C0C09090F990",
  9920 => x"C0C0C0C09090A4C0",
  9921 => x"C0C0C0C09090A4F9",
  9922 => x"C0C0C0C09090A4A4",
  9923 => x"C0C0C0C09090A4B0",
  9924 => x"C0C0C0C09090A499",
  9925 => x"C0C0C0C09090A492",
  9926 => x"C0C0C0C09090A482",
  9927 => x"C0C0C0C09090A4F8",
  9928 => x"C0C0C0C09090A480",
  9929 => x"C0C0C0C09090A490",
  9930 => x"C0C0C0C09090B0C0",
  9931 => x"C0C0C0C09090B0F9",
  9932 => x"C0C0C0C09090B0A4",
  9933 => x"C0C0C0C09090B0B0",
  9934 => x"C0C0C0C09090B099",
  9935 => x"C0C0C0C09090B092",
  9936 => x"C0C0C0C09090B082",
  9937 => x"C0C0C0C09090B0F8",
  9938 => x"C0C0C0C09090B080",
  9939 => x"C0C0C0C09090B090",
  9940 => x"C0C0C0C0909099C0",
  9941 => x"C0C0C0C0909099F9",
  9942 => x"C0C0C0C0909099A4",
  9943 => x"C0C0C0C0909099B0",
  9944 => x"C0C0C0C090909999",
  9945 => x"C0C0C0C090909992",
  9946 => x"C0C0C0C090909982",
  9947 => x"C0C0C0C0909099F8",
  9948 => x"C0C0C0C090909980",
  9949 => x"C0C0C0C090909990",
  9950 => x"C0C0C0C0909092C0",
  9951 => x"C0C0C0C0909092F9",
  9952 => x"C0C0C0C0909092A4",
  9953 => x"C0C0C0C0909092B0",
  9954 => x"C0C0C0C090909299",
  9955 => x"C0C0C0C090909292",
  9956 => x"C0C0C0C090909282",
  9957 => x"C0C0C0C0909092F8",
  9958 => x"C0C0C0C090909280",
  9959 => x"C0C0C0C090909290",
  9960 => x"C0C0C0C0909082C0",
  9961 => x"C0C0C0C0909082F9",
  9962 => x"C0C0C0C0909082A4",
  9963 => x"C0C0C0C0909082B0",
  9964 => x"C0C0C0C090908299",
  9965 => x"C0C0C0C090908292",
  9966 => x"C0C0C0C090908282",
  9967 => x"C0C0C0C0909082F8",
  9968 => x"C0C0C0C090908280",
  9969 => x"C0C0C0C090908290",
  9970 => x"C0C0C0C09090F8C0",
  9971 => x"C0C0C0C09090F8F9",
  9972 => x"C0C0C0C09090F8A4",
  9973 => x"C0C0C0C09090F8B0",
  9974 => x"C0C0C0C09090F899",
  9975 => x"C0C0C0C09090F892",
  9976 => x"C0C0C0C09090F882",
  9977 => x"C0C0C0C09090F8F8",
  9978 => x"C0C0C0C09090F880",
  9979 => x"C0C0C0C09090F890",
  9980 => x"C0C0C0C0909080C0",
  9981 => x"C0C0C0C0909080F9",
  9982 => x"C0C0C0C0909080A4",
  9983 => x"C0C0C0C0909080B0",
  9984 => x"C0C0C0C090908099",
  9985 => x"C0C0C0C090908092",
  9986 => x"C0C0C0C090908082",
  9987 => x"C0C0C0C0909080F8",
  9988 => x"C0C0C0C090908080",
  9989 => x"C0C0C0C090908090",
  9990 => x"C0C0C0C0909090C0",
  9991 => x"C0C0C0C0909090F9",
  9992 => x"C0C0C0C0909090A4",
  9993 => x"C0C0C0C0909090B0",
  9994 => x"C0C0C0C090909099",
  9995 => x"C0C0C0C090909092",
  9996 => x"C0C0C0C090909082",
  9997 => x"C0C0C0C0909090F8",
  9998 => x"C0C0C0C090909080",
  9999 => x"C0C0C0C090909090",
 10000 => x"C0C0C0F9C0C0C0C0",
 10001 => x"C0C0C0F9C0C0C0F9",
 10002 => x"C0C0C0F9C0C0C0A4",
 10003 => x"C0C0C0F9C0C0C0B0",
 10004 => x"C0C0C0F9C0C0C099",
 10005 => x"C0C0C0F9C0C0C092",
 10006 => x"C0C0C0F9C0C0C082",
 10007 => x"C0C0C0F9C0C0C0F8",
 10008 => x"C0C0C0F9C0C0C080",
 10009 => x"C0C0C0F9C0C0C090",
 10010 => x"C0C0C0F9C0C0F9C0",
 10011 => x"C0C0C0F9C0C0F9F9",
 10012 => x"C0C0C0F9C0C0F9A4",
 10013 => x"C0C0C0F9C0C0F9B0",
 10014 => x"C0C0C0F9C0C0F999",
 10015 => x"C0C0C0F9C0C0F992",
 10016 => x"C0C0C0F9C0C0F982",
 10017 => x"C0C0C0F9C0C0F9F8",
 10018 => x"C0C0C0F9C0C0F980",
 10019 => x"C0C0C0F9C0C0F990",
 10020 => x"C0C0C0F9C0C0A4C0",
 10021 => x"C0C0C0F9C0C0A4F9",
 10022 => x"C0C0C0F9C0C0A4A4",
 10023 => x"C0C0C0F9C0C0A4B0",
 10024 => x"C0C0C0F9C0C0A499",
 10025 => x"C0C0C0F9C0C0A492",
 10026 => x"C0C0C0F9C0C0A482",
 10027 => x"C0C0C0F9C0C0A4F8",
 10028 => x"C0C0C0F9C0C0A480",
 10029 => x"C0C0C0F9C0C0A490",
 10030 => x"C0C0C0F9C0C0B0C0",
 10031 => x"C0C0C0F9C0C0B0F9",
 10032 => x"C0C0C0F9C0C0B0A4",
 10033 => x"C0C0C0F9C0C0B0B0",
 10034 => x"C0C0C0F9C0C0B099",
 10035 => x"C0C0C0F9C0C0B092",
 10036 => x"C0C0C0F9C0C0B082",
 10037 => x"C0C0C0F9C0C0B0F8",
 10038 => x"C0C0C0F9C0C0B080",
 10039 => x"C0C0C0F9C0C0B090",
 10040 => x"C0C0C0F9C0C099C0",
 10041 => x"C0C0C0F9C0C099F9",
 10042 => x"C0C0C0F9C0C099A4",
 10043 => x"C0C0C0F9C0C099B0",
 10044 => x"C0C0C0F9C0C09999",
 10045 => x"C0C0C0F9C0C09992",
 10046 => x"C0C0C0F9C0C09982",
 10047 => x"C0C0C0F9C0C099F8",
 10048 => x"C0C0C0F9C0C09980",
 10049 => x"C0C0C0F9C0C09990",
 10050 => x"C0C0C0F9C0C092C0",
 10051 => x"C0C0C0F9C0C092F9",
 10052 => x"C0C0C0F9C0C092A4",
 10053 => x"C0C0C0F9C0C092B0",
 10054 => x"C0C0C0F9C0C09299",
 10055 => x"C0C0C0F9C0C09292",
 10056 => x"C0C0C0F9C0C09282",
 10057 => x"C0C0C0F9C0C092F8",
 10058 => x"C0C0C0F9C0C09280",
 10059 => x"C0C0C0F9C0C09290",
 10060 => x"C0C0C0F9C0C082C0",
 10061 => x"C0C0C0F9C0C082F9",
 10062 => x"C0C0C0F9C0C082A4",
 10063 => x"C0C0C0F9C0C082B0",
 10064 => x"C0C0C0F9C0C08299",
 10065 => x"C0C0C0F9C0C08292",
 10066 => x"C0C0C0F9C0C08282",
 10067 => x"C0C0C0F9C0C082F8",
 10068 => x"C0C0C0F9C0C08280",
 10069 => x"C0C0C0F9C0C08290",
 10070 => x"C0C0C0F9C0C0F8C0",
 10071 => x"C0C0C0F9C0C0F8F9",
 10072 => x"C0C0C0F9C0C0F8A4",
 10073 => x"C0C0C0F9C0C0F8B0",
 10074 => x"C0C0C0F9C0C0F899",
 10075 => x"C0C0C0F9C0C0F892",
 10076 => x"C0C0C0F9C0C0F882",
 10077 => x"C0C0C0F9C0C0F8F8",
 10078 => x"C0C0C0F9C0C0F880",
 10079 => x"C0C0C0F9C0C0F890",
 10080 => x"C0C0C0F9C0C080C0",
 10081 => x"C0C0C0F9C0C080F9",
 10082 => x"C0C0C0F9C0C080A4",
 10083 => x"C0C0C0F9C0C080B0",
 10084 => x"C0C0C0F9C0C08099",
 10085 => x"C0C0C0F9C0C08092",
 10086 => x"C0C0C0F9C0C08082",
 10087 => x"C0C0C0F9C0C080F8",
 10088 => x"C0C0C0F9C0C08080",
 10089 => x"C0C0C0F9C0C08090",
 10090 => x"C0C0C0F9C0C090C0",
 10091 => x"C0C0C0F9C0C090F9",
 10092 => x"C0C0C0F9C0C090A4",
 10093 => x"C0C0C0F9C0C090B0",
 10094 => x"C0C0C0F9C0C09099",
 10095 => x"C0C0C0F9C0C09092",
 10096 => x"C0C0C0F9C0C09082",
 10097 => x"C0C0C0F9C0C090F8",
 10098 => x"C0C0C0F9C0C09080",
 10099 => x"C0C0C0F9C0C09090",
 10100 => x"C0C0C0F9C0F9C0C0",
 10101 => x"C0C0C0F9C0F9C0F9",
 10102 => x"C0C0C0F9C0F9C0A4",
 10103 => x"C0C0C0F9C0F9C0B0",
 10104 => x"C0C0C0F9C0F9C099",
 10105 => x"C0C0C0F9C0F9C092",
 10106 => x"C0C0C0F9C0F9C082",
 10107 => x"C0C0C0F9C0F9C0F8",
 10108 => x"C0C0C0F9C0F9C080",
 10109 => x"C0C0C0F9C0F9C090",
 10110 => x"C0C0C0F9C0F9F9C0",
 10111 => x"C0C0C0F9C0F9F9F9",
 10112 => x"C0C0C0F9C0F9F9A4",
 10113 => x"C0C0C0F9C0F9F9B0",
 10114 => x"C0C0C0F9C0F9F999",
 10115 => x"C0C0C0F9C0F9F992",
 10116 => x"C0C0C0F9C0F9F982",
 10117 => x"C0C0C0F9C0F9F9F8",
 10118 => x"C0C0C0F9C0F9F980",
 10119 => x"C0C0C0F9C0F9F990",
 10120 => x"C0C0C0F9C0F9A4C0",
 10121 => x"C0C0C0F9C0F9A4F9",
 10122 => x"C0C0C0F9C0F9A4A4",
 10123 => x"C0C0C0F9C0F9A4B0",
 10124 => x"C0C0C0F9C0F9A499",
 10125 => x"C0C0C0F9C0F9A492",
 10126 => x"C0C0C0F9C0F9A482",
 10127 => x"C0C0C0F9C0F9A4F8",
 10128 => x"C0C0C0F9C0F9A480",
 10129 => x"C0C0C0F9C0F9A490",
 10130 => x"C0C0C0F9C0F9B0C0",
 10131 => x"C0C0C0F9C0F9B0F9",
 10132 => x"C0C0C0F9C0F9B0A4",
 10133 => x"C0C0C0F9C0F9B0B0",
 10134 => x"C0C0C0F9C0F9B099",
 10135 => x"C0C0C0F9C0F9B092",
 10136 => x"C0C0C0F9C0F9B082",
 10137 => x"C0C0C0F9C0F9B0F8",
 10138 => x"C0C0C0F9C0F9B080",
 10139 => x"C0C0C0F9C0F9B090",
 10140 => x"C0C0C0F9C0F999C0",
 10141 => x"C0C0C0F9C0F999F9",
 10142 => x"C0C0C0F9C0F999A4",
 10143 => x"C0C0C0F9C0F999B0",
 10144 => x"C0C0C0F9C0F99999",
 10145 => x"C0C0C0F9C0F99992",
 10146 => x"C0C0C0F9C0F99982",
 10147 => x"C0C0C0F9C0F999F8",
 10148 => x"C0C0C0F9C0F99980",
 10149 => x"C0C0C0F9C0F99990",
 10150 => x"C0C0C0F9C0F992C0",
 10151 => x"C0C0C0F9C0F992F9",
 10152 => x"C0C0C0F9C0F992A4",
 10153 => x"C0C0C0F9C0F992B0",
 10154 => x"C0C0C0F9C0F99299",
 10155 => x"C0C0C0F9C0F99292",
 10156 => x"C0C0C0F9C0F99282",
 10157 => x"C0C0C0F9C0F992F8",
 10158 => x"C0C0C0F9C0F99280",
 10159 => x"C0C0C0F9C0F99290",
 10160 => x"C0C0C0F9C0F982C0",
 10161 => x"C0C0C0F9C0F982F9",
 10162 => x"C0C0C0F9C0F982A4",
 10163 => x"C0C0C0F9C0F982B0",
 10164 => x"C0C0C0F9C0F98299",
 10165 => x"C0C0C0F9C0F98292",
 10166 => x"C0C0C0F9C0F98282",
 10167 => x"C0C0C0F9C0F982F8",
 10168 => x"C0C0C0F9C0F98280",
 10169 => x"C0C0C0F9C0F98290",
 10170 => x"C0C0C0F9C0F9F8C0",
 10171 => x"C0C0C0F9C0F9F8F9",
 10172 => x"C0C0C0F9C0F9F8A4",
 10173 => x"C0C0C0F9C0F9F8B0",
 10174 => x"C0C0C0F9C0F9F899",
 10175 => x"C0C0C0F9C0F9F892",
 10176 => x"C0C0C0F9C0F9F882",
 10177 => x"C0C0C0F9C0F9F8F8",
 10178 => x"C0C0C0F9C0F9F880",
 10179 => x"C0C0C0F9C0F9F890",
 10180 => x"C0C0C0F9C0F980C0",
 10181 => x"C0C0C0F9C0F980F9",
 10182 => x"C0C0C0F9C0F980A4",
 10183 => x"C0C0C0F9C0F980B0",
 10184 => x"C0C0C0F9C0F98099",
 10185 => x"C0C0C0F9C0F98092",
 10186 => x"C0C0C0F9C0F98082",
 10187 => x"C0C0C0F9C0F980F8",
 10188 => x"C0C0C0F9C0F98080",
 10189 => x"C0C0C0F9C0F98090",
 10190 => x"C0C0C0F9C0F990C0",
 10191 => x"C0C0C0F9C0F990F9",
 10192 => x"C0C0C0F9C0F990A4",
 10193 => x"C0C0C0F9C0F990B0",
 10194 => x"C0C0C0F9C0F99099",
 10195 => x"C0C0C0F9C0F99092",
 10196 => x"C0C0C0F9C0F99082",
 10197 => x"C0C0C0F9C0F990F8",
 10198 => x"C0C0C0F9C0F99080",
 10199 => x"C0C0C0F9C0F99090",
 10200 => x"C0C0C0F9C0A4C0C0",
 10201 => x"C0C0C0F9C0A4C0F9",
 10202 => x"C0C0C0F9C0A4C0A4",
 10203 => x"C0C0C0F9C0A4C0B0",
 10204 => x"C0C0C0F9C0A4C099",
 10205 => x"C0C0C0F9C0A4C092",
 10206 => x"C0C0C0F9C0A4C082",
 10207 => x"C0C0C0F9C0A4C0F8",
 10208 => x"C0C0C0F9C0A4C080",
 10209 => x"C0C0C0F9C0A4C090",
 10210 => x"C0C0C0F9C0A4F9C0",
 10211 => x"C0C0C0F9C0A4F9F9",
 10212 => x"C0C0C0F9C0A4F9A4",
 10213 => x"C0C0C0F9C0A4F9B0",
 10214 => x"C0C0C0F9C0A4F999",
 10215 => x"C0C0C0F9C0A4F992",
 10216 => x"C0C0C0F9C0A4F982",
 10217 => x"C0C0C0F9C0A4F9F8",
 10218 => x"C0C0C0F9C0A4F980",
 10219 => x"C0C0C0F9C0A4F990",
 10220 => x"C0C0C0F9C0A4A4C0",
 10221 => x"C0C0C0F9C0A4A4F9",
 10222 => x"C0C0C0F9C0A4A4A4",
 10223 => x"C0C0C0F9C0A4A4B0",
 10224 => x"C0C0C0F9C0A4A499",
 10225 => x"C0C0C0F9C0A4A492",
 10226 => x"C0C0C0F9C0A4A482",
 10227 => x"C0C0C0F9C0A4A4F8",
 10228 => x"C0C0C0F9C0A4A480",
 10229 => x"C0C0C0F9C0A4A490",
 10230 => x"C0C0C0F9C0A4B0C0",
 10231 => x"C0C0C0F9C0A4B0F9",
 10232 => x"C0C0C0F9C0A4B0A4",
 10233 => x"C0C0C0F9C0A4B0B0",
 10234 => x"C0C0C0F9C0A4B099",
 10235 => x"C0C0C0F9C0A4B092",
 10236 => x"C0C0C0F9C0A4B082",
 10237 => x"C0C0C0F9C0A4B0F8",
 10238 => x"C0C0C0F9C0A4B080",
 10239 => x"C0C0C0F9C0A4B090",
 10240 => x"C0C0C0F9C0A499C0",
 10241 => x"C0C0C0F9C0A499F9",
 10242 => x"C0C0C0F9C0A499A4",
 10243 => x"C0C0C0F9C0A499B0",
 10244 => x"C0C0C0F9C0A49999",
 10245 => x"C0C0C0F9C0A49992",
 10246 => x"C0C0C0F9C0A49982",
 10247 => x"C0C0C0F9C0A499F8",
 10248 => x"C0C0C0F9C0A49980",
 10249 => x"C0C0C0F9C0A49990",
 10250 => x"C0C0C0F9C0A492C0",
 10251 => x"C0C0C0F9C0A492F9",
 10252 => x"C0C0C0F9C0A492A4",
 10253 => x"C0C0C0F9C0A492B0",
 10254 => x"C0C0C0F9C0A49299",
 10255 => x"C0C0C0F9C0A49292",
 10256 => x"C0C0C0F9C0A49282",
 10257 => x"C0C0C0F9C0A492F8",
 10258 => x"C0C0C0F9C0A49280",
 10259 => x"C0C0C0F9C0A49290",
 10260 => x"C0C0C0F9C0A482C0",
 10261 => x"C0C0C0F9C0A482F9",
 10262 => x"C0C0C0F9C0A482A4",
 10263 => x"C0C0C0F9C0A482B0",
 10264 => x"C0C0C0F9C0A48299",
 10265 => x"C0C0C0F9C0A48292",
 10266 => x"C0C0C0F9C0A48282",
 10267 => x"C0C0C0F9C0A482F8",
 10268 => x"C0C0C0F9C0A48280",
 10269 => x"C0C0C0F9C0A48290",
 10270 => x"C0C0C0F9C0A4F8C0",
 10271 => x"C0C0C0F9C0A4F8F9",
 10272 => x"C0C0C0F9C0A4F8A4",
 10273 => x"C0C0C0F9C0A4F8B0",
 10274 => x"C0C0C0F9C0A4F899",
 10275 => x"C0C0C0F9C0A4F892",
 10276 => x"C0C0C0F9C0A4F882",
 10277 => x"C0C0C0F9C0A4F8F8",
 10278 => x"C0C0C0F9C0A4F880",
 10279 => x"C0C0C0F9C0A4F890",
 10280 => x"C0C0C0F9C0A480C0",
 10281 => x"C0C0C0F9C0A480F9",
 10282 => x"C0C0C0F9C0A480A4",
 10283 => x"C0C0C0F9C0A480B0",
 10284 => x"C0C0C0F9C0A48099",
 10285 => x"C0C0C0F9C0A48092",
 10286 => x"C0C0C0F9C0A48082",
 10287 => x"C0C0C0F9C0A480F8",
 10288 => x"C0C0C0F9C0A48080",
 10289 => x"C0C0C0F9C0A48090",
 10290 => x"C0C0C0F9C0A490C0",
 10291 => x"C0C0C0F9C0A490F9",
 10292 => x"C0C0C0F9C0A490A4",
 10293 => x"C0C0C0F9C0A490B0",
 10294 => x"C0C0C0F9C0A49099",
 10295 => x"C0C0C0F9C0A49092",
 10296 => x"C0C0C0F9C0A49082",
 10297 => x"C0C0C0F9C0A490F8",
 10298 => x"C0C0C0F9C0A49080",
 10299 => x"C0C0C0F9C0A49090",
 10300 => x"C0C0C0F9C0B0C0C0",
 10301 => x"C0C0C0F9C0B0C0F9",
 10302 => x"C0C0C0F9C0B0C0A4",
 10303 => x"C0C0C0F9C0B0C0B0",
 10304 => x"C0C0C0F9C0B0C099",
 10305 => x"C0C0C0F9C0B0C092",
 10306 => x"C0C0C0F9C0B0C082",
 10307 => x"C0C0C0F9C0B0C0F8",
 10308 => x"C0C0C0F9C0B0C080",
 10309 => x"C0C0C0F9C0B0C090",
 10310 => x"C0C0C0F9C0B0F9C0",
 10311 => x"C0C0C0F9C0B0F9F9",
 10312 => x"C0C0C0F9C0B0F9A4",
 10313 => x"C0C0C0F9C0B0F9B0",
 10314 => x"C0C0C0F9C0B0F999",
 10315 => x"C0C0C0F9C0B0F992",
 10316 => x"C0C0C0F9C0B0F982",
 10317 => x"C0C0C0F9C0B0F9F8",
 10318 => x"C0C0C0F9C0B0F980",
 10319 => x"C0C0C0F9C0B0F990",
 10320 => x"C0C0C0F9C0B0A4C0",
 10321 => x"C0C0C0F9C0B0A4F9",
 10322 => x"C0C0C0F9C0B0A4A4",
 10323 => x"C0C0C0F9C0B0A4B0",
 10324 => x"C0C0C0F9C0B0A499",
 10325 => x"C0C0C0F9C0B0A492",
 10326 => x"C0C0C0F9C0B0A482",
 10327 => x"C0C0C0F9C0B0A4F8",
 10328 => x"C0C0C0F9C0B0A480",
 10329 => x"C0C0C0F9C0B0A490",
 10330 => x"C0C0C0F9C0B0B0C0",
 10331 => x"C0C0C0F9C0B0B0F9",
 10332 => x"C0C0C0F9C0B0B0A4",
 10333 => x"C0C0C0F9C0B0B0B0",
 10334 => x"C0C0C0F9C0B0B099",
 10335 => x"C0C0C0F9C0B0B092",
 10336 => x"C0C0C0F9C0B0B082",
 10337 => x"C0C0C0F9C0B0B0F8",
 10338 => x"C0C0C0F9C0B0B080",
 10339 => x"C0C0C0F9C0B0B090",
 10340 => x"C0C0C0F9C0B099C0",
 10341 => x"C0C0C0F9C0B099F9",
 10342 => x"C0C0C0F9C0B099A4",
 10343 => x"C0C0C0F9C0B099B0",
 10344 => x"C0C0C0F9C0B09999",
 10345 => x"C0C0C0F9C0B09992",
 10346 => x"C0C0C0F9C0B09982",
 10347 => x"C0C0C0F9C0B099F8",
 10348 => x"C0C0C0F9C0B09980",
 10349 => x"C0C0C0F9C0B09990",
 10350 => x"C0C0C0F9C0B092C0",
 10351 => x"C0C0C0F9C0B092F9",
 10352 => x"C0C0C0F9C0B092A4",
 10353 => x"C0C0C0F9C0B092B0",
 10354 => x"C0C0C0F9C0B09299",
 10355 => x"C0C0C0F9C0B09292",
 10356 => x"C0C0C0F9C0B09282",
 10357 => x"C0C0C0F9C0B092F8",
 10358 => x"C0C0C0F9C0B09280",
 10359 => x"C0C0C0F9C0B09290",
 10360 => x"C0C0C0F9C0B082C0",
 10361 => x"C0C0C0F9C0B082F9",
 10362 => x"C0C0C0F9C0B082A4",
 10363 => x"C0C0C0F9C0B082B0",
 10364 => x"C0C0C0F9C0B08299",
 10365 => x"C0C0C0F9C0B08292",
 10366 => x"C0C0C0F9C0B08282",
 10367 => x"C0C0C0F9C0B082F8",
 10368 => x"C0C0C0F9C0B08280",
 10369 => x"C0C0C0F9C0B08290",
 10370 => x"C0C0C0F9C0B0F8C0",
 10371 => x"C0C0C0F9C0B0F8F9",
 10372 => x"C0C0C0F9C0B0F8A4",
 10373 => x"C0C0C0F9C0B0F8B0",
 10374 => x"C0C0C0F9C0B0F899",
 10375 => x"C0C0C0F9C0B0F892",
 10376 => x"C0C0C0F9C0B0F882",
 10377 => x"C0C0C0F9C0B0F8F8",
 10378 => x"C0C0C0F9C0B0F880",
 10379 => x"C0C0C0F9C0B0F890",
 10380 => x"C0C0C0F9C0B080C0",
 10381 => x"C0C0C0F9C0B080F9",
 10382 => x"C0C0C0F9C0B080A4",
 10383 => x"C0C0C0F9C0B080B0",
 10384 => x"C0C0C0F9C0B08099",
 10385 => x"C0C0C0F9C0B08092",
 10386 => x"C0C0C0F9C0B08082",
 10387 => x"C0C0C0F9C0B080F8",
 10388 => x"C0C0C0F9C0B08080",
 10389 => x"C0C0C0F9C0B08090",
 10390 => x"C0C0C0F9C0B090C0",
 10391 => x"C0C0C0F9C0B090F9",
 10392 => x"C0C0C0F9C0B090A4",
 10393 => x"C0C0C0F9C0B090B0",
 10394 => x"C0C0C0F9C0B09099",
 10395 => x"C0C0C0F9C0B09092",
 10396 => x"C0C0C0F9C0B09082",
 10397 => x"C0C0C0F9C0B090F8",
 10398 => x"C0C0C0F9C0B09080",
 10399 => x"C0C0C0F9C0B09090",
 10400 => x"C0C0C0F9C099C0C0",
 10401 => x"C0C0C0F9C099C0F9",
 10402 => x"C0C0C0F9C099C0A4",
 10403 => x"C0C0C0F9C099C0B0",
 10404 => x"C0C0C0F9C099C099",
 10405 => x"C0C0C0F9C099C092",
 10406 => x"C0C0C0F9C099C082",
 10407 => x"C0C0C0F9C099C0F8",
 10408 => x"C0C0C0F9C099C080",
 10409 => x"C0C0C0F9C099C090",
 10410 => x"C0C0C0F9C099F9C0",
 10411 => x"C0C0C0F9C099F9F9",
 10412 => x"C0C0C0F9C099F9A4",
 10413 => x"C0C0C0F9C099F9B0",
 10414 => x"C0C0C0F9C099F999",
 10415 => x"C0C0C0F9C099F992",
 10416 => x"C0C0C0F9C099F982",
 10417 => x"C0C0C0F9C099F9F8",
 10418 => x"C0C0C0F9C099F980",
 10419 => x"C0C0C0F9C099F990",
 10420 => x"C0C0C0F9C099A4C0",
 10421 => x"C0C0C0F9C099A4F9",
 10422 => x"C0C0C0F9C099A4A4",
 10423 => x"C0C0C0F9C099A4B0",
 10424 => x"C0C0C0F9C099A499",
 10425 => x"C0C0C0F9C099A492",
 10426 => x"C0C0C0F9C099A482",
 10427 => x"C0C0C0F9C099A4F8",
 10428 => x"C0C0C0F9C099A480",
 10429 => x"C0C0C0F9C099A490",
 10430 => x"C0C0C0F9C099B0C0",
 10431 => x"C0C0C0F9C099B0F9",
 10432 => x"C0C0C0F9C099B0A4",
 10433 => x"C0C0C0F9C099B0B0",
 10434 => x"C0C0C0F9C099B099",
 10435 => x"C0C0C0F9C099B092",
 10436 => x"C0C0C0F9C099B082",
 10437 => x"C0C0C0F9C099B0F8",
 10438 => x"C0C0C0F9C099B080",
 10439 => x"C0C0C0F9C099B090",
 10440 => x"C0C0C0F9C09999C0",
 10441 => x"C0C0C0F9C09999F9",
 10442 => x"C0C0C0F9C09999A4",
 10443 => x"C0C0C0F9C09999B0",
 10444 => x"C0C0C0F9C0999999",
 10445 => x"C0C0C0F9C0999992",
 10446 => x"C0C0C0F9C0999982",
 10447 => x"C0C0C0F9C09999F8",
 10448 => x"C0C0C0F9C0999980",
 10449 => x"C0C0C0F9C0999990",
 10450 => x"C0C0C0F9C09992C0",
 10451 => x"C0C0C0F9C09992F9",
 10452 => x"C0C0C0F9C09992A4",
 10453 => x"C0C0C0F9C09992B0",
 10454 => x"C0C0C0F9C0999299",
 10455 => x"C0C0C0F9C0999292",
 10456 => x"C0C0C0F9C0999282",
 10457 => x"C0C0C0F9C09992F8",
 10458 => x"C0C0C0F9C0999280",
 10459 => x"C0C0C0F9C0999290",
 10460 => x"C0C0C0F9C09982C0",
 10461 => x"C0C0C0F9C09982F9",
 10462 => x"C0C0C0F9C09982A4",
 10463 => x"C0C0C0F9C09982B0",
 10464 => x"C0C0C0F9C0998299",
 10465 => x"C0C0C0F9C0998292",
 10466 => x"C0C0C0F9C0998282",
 10467 => x"C0C0C0F9C09982F8",
 10468 => x"C0C0C0F9C0998280",
 10469 => x"C0C0C0F9C0998290",
 10470 => x"C0C0C0F9C099F8C0",
 10471 => x"C0C0C0F9C099F8F9",
 10472 => x"C0C0C0F9C099F8A4",
 10473 => x"C0C0C0F9C099F8B0",
 10474 => x"C0C0C0F9C099F899",
 10475 => x"C0C0C0F9C099F892",
 10476 => x"C0C0C0F9C099F882",
 10477 => x"C0C0C0F9C099F8F8",
 10478 => x"C0C0C0F9C099F880",
 10479 => x"C0C0C0F9C099F890",
 10480 => x"C0C0C0F9C09980C0",
 10481 => x"C0C0C0F9C09980F9",
 10482 => x"C0C0C0F9C09980A4",
 10483 => x"C0C0C0F9C09980B0",
 10484 => x"C0C0C0F9C0998099",
 10485 => x"C0C0C0F9C0998092",
 10486 => x"C0C0C0F9C0998082",
 10487 => x"C0C0C0F9C09980F8",
 10488 => x"C0C0C0F9C0998080",
 10489 => x"C0C0C0F9C0998090",
 10490 => x"C0C0C0F9C09990C0",
 10491 => x"C0C0C0F9C09990F9",
 10492 => x"C0C0C0F9C09990A4",
 10493 => x"C0C0C0F9C09990B0",
 10494 => x"C0C0C0F9C0999099",
 10495 => x"C0C0C0F9C0999092",
 10496 => x"C0C0C0F9C0999082",
 10497 => x"C0C0C0F9C09990F8",
 10498 => x"C0C0C0F9C0999080",
 10499 => x"C0C0C0F9C0999090",
 10500 => x"C0C0C0F9C092C0C0",
 10501 => x"C0C0C0F9C092C0F9",
 10502 => x"C0C0C0F9C092C0A4",
 10503 => x"C0C0C0F9C092C0B0",
 10504 => x"C0C0C0F9C092C099",
 10505 => x"C0C0C0F9C092C092",
 10506 => x"C0C0C0F9C092C082",
 10507 => x"C0C0C0F9C092C0F8",
 10508 => x"C0C0C0F9C092C080",
 10509 => x"C0C0C0F9C092C090",
 10510 => x"C0C0C0F9C092F9C0",
 10511 => x"C0C0C0F9C092F9F9",
 10512 => x"C0C0C0F9C092F9A4",
 10513 => x"C0C0C0F9C092F9B0",
 10514 => x"C0C0C0F9C092F999",
 10515 => x"C0C0C0F9C092F992",
 10516 => x"C0C0C0F9C092F982",
 10517 => x"C0C0C0F9C092F9F8",
 10518 => x"C0C0C0F9C092F980",
 10519 => x"C0C0C0F9C092F990",
 10520 => x"C0C0C0F9C092A4C0",
 10521 => x"C0C0C0F9C092A4F9",
 10522 => x"C0C0C0F9C092A4A4",
 10523 => x"C0C0C0F9C092A4B0",
 10524 => x"C0C0C0F9C092A499",
 10525 => x"C0C0C0F9C092A492",
 10526 => x"C0C0C0F9C092A482",
 10527 => x"C0C0C0F9C092A4F8",
 10528 => x"C0C0C0F9C092A480",
 10529 => x"C0C0C0F9C092A490",
 10530 => x"C0C0C0F9C092B0C0",
 10531 => x"C0C0C0F9C092B0F9",
 10532 => x"C0C0C0F9C092B0A4",
 10533 => x"C0C0C0F9C092B0B0",
 10534 => x"C0C0C0F9C092B099",
 10535 => x"C0C0C0F9C092B092",
 10536 => x"C0C0C0F9C092B082",
 10537 => x"C0C0C0F9C092B0F8",
 10538 => x"C0C0C0F9C092B080",
 10539 => x"C0C0C0F9C092B090",
 10540 => x"C0C0C0F9C09299C0",
 10541 => x"C0C0C0F9C09299F9",
 10542 => x"C0C0C0F9C09299A4",
 10543 => x"C0C0C0F9C09299B0",
 10544 => x"C0C0C0F9C0929999",
 10545 => x"C0C0C0F9C0929992",
 10546 => x"C0C0C0F9C0929982",
 10547 => x"C0C0C0F9C09299F8",
 10548 => x"C0C0C0F9C0929980",
 10549 => x"C0C0C0F9C0929990",
 10550 => x"C0C0C0F9C09292C0",
 10551 => x"C0C0C0F9C09292F9",
 10552 => x"C0C0C0F9C09292A4",
 10553 => x"C0C0C0F9C09292B0",
 10554 => x"C0C0C0F9C0929299",
 10555 => x"C0C0C0F9C0929292",
 10556 => x"C0C0C0F9C0929282",
 10557 => x"C0C0C0F9C09292F8",
 10558 => x"C0C0C0F9C0929280",
 10559 => x"C0C0C0F9C0929290",
 10560 => x"C0C0C0F9C09282C0",
 10561 => x"C0C0C0F9C09282F9",
 10562 => x"C0C0C0F9C09282A4",
 10563 => x"C0C0C0F9C09282B0",
 10564 => x"C0C0C0F9C0928299",
 10565 => x"C0C0C0F9C0928292",
 10566 => x"C0C0C0F9C0928282",
 10567 => x"C0C0C0F9C09282F8",
 10568 => x"C0C0C0F9C0928280",
 10569 => x"C0C0C0F9C0928290",
 10570 => x"C0C0C0F9C092F8C0",
 10571 => x"C0C0C0F9C092F8F9",
 10572 => x"C0C0C0F9C092F8A4",
 10573 => x"C0C0C0F9C092F8B0",
 10574 => x"C0C0C0F9C092F899",
 10575 => x"C0C0C0F9C092F892",
 10576 => x"C0C0C0F9C092F882",
 10577 => x"C0C0C0F9C092F8F8",
 10578 => x"C0C0C0F9C092F880",
 10579 => x"C0C0C0F9C092F890",
 10580 => x"C0C0C0F9C09280C0",
 10581 => x"C0C0C0F9C09280F9",
 10582 => x"C0C0C0F9C09280A4",
 10583 => x"C0C0C0F9C09280B0",
 10584 => x"C0C0C0F9C0928099",
 10585 => x"C0C0C0F9C0928092",
 10586 => x"C0C0C0F9C0928082",
 10587 => x"C0C0C0F9C09280F8",
 10588 => x"C0C0C0F9C0928080",
 10589 => x"C0C0C0F9C0928090",
 10590 => x"C0C0C0F9C09290C0",
 10591 => x"C0C0C0F9C09290F9",
 10592 => x"C0C0C0F9C09290A4",
 10593 => x"C0C0C0F9C09290B0",
 10594 => x"C0C0C0F9C0929099",
 10595 => x"C0C0C0F9C0929092",
 10596 => x"C0C0C0F9C0929082",
 10597 => x"C0C0C0F9C09290F8",
 10598 => x"C0C0C0F9C0929080",
 10599 => x"C0C0C0F9C0929090",
 10600 => x"C0C0C0F9C082C0C0",
 10601 => x"C0C0C0F9C082C0F9",
 10602 => x"C0C0C0F9C082C0A4",
 10603 => x"C0C0C0F9C082C0B0",
 10604 => x"C0C0C0F9C082C099",
 10605 => x"C0C0C0F9C082C092",
 10606 => x"C0C0C0F9C082C082",
 10607 => x"C0C0C0F9C082C0F8",
 10608 => x"C0C0C0F9C082C080",
 10609 => x"C0C0C0F9C082C090",
 10610 => x"C0C0C0F9C082F9C0",
 10611 => x"C0C0C0F9C082F9F9",
 10612 => x"C0C0C0F9C082F9A4",
 10613 => x"C0C0C0F9C082F9B0",
 10614 => x"C0C0C0F9C082F999",
 10615 => x"C0C0C0F9C082F992",
 10616 => x"C0C0C0F9C082F982",
 10617 => x"C0C0C0F9C082F9F8",
 10618 => x"C0C0C0F9C082F980",
 10619 => x"C0C0C0F9C082F990",
 10620 => x"C0C0C0F9C082A4C0",
 10621 => x"C0C0C0F9C082A4F9",
 10622 => x"C0C0C0F9C082A4A4",
 10623 => x"C0C0C0F9C082A4B0",
 10624 => x"C0C0C0F9C082A499",
 10625 => x"C0C0C0F9C082A492",
 10626 => x"C0C0C0F9C082A482",
 10627 => x"C0C0C0F9C082A4F8",
 10628 => x"C0C0C0F9C082A480",
 10629 => x"C0C0C0F9C082A490",
 10630 => x"C0C0C0F9C082B0C0",
 10631 => x"C0C0C0F9C082B0F9",
 10632 => x"C0C0C0F9C082B0A4",
 10633 => x"C0C0C0F9C082B0B0",
 10634 => x"C0C0C0F9C082B099",
 10635 => x"C0C0C0F9C082B092",
 10636 => x"C0C0C0F9C082B082",
 10637 => x"C0C0C0F9C082B0F8",
 10638 => x"C0C0C0F9C082B080",
 10639 => x"C0C0C0F9C082B090",
 10640 => x"C0C0C0F9C08299C0",
 10641 => x"C0C0C0F9C08299F9",
 10642 => x"C0C0C0F9C08299A4",
 10643 => x"C0C0C0F9C08299B0",
 10644 => x"C0C0C0F9C0829999",
 10645 => x"C0C0C0F9C0829992",
 10646 => x"C0C0C0F9C0829982",
 10647 => x"C0C0C0F9C08299F8",
 10648 => x"C0C0C0F9C0829980",
 10649 => x"C0C0C0F9C0829990",
 10650 => x"C0C0C0F9C08292C0",
 10651 => x"C0C0C0F9C08292F9",
 10652 => x"C0C0C0F9C08292A4",
 10653 => x"C0C0C0F9C08292B0",
 10654 => x"C0C0C0F9C0829299",
 10655 => x"C0C0C0F9C0829292",
 10656 => x"C0C0C0F9C0829282",
 10657 => x"C0C0C0F9C08292F8",
 10658 => x"C0C0C0F9C0829280",
 10659 => x"C0C0C0F9C0829290",
 10660 => x"C0C0C0F9C08282C0",
 10661 => x"C0C0C0F9C08282F9",
 10662 => x"C0C0C0F9C08282A4",
 10663 => x"C0C0C0F9C08282B0",
 10664 => x"C0C0C0F9C0828299",
 10665 => x"C0C0C0F9C0828292",
 10666 => x"C0C0C0F9C0828282",
 10667 => x"C0C0C0F9C08282F8",
 10668 => x"C0C0C0F9C0828280",
 10669 => x"C0C0C0F9C0828290",
 10670 => x"C0C0C0F9C082F8C0",
 10671 => x"C0C0C0F9C082F8F9",
 10672 => x"C0C0C0F9C082F8A4",
 10673 => x"C0C0C0F9C082F8B0",
 10674 => x"C0C0C0F9C082F899",
 10675 => x"C0C0C0F9C082F892",
 10676 => x"C0C0C0F9C082F882",
 10677 => x"C0C0C0F9C082F8F8",
 10678 => x"C0C0C0F9C082F880",
 10679 => x"C0C0C0F9C082F890",
 10680 => x"C0C0C0F9C08280C0",
 10681 => x"C0C0C0F9C08280F9",
 10682 => x"C0C0C0F9C08280A4",
 10683 => x"C0C0C0F9C08280B0",
 10684 => x"C0C0C0F9C0828099",
 10685 => x"C0C0C0F9C0828092",
 10686 => x"C0C0C0F9C0828082",
 10687 => x"C0C0C0F9C08280F8",
 10688 => x"C0C0C0F9C0828080",
 10689 => x"C0C0C0F9C0828090",
 10690 => x"C0C0C0F9C08290C0",
 10691 => x"C0C0C0F9C08290F9",
 10692 => x"C0C0C0F9C08290A4",
 10693 => x"C0C0C0F9C08290B0",
 10694 => x"C0C0C0F9C0829099",
 10695 => x"C0C0C0F9C0829092",
 10696 => x"C0C0C0F9C0829082",
 10697 => x"C0C0C0F9C08290F8",
 10698 => x"C0C0C0F9C0829080",
 10699 => x"C0C0C0F9C0829090",
 10700 => x"C0C0C0F9C0F8C0C0",
 10701 => x"C0C0C0F9C0F8C0F9",
 10702 => x"C0C0C0F9C0F8C0A4",
 10703 => x"C0C0C0F9C0F8C0B0",
 10704 => x"C0C0C0F9C0F8C099",
 10705 => x"C0C0C0F9C0F8C092",
 10706 => x"C0C0C0F9C0F8C082",
 10707 => x"C0C0C0F9C0F8C0F8",
 10708 => x"C0C0C0F9C0F8C080",
 10709 => x"C0C0C0F9C0F8C090",
 10710 => x"C0C0C0F9C0F8F9C0",
 10711 => x"C0C0C0F9C0F8F9F9",
 10712 => x"C0C0C0F9C0F8F9A4",
 10713 => x"C0C0C0F9C0F8F9B0",
 10714 => x"C0C0C0F9C0F8F999",
 10715 => x"C0C0C0F9C0F8F992",
 10716 => x"C0C0C0F9C0F8F982",
 10717 => x"C0C0C0F9C0F8F9F8",
 10718 => x"C0C0C0F9C0F8F980",
 10719 => x"C0C0C0F9C0F8F990",
 10720 => x"C0C0C0F9C0F8A4C0",
 10721 => x"C0C0C0F9C0F8A4F9",
 10722 => x"C0C0C0F9C0F8A4A4",
 10723 => x"C0C0C0F9C0F8A4B0",
 10724 => x"C0C0C0F9C0F8A499",
 10725 => x"C0C0C0F9C0F8A492",
 10726 => x"C0C0C0F9C0F8A482",
 10727 => x"C0C0C0F9C0F8A4F8",
 10728 => x"C0C0C0F9C0F8A480",
 10729 => x"C0C0C0F9C0F8A490",
 10730 => x"C0C0C0F9C0F8B0C0",
 10731 => x"C0C0C0F9C0F8B0F9",
 10732 => x"C0C0C0F9C0F8B0A4",
 10733 => x"C0C0C0F9C0F8B0B0",
 10734 => x"C0C0C0F9C0F8B099",
 10735 => x"C0C0C0F9C0F8B092",
 10736 => x"C0C0C0F9C0F8B082",
 10737 => x"C0C0C0F9C0F8B0F8",
 10738 => x"C0C0C0F9C0F8B080",
 10739 => x"C0C0C0F9C0F8B090",
 10740 => x"C0C0C0F9C0F899C0",
 10741 => x"C0C0C0F9C0F899F9",
 10742 => x"C0C0C0F9C0F899A4",
 10743 => x"C0C0C0F9C0F899B0",
 10744 => x"C0C0C0F9C0F89999",
 10745 => x"C0C0C0F9C0F89992",
 10746 => x"C0C0C0F9C0F89982",
 10747 => x"C0C0C0F9C0F899F8",
 10748 => x"C0C0C0F9C0F89980",
 10749 => x"C0C0C0F9C0F89990",
 10750 => x"C0C0C0F9C0F892C0",
 10751 => x"C0C0C0F9C0F892F9",
 10752 => x"C0C0C0F9C0F892A4",
 10753 => x"C0C0C0F9C0F892B0",
 10754 => x"C0C0C0F9C0F89299",
 10755 => x"C0C0C0F9C0F89292",
 10756 => x"C0C0C0F9C0F89282",
 10757 => x"C0C0C0F9C0F892F8",
 10758 => x"C0C0C0F9C0F89280",
 10759 => x"C0C0C0F9C0F89290",
 10760 => x"C0C0C0F9C0F882C0",
 10761 => x"C0C0C0F9C0F882F9",
 10762 => x"C0C0C0F9C0F882A4",
 10763 => x"C0C0C0F9C0F882B0",
 10764 => x"C0C0C0F9C0F88299",
 10765 => x"C0C0C0F9C0F88292",
 10766 => x"C0C0C0F9C0F88282",
 10767 => x"C0C0C0F9C0F882F8",
 10768 => x"C0C0C0F9C0F88280",
 10769 => x"C0C0C0F9C0F88290",
 10770 => x"C0C0C0F9C0F8F8C0",
 10771 => x"C0C0C0F9C0F8F8F9",
 10772 => x"C0C0C0F9C0F8F8A4",
 10773 => x"C0C0C0F9C0F8F8B0",
 10774 => x"C0C0C0F9C0F8F899",
 10775 => x"C0C0C0F9C0F8F892",
 10776 => x"C0C0C0F9C0F8F882",
 10777 => x"C0C0C0F9C0F8F8F8",
 10778 => x"C0C0C0F9C0F8F880",
 10779 => x"C0C0C0F9C0F8F890",
 10780 => x"C0C0C0F9C0F880C0",
 10781 => x"C0C0C0F9C0F880F9",
 10782 => x"C0C0C0F9C0F880A4",
 10783 => x"C0C0C0F9C0F880B0",
 10784 => x"C0C0C0F9C0F88099",
 10785 => x"C0C0C0F9C0F88092",
 10786 => x"C0C0C0F9C0F88082",
 10787 => x"C0C0C0F9C0F880F8",
 10788 => x"C0C0C0F9C0F88080",
 10789 => x"C0C0C0F9C0F88090",
 10790 => x"C0C0C0F9C0F890C0",
 10791 => x"C0C0C0F9C0F890F9",
 10792 => x"C0C0C0F9C0F890A4",
 10793 => x"C0C0C0F9C0F890B0",
 10794 => x"C0C0C0F9C0F89099",
 10795 => x"C0C0C0F9C0F89092",
 10796 => x"C0C0C0F9C0F89082",
 10797 => x"C0C0C0F9C0F890F8",
 10798 => x"C0C0C0F9C0F89080",
 10799 => x"C0C0C0F9C0F89090",
 10800 => x"C0C0C0F9C080C0C0",
 10801 => x"C0C0C0F9C080C0F9",
 10802 => x"C0C0C0F9C080C0A4",
 10803 => x"C0C0C0F9C080C0B0",
 10804 => x"C0C0C0F9C080C099",
 10805 => x"C0C0C0F9C080C092",
 10806 => x"C0C0C0F9C080C082",
 10807 => x"C0C0C0F9C080C0F8",
 10808 => x"C0C0C0F9C080C080",
 10809 => x"C0C0C0F9C080C090",
 10810 => x"C0C0C0F9C080F9C0",
 10811 => x"C0C0C0F9C080F9F9",
 10812 => x"C0C0C0F9C080F9A4",
 10813 => x"C0C0C0F9C080F9B0",
 10814 => x"C0C0C0F9C080F999",
 10815 => x"C0C0C0F9C080F992",
 10816 => x"C0C0C0F9C080F982",
 10817 => x"C0C0C0F9C080F9F8",
 10818 => x"C0C0C0F9C080F980",
 10819 => x"C0C0C0F9C080F990",
 10820 => x"C0C0C0F9C080A4C0",
 10821 => x"C0C0C0F9C080A4F9",
 10822 => x"C0C0C0F9C080A4A4",
 10823 => x"C0C0C0F9C080A4B0",
 10824 => x"C0C0C0F9C080A499",
 10825 => x"C0C0C0F9C080A492",
 10826 => x"C0C0C0F9C080A482",
 10827 => x"C0C0C0F9C080A4F8",
 10828 => x"C0C0C0F9C080A480",
 10829 => x"C0C0C0F9C080A490",
 10830 => x"C0C0C0F9C080B0C0",
 10831 => x"C0C0C0F9C080B0F9",
 10832 => x"C0C0C0F9C080B0A4",
 10833 => x"C0C0C0F9C080B0B0",
 10834 => x"C0C0C0F9C080B099",
 10835 => x"C0C0C0F9C080B092",
 10836 => x"C0C0C0F9C080B082",
 10837 => x"C0C0C0F9C080B0F8",
 10838 => x"C0C0C0F9C080B080",
 10839 => x"C0C0C0F9C080B090",
 10840 => x"C0C0C0F9C08099C0",
 10841 => x"C0C0C0F9C08099F9",
 10842 => x"C0C0C0F9C08099A4",
 10843 => x"C0C0C0F9C08099B0",
 10844 => x"C0C0C0F9C0809999",
 10845 => x"C0C0C0F9C0809992",
 10846 => x"C0C0C0F9C0809982",
 10847 => x"C0C0C0F9C08099F8",
 10848 => x"C0C0C0F9C0809980",
 10849 => x"C0C0C0F9C0809990",
 10850 => x"C0C0C0F9C08092C0",
 10851 => x"C0C0C0F9C08092F9",
 10852 => x"C0C0C0F9C08092A4",
 10853 => x"C0C0C0F9C08092B0",
 10854 => x"C0C0C0F9C0809299",
 10855 => x"C0C0C0F9C0809292",
 10856 => x"C0C0C0F9C0809282",
 10857 => x"C0C0C0F9C08092F8",
 10858 => x"C0C0C0F9C0809280",
 10859 => x"C0C0C0F9C0809290",
 10860 => x"C0C0C0F9C08082C0",
 10861 => x"C0C0C0F9C08082F9",
 10862 => x"C0C0C0F9C08082A4",
 10863 => x"C0C0C0F9C08082B0",
 10864 => x"C0C0C0F9C0808299",
 10865 => x"C0C0C0F9C0808292",
 10866 => x"C0C0C0F9C0808282",
 10867 => x"C0C0C0F9C08082F8",
 10868 => x"C0C0C0F9C0808280",
 10869 => x"C0C0C0F9C0808290",
 10870 => x"C0C0C0F9C080F8C0",
 10871 => x"C0C0C0F9C080F8F9",
 10872 => x"C0C0C0F9C080F8A4",
 10873 => x"C0C0C0F9C080F8B0",
 10874 => x"C0C0C0F9C080F899",
 10875 => x"C0C0C0F9C080F892",
 10876 => x"C0C0C0F9C080F882",
 10877 => x"C0C0C0F9C080F8F8",
 10878 => x"C0C0C0F9C080F880",
 10879 => x"C0C0C0F9C080F890",
 10880 => x"C0C0C0F9C08080C0",
 10881 => x"C0C0C0F9C08080F9",
 10882 => x"C0C0C0F9C08080A4",
 10883 => x"C0C0C0F9C08080B0",
 10884 => x"C0C0C0F9C0808099",
 10885 => x"C0C0C0F9C0808092",
 10886 => x"C0C0C0F9C0808082",
 10887 => x"C0C0C0F9C08080F8",
 10888 => x"C0C0C0F9C0808080",
 10889 => x"C0C0C0F9C0808090",
 10890 => x"C0C0C0F9C08090C0",
 10891 => x"C0C0C0F9C08090F9",
 10892 => x"C0C0C0F9C08090A4",
 10893 => x"C0C0C0F9C08090B0",
 10894 => x"C0C0C0F9C0809099",
 10895 => x"C0C0C0F9C0809092",
 10896 => x"C0C0C0F9C0809082",
 10897 => x"C0C0C0F9C08090F8",
 10898 => x"C0C0C0F9C0809080",
 10899 => x"C0C0C0F9C0809090",
 10900 => x"C0C0C0F9C090C0C0",
 10901 => x"C0C0C0F9C090C0F9",
 10902 => x"C0C0C0F9C090C0A4",
 10903 => x"C0C0C0F9C090C0B0",
 10904 => x"C0C0C0F9C090C099",
 10905 => x"C0C0C0F9C090C092",
 10906 => x"C0C0C0F9C090C082",
 10907 => x"C0C0C0F9C090C0F8",
 10908 => x"C0C0C0F9C090C080",
 10909 => x"C0C0C0F9C090C090",
 10910 => x"C0C0C0F9C090F9C0",
 10911 => x"C0C0C0F9C090F9F9",
 10912 => x"C0C0C0F9C090F9A4",
 10913 => x"C0C0C0F9C090F9B0",
 10914 => x"C0C0C0F9C090F999",
 10915 => x"C0C0C0F9C090F992",
 10916 => x"C0C0C0F9C090F982",
 10917 => x"C0C0C0F9C090F9F8",
 10918 => x"C0C0C0F9C090F980",
 10919 => x"C0C0C0F9C090F990",
 10920 => x"C0C0C0F9C090A4C0",
 10921 => x"C0C0C0F9C090A4F9",
 10922 => x"C0C0C0F9C090A4A4",
 10923 => x"C0C0C0F9C090A4B0",
 10924 => x"C0C0C0F9C090A499",
 10925 => x"C0C0C0F9C090A492",
 10926 => x"C0C0C0F9C090A482",
 10927 => x"C0C0C0F9C090A4F8",
 10928 => x"C0C0C0F9C090A480",
 10929 => x"C0C0C0F9C090A490",
 10930 => x"C0C0C0F9C090B0C0",
 10931 => x"C0C0C0F9C090B0F9",
 10932 => x"C0C0C0F9C090B0A4",
 10933 => x"C0C0C0F9C090B0B0",
 10934 => x"C0C0C0F9C090B099",
 10935 => x"C0C0C0F9C090B092",
 10936 => x"C0C0C0F9C090B082",
 10937 => x"C0C0C0F9C090B0F8",
 10938 => x"C0C0C0F9C090B080",
 10939 => x"C0C0C0F9C090B090",
 10940 => x"C0C0C0F9C09099C0",
 10941 => x"C0C0C0F9C09099F9",
 10942 => x"C0C0C0F9C09099A4",
 10943 => x"C0C0C0F9C09099B0",
 10944 => x"C0C0C0F9C0909999",
 10945 => x"C0C0C0F9C0909992",
 10946 => x"C0C0C0F9C0909982",
 10947 => x"C0C0C0F9C09099F8",
 10948 => x"C0C0C0F9C0909980",
 10949 => x"C0C0C0F9C0909990",
 10950 => x"C0C0C0F9C09092C0",
 10951 => x"C0C0C0F9C09092F9",
 10952 => x"C0C0C0F9C09092A4",
 10953 => x"C0C0C0F9C09092B0",
 10954 => x"C0C0C0F9C0909299",
 10955 => x"C0C0C0F9C0909292",
 10956 => x"C0C0C0F9C0909282",
 10957 => x"C0C0C0F9C09092F8",
 10958 => x"C0C0C0F9C0909280",
 10959 => x"C0C0C0F9C0909290",
 10960 => x"C0C0C0F9C09082C0",
 10961 => x"C0C0C0F9C09082F9",
 10962 => x"C0C0C0F9C09082A4",
 10963 => x"C0C0C0F9C09082B0",
 10964 => x"C0C0C0F9C0908299",
 10965 => x"C0C0C0F9C0908292",
 10966 => x"C0C0C0F9C0908282",
 10967 => x"C0C0C0F9C09082F8",
 10968 => x"C0C0C0F9C0908280",
 10969 => x"C0C0C0F9C0908290",
 10970 => x"C0C0C0F9C090F8C0",
 10971 => x"C0C0C0F9C090F8F9",
 10972 => x"C0C0C0F9C090F8A4",
 10973 => x"C0C0C0F9C090F8B0",
 10974 => x"C0C0C0F9C090F899",
 10975 => x"C0C0C0F9C090F892",
 10976 => x"C0C0C0F9C090F882",
 10977 => x"C0C0C0F9C090F8F8",
 10978 => x"C0C0C0F9C090F880",
 10979 => x"C0C0C0F9C090F890",
 10980 => x"C0C0C0F9C09080C0",
 10981 => x"C0C0C0F9C09080F9",
 10982 => x"C0C0C0F9C09080A4",
 10983 => x"C0C0C0F9C09080B0",
 10984 => x"C0C0C0F9C0908099",
 10985 => x"C0C0C0F9C0908092",
 10986 => x"C0C0C0F9C0908082",
 10987 => x"C0C0C0F9C09080F8",
 10988 => x"C0C0C0F9C0908080",
 10989 => x"C0C0C0F9C0908090",
 10990 => x"C0C0C0F9C09090C0",
 10991 => x"C0C0C0F9C09090F9",
 10992 => x"C0C0C0F9C09090A4",
 10993 => x"C0C0C0F9C09090B0",
 10994 => x"C0C0C0F9C0909099",
 10995 => x"C0C0C0F9C0909092",
 10996 => x"C0C0C0F9C0909082",
 10997 => x"C0C0C0F9C09090F8",
 10998 => x"C0C0C0F9C0909080",
 10999 => x"C0C0C0F9C0909090",
 11000 => x"C0C0C0F9F9C0C0C0",
 11001 => x"C0C0C0F9F9C0C0F9",
 11002 => x"C0C0C0F9F9C0C0A4",
 11003 => x"C0C0C0F9F9C0C0B0",
 11004 => x"C0C0C0F9F9C0C099",
 11005 => x"C0C0C0F9F9C0C092",
 11006 => x"C0C0C0F9F9C0C082",
 11007 => x"C0C0C0F9F9C0C0F8",
 11008 => x"C0C0C0F9F9C0C080",
 11009 => x"C0C0C0F9F9C0C090",
 11010 => x"C0C0C0F9F9C0F9C0",
 11011 => x"C0C0C0F9F9C0F9F9",
 11012 => x"C0C0C0F9F9C0F9A4",
 11013 => x"C0C0C0F9F9C0F9B0",
 11014 => x"C0C0C0F9F9C0F999",
 11015 => x"C0C0C0F9F9C0F992",
 11016 => x"C0C0C0F9F9C0F982",
 11017 => x"C0C0C0F9F9C0F9F8",
 11018 => x"C0C0C0F9F9C0F980",
 11019 => x"C0C0C0F9F9C0F990",
 11020 => x"C0C0C0F9F9C0A4C0",
 11021 => x"C0C0C0F9F9C0A4F9",
 11022 => x"C0C0C0F9F9C0A4A4",
 11023 => x"C0C0C0F9F9C0A4B0",
 11024 => x"C0C0C0F9F9C0A499",
 11025 => x"C0C0C0F9F9C0A492",
 11026 => x"C0C0C0F9F9C0A482",
 11027 => x"C0C0C0F9F9C0A4F8",
 11028 => x"C0C0C0F9F9C0A480",
 11029 => x"C0C0C0F9F9C0A490",
 11030 => x"C0C0C0F9F9C0B0C0",
 11031 => x"C0C0C0F9F9C0B0F9",
 11032 => x"C0C0C0F9F9C0B0A4",
 11033 => x"C0C0C0F9F9C0B0B0",
 11034 => x"C0C0C0F9F9C0B099",
 11035 => x"C0C0C0F9F9C0B092",
 11036 => x"C0C0C0F9F9C0B082",
 11037 => x"C0C0C0F9F9C0B0F8",
 11038 => x"C0C0C0F9F9C0B080",
 11039 => x"C0C0C0F9F9C0B090",
 11040 => x"C0C0C0F9F9C099C0",
 11041 => x"C0C0C0F9F9C099F9",
 11042 => x"C0C0C0F9F9C099A4",
 11043 => x"C0C0C0F9F9C099B0",
 11044 => x"C0C0C0F9F9C09999",
 11045 => x"C0C0C0F9F9C09992",
 11046 => x"C0C0C0F9F9C09982",
 11047 => x"C0C0C0F9F9C099F8",
 11048 => x"C0C0C0F9F9C09980",
 11049 => x"C0C0C0F9F9C09990",
 11050 => x"C0C0C0F9F9C092C0",
 11051 => x"C0C0C0F9F9C092F9",
 11052 => x"C0C0C0F9F9C092A4",
 11053 => x"C0C0C0F9F9C092B0",
 11054 => x"C0C0C0F9F9C09299",
 11055 => x"C0C0C0F9F9C09292",
 11056 => x"C0C0C0F9F9C09282",
 11057 => x"C0C0C0F9F9C092F8",
 11058 => x"C0C0C0F9F9C09280",
 11059 => x"C0C0C0F9F9C09290",
 11060 => x"C0C0C0F9F9C082C0",
 11061 => x"C0C0C0F9F9C082F9",
 11062 => x"C0C0C0F9F9C082A4",
 11063 => x"C0C0C0F9F9C082B0",
 11064 => x"C0C0C0F9F9C08299",
 11065 => x"C0C0C0F9F9C08292",
 11066 => x"C0C0C0F9F9C08282",
 11067 => x"C0C0C0F9F9C082F8",
 11068 => x"C0C0C0F9F9C08280",
 11069 => x"C0C0C0F9F9C08290",
 11070 => x"C0C0C0F9F9C0F8C0",
 11071 => x"C0C0C0F9F9C0F8F9",
 11072 => x"C0C0C0F9F9C0F8A4",
 11073 => x"C0C0C0F9F9C0F8B0",
 11074 => x"C0C0C0F9F9C0F899",
 11075 => x"C0C0C0F9F9C0F892",
 11076 => x"C0C0C0F9F9C0F882",
 11077 => x"C0C0C0F9F9C0F8F8",
 11078 => x"C0C0C0F9F9C0F880",
 11079 => x"C0C0C0F9F9C0F890",
 11080 => x"C0C0C0F9F9C080C0",
 11081 => x"C0C0C0F9F9C080F9",
 11082 => x"C0C0C0F9F9C080A4",
 11083 => x"C0C0C0F9F9C080B0",
 11084 => x"C0C0C0F9F9C08099",
 11085 => x"C0C0C0F9F9C08092",
 11086 => x"C0C0C0F9F9C08082",
 11087 => x"C0C0C0F9F9C080F8",
 11088 => x"C0C0C0F9F9C08080",
 11089 => x"C0C0C0F9F9C08090",
 11090 => x"C0C0C0F9F9C090C0",
 11091 => x"C0C0C0F9F9C090F9",
 11092 => x"C0C0C0F9F9C090A4",
 11093 => x"C0C0C0F9F9C090B0",
 11094 => x"C0C0C0F9F9C09099",
 11095 => x"C0C0C0F9F9C09092",
 11096 => x"C0C0C0F9F9C09082",
 11097 => x"C0C0C0F9F9C090F8",
 11098 => x"C0C0C0F9F9C09080",
 11099 => x"C0C0C0F9F9C09090",
 11100 => x"C0C0C0F9F9F9C0C0",
 11101 => x"C0C0C0F9F9F9C0F9",
 11102 => x"C0C0C0F9F9F9C0A4",
 11103 => x"C0C0C0F9F9F9C0B0",
 11104 => x"C0C0C0F9F9F9C099",
 11105 => x"C0C0C0F9F9F9C092",
 11106 => x"C0C0C0F9F9F9C082",
 11107 => x"C0C0C0F9F9F9C0F8",
 11108 => x"C0C0C0F9F9F9C080",
 11109 => x"C0C0C0F9F9F9C090",
 11110 => x"C0C0C0F9F9F9F9C0",
 11111 => x"C0C0C0F9F9F9F9F9",
 11112 => x"C0C0C0F9F9F9F9A4",
 11113 => x"C0C0C0F9F9F9F9B0",
 11114 => x"C0C0C0F9F9F9F999",
 11115 => x"C0C0C0F9F9F9F992",
 11116 => x"C0C0C0F9F9F9F982",
 11117 => x"C0C0C0F9F9F9F9F8",
 11118 => x"C0C0C0F9F9F9F980",
 11119 => x"C0C0C0F9F9F9F990",
 11120 => x"C0C0C0F9F9F9A4C0",
 11121 => x"C0C0C0F9F9F9A4F9",
 11122 => x"C0C0C0F9F9F9A4A4",
 11123 => x"C0C0C0F9F9F9A4B0",
 11124 => x"C0C0C0F9F9F9A499",
 11125 => x"C0C0C0F9F9F9A492",
 11126 => x"C0C0C0F9F9F9A482",
 11127 => x"C0C0C0F9F9F9A4F8",
 11128 => x"C0C0C0F9F9F9A480",
 11129 => x"C0C0C0F9F9F9A490",
 11130 => x"C0C0C0F9F9F9B0C0",
 11131 => x"C0C0C0F9F9F9B0F9",
 11132 => x"C0C0C0F9F9F9B0A4",
 11133 => x"C0C0C0F9F9F9B0B0",
 11134 => x"C0C0C0F9F9F9B099",
 11135 => x"C0C0C0F9F9F9B092",
 11136 => x"C0C0C0F9F9F9B082",
 11137 => x"C0C0C0F9F9F9B0F8",
 11138 => x"C0C0C0F9F9F9B080",
 11139 => x"C0C0C0F9F9F9B090",
 11140 => x"C0C0C0F9F9F999C0",
 11141 => x"C0C0C0F9F9F999F9",
 11142 => x"C0C0C0F9F9F999A4",
 11143 => x"C0C0C0F9F9F999B0",
 11144 => x"C0C0C0F9F9F99999",
 11145 => x"C0C0C0F9F9F99992",
 11146 => x"C0C0C0F9F9F99982",
 11147 => x"C0C0C0F9F9F999F8",
 11148 => x"C0C0C0F9F9F99980",
 11149 => x"C0C0C0F9F9F99990",
 11150 => x"C0C0C0F9F9F992C0",
 11151 => x"C0C0C0F9F9F992F9",
 11152 => x"C0C0C0F9F9F992A4",
 11153 => x"C0C0C0F9F9F992B0",
 11154 => x"C0C0C0F9F9F99299",
 11155 => x"C0C0C0F9F9F99292",
 11156 => x"C0C0C0F9F9F99282",
 11157 => x"C0C0C0F9F9F992F8",
 11158 => x"C0C0C0F9F9F99280",
 11159 => x"C0C0C0F9F9F99290",
 11160 => x"C0C0C0F9F9F982C0",
 11161 => x"C0C0C0F9F9F982F9",
 11162 => x"C0C0C0F9F9F982A4",
 11163 => x"C0C0C0F9F9F982B0",
 11164 => x"C0C0C0F9F9F98299",
 11165 => x"C0C0C0F9F9F98292",
 11166 => x"C0C0C0F9F9F98282",
 11167 => x"C0C0C0F9F9F982F8",
 11168 => x"C0C0C0F9F9F98280",
 11169 => x"C0C0C0F9F9F98290",
 11170 => x"C0C0C0F9F9F9F8C0",
 11171 => x"C0C0C0F9F9F9F8F9",
 11172 => x"C0C0C0F9F9F9F8A4",
 11173 => x"C0C0C0F9F9F9F8B0",
 11174 => x"C0C0C0F9F9F9F899",
 11175 => x"C0C0C0F9F9F9F892",
 11176 => x"C0C0C0F9F9F9F882",
 11177 => x"C0C0C0F9F9F9F8F8",
 11178 => x"C0C0C0F9F9F9F880",
 11179 => x"C0C0C0F9F9F9F890",
 11180 => x"C0C0C0F9F9F980C0",
 11181 => x"C0C0C0F9F9F980F9",
 11182 => x"C0C0C0F9F9F980A4",
 11183 => x"C0C0C0F9F9F980B0",
 11184 => x"C0C0C0F9F9F98099",
 11185 => x"C0C0C0F9F9F98092",
 11186 => x"C0C0C0F9F9F98082",
 11187 => x"C0C0C0F9F9F980F8",
 11188 => x"C0C0C0F9F9F98080",
 11189 => x"C0C0C0F9F9F98090",
 11190 => x"C0C0C0F9F9F990C0",
 11191 => x"C0C0C0F9F9F990F9",
 11192 => x"C0C0C0F9F9F990A4",
 11193 => x"C0C0C0F9F9F990B0",
 11194 => x"C0C0C0F9F9F99099",
 11195 => x"C0C0C0F9F9F99092",
 11196 => x"C0C0C0F9F9F99082",
 11197 => x"C0C0C0F9F9F990F8",
 11198 => x"C0C0C0F9F9F99080",
 11199 => x"C0C0C0F9F9F99090",
 11200 => x"C0C0C0F9F9A4C0C0",
 11201 => x"C0C0C0F9F9A4C0F9",
 11202 => x"C0C0C0F9F9A4C0A4",
 11203 => x"C0C0C0F9F9A4C0B0",
 11204 => x"C0C0C0F9F9A4C099",
 11205 => x"C0C0C0F9F9A4C092",
 11206 => x"C0C0C0F9F9A4C082",
 11207 => x"C0C0C0F9F9A4C0F8",
 11208 => x"C0C0C0F9F9A4C080",
 11209 => x"C0C0C0F9F9A4C090",
 11210 => x"C0C0C0F9F9A4F9C0",
 11211 => x"C0C0C0F9F9A4F9F9",
 11212 => x"C0C0C0F9F9A4F9A4",
 11213 => x"C0C0C0F9F9A4F9B0",
 11214 => x"C0C0C0F9F9A4F999",
 11215 => x"C0C0C0F9F9A4F992",
 11216 => x"C0C0C0F9F9A4F982",
 11217 => x"C0C0C0F9F9A4F9F8",
 11218 => x"C0C0C0F9F9A4F980",
 11219 => x"C0C0C0F9F9A4F990",
 11220 => x"C0C0C0F9F9A4A4C0",
 11221 => x"C0C0C0F9F9A4A4F9",
 11222 => x"C0C0C0F9F9A4A4A4",
 11223 => x"C0C0C0F9F9A4A4B0",
 11224 => x"C0C0C0F9F9A4A499",
 11225 => x"C0C0C0F9F9A4A492",
 11226 => x"C0C0C0F9F9A4A482",
 11227 => x"C0C0C0F9F9A4A4F8",
 11228 => x"C0C0C0F9F9A4A480",
 11229 => x"C0C0C0F9F9A4A490",
 11230 => x"C0C0C0F9F9A4B0C0",
 11231 => x"C0C0C0F9F9A4B0F9",
 11232 => x"C0C0C0F9F9A4B0A4",
 11233 => x"C0C0C0F9F9A4B0B0",
 11234 => x"C0C0C0F9F9A4B099",
 11235 => x"C0C0C0F9F9A4B092",
 11236 => x"C0C0C0F9F9A4B082",
 11237 => x"C0C0C0F9F9A4B0F8",
 11238 => x"C0C0C0F9F9A4B080",
 11239 => x"C0C0C0F9F9A4B090",
 11240 => x"C0C0C0F9F9A499C0",
 11241 => x"C0C0C0F9F9A499F9",
 11242 => x"C0C0C0F9F9A499A4",
 11243 => x"C0C0C0F9F9A499B0",
 11244 => x"C0C0C0F9F9A49999",
 11245 => x"C0C0C0F9F9A49992",
 11246 => x"C0C0C0F9F9A49982",
 11247 => x"C0C0C0F9F9A499F8",
 11248 => x"C0C0C0F9F9A49980",
 11249 => x"C0C0C0F9F9A49990",
 11250 => x"C0C0C0F9F9A492C0",
 11251 => x"C0C0C0F9F9A492F9",
 11252 => x"C0C0C0F9F9A492A4",
 11253 => x"C0C0C0F9F9A492B0",
 11254 => x"C0C0C0F9F9A49299",
 11255 => x"C0C0C0F9F9A49292",
 11256 => x"C0C0C0F9F9A49282",
 11257 => x"C0C0C0F9F9A492F8",
 11258 => x"C0C0C0F9F9A49280",
 11259 => x"C0C0C0F9F9A49290",
 11260 => x"C0C0C0F9F9A482C0",
 11261 => x"C0C0C0F9F9A482F9",
 11262 => x"C0C0C0F9F9A482A4",
 11263 => x"C0C0C0F9F9A482B0",
 11264 => x"C0C0C0F9F9A48299",
 11265 => x"C0C0C0F9F9A48292",
 11266 => x"C0C0C0F9F9A48282",
 11267 => x"C0C0C0F9F9A482F8",
 11268 => x"C0C0C0F9F9A48280",
 11269 => x"C0C0C0F9F9A48290",
 11270 => x"C0C0C0F9F9A4F8C0",
 11271 => x"C0C0C0F9F9A4F8F9",
 11272 => x"C0C0C0F9F9A4F8A4",
 11273 => x"C0C0C0F9F9A4F8B0",
 11274 => x"C0C0C0F9F9A4F899",
 11275 => x"C0C0C0F9F9A4F892",
 11276 => x"C0C0C0F9F9A4F882",
 11277 => x"C0C0C0F9F9A4F8F8",
 11278 => x"C0C0C0F9F9A4F880",
 11279 => x"C0C0C0F9F9A4F890",
 11280 => x"C0C0C0F9F9A480C0",
 11281 => x"C0C0C0F9F9A480F9",
 11282 => x"C0C0C0F9F9A480A4",
 11283 => x"C0C0C0F9F9A480B0",
 11284 => x"C0C0C0F9F9A48099",
 11285 => x"C0C0C0F9F9A48092",
 11286 => x"C0C0C0F9F9A48082",
 11287 => x"C0C0C0F9F9A480F8",
 11288 => x"C0C0C0F9F9A48080",
 11289 => x"C0C0C0F9F9A48090",
 11290 => x"C0C0C0F9F9A490C0",
 11291 => x"C0C0C0F9F9A490F9",
 11292 => x"C0C0C0F9F9A490A4",
 11293 => x"C0C0C0F9F9A490B0",
 11294 => x"C0C0C0F9F9A49099",
 11295 => x"C0C0C0F9F9A49092",
 11296 => x"C0C0C0F9F9A49082",
 11297 => x"C0C0C0F9F9A490F8",
 11298 => x"C0C0C0F9F9A49080",
 11299 => x"C0C0C0F9F9A49090",
 11300 => x"C0C0C0F9F9B0C0C0",
 11301 => x"C0C0C0F9F9B0C0F9",
 11302 => x"C0C0C0F9F9B0C0A4",
 11303 => x"C0C0C0F9F9B0C0B0",
 11304 => x"C0C0C0F9F9B0C099",
 11305 => x"C0C0C0F9F9B0C092",
 11306 => x"C0C0C0F9F9B0C082",
 11307 => x"C0C0C0F9F9B0C0F8",
 11308 => x"C0C0C0F9F9B0C080",
 11309 => x"C0C0C0F9F9B0C090",
 11310 => x"C0C0C0F9F9B0F9C0",
 11311 => x"C0C0C0F9F9B0F9F9",
 11312 => x"C0C0C0F9F9B0F9A4",
 11313 => x"C0C0C0F9F9B0F9B0",
 11314 => x"C0C0C0F9F9B0F999",
 11315 => x"C0C0C0F9F9B0F992",
 11316 => x"C0C0C0F9F9B0F982",
 11317 => x"C0C0C0F9F9B0F9F8",
 11318 => x"C0C0C0F9F9B0F980",
 11319 => x"C0C0C0F9F9B0F990",
 11320 => x"C0C0C0F9F9B0A4C0",
 11321 => x"C0C0C0F9F9B0A4F9",
 11322 => x"C0C0C0F9F9B0A4A4",
 11323 => x"C0C0C0F9F9B0A4B0",
 11324 => x"C0C0C0F9F9B0A499",
 11325 => x"C0C0C0F9F9B0A492",
 11326 => x"C0C0C0F9F9B0A482",
 11327 => x"C0C0C0F9F9B0A4F8",
 11328 => x"C0C0C0F9F9B0A480",
 11329 => x"C0C0C0F9F9B0A490",
 11330 => x"C0C0C0F9F9B0B0C0",
 11331 => x"C0C0C0F9F9B0B0F9",
 11332 => x"C0C0C0F9F9B0B0A4",
 11333 => x"C0C0C0F9F9B0B0B0",
 11334 => x"C0C0C0F9F9B0B099",
 11335 => x"C0C0C0F9F9B0B092",
 11336 => x"C0C0C0F9F9B0B082",
 11337 => x"C0C0C0F9F9B0B0F8",
 11338 => x"C0C0C0F9F9B0B080",
 11339 => x"C0C0C0F9F9B0B090",
 11340 => x"C0C0C0F9F9B099C0",
 11341 => x"C0C0C0F9F9B099F9",
 11342 => x"C0C0C0F9F9B099A4",
 11343 => x"C0C0C0F9F9B099B0",
 11344 => x"C0C0C0F9F9B09999",
 11345 => x"C0C0C0F9F9B09992",
 11346 => x"C0C0C0F9F9B09982",
 11347 => x"C0C0C0F9F9B099F8",
 11348 => x"C0C0C0F9F9B09980",
 11349 => x"C0C0C0F9F9B09990",
 11350 => x"C0C0C0F9F9B092C0",
 11351 => x"C0C0C0F9F9B092F9",
 11352 => x"C0C0C0F9F9B092A4",
 11353 => x"C0C0C0F9F9B092B0",
 11354 => x"C0C0C0F9F9B09299",
 11355 => x"C0C0C0F9F9B09292",
 11356 => x"C0C0C0F9F9B09282",
 11357 => x"C0C0C0F9F9B092F8",
 11358 => x"C0C0C0F9F9B09280",
 11359 => x"C0C0C0F9F9B09290",
 11360 => x"C0C0C0F9F9B082C0",
 11361 => x"C0C0C0F9F9B082F9",
 11362 => x"C0C0C0F9F9B082A4",
 11363 => x"C0C0C0F9F9B082B0",
 11364 => x"C0C0C0F9F9B08299",
 11365 => x"C0C0C0F9F9B08292",
 11366 => x"C0C0C0F9F9B08282",
 11367 => x"C0C0C0F9F9B082F8",
 11368 => x"C0C0C0F9F9B08280",
 11369 => x"C0C0C0F9F9B08290",
 11370 => x"C0C0C0F9F9B0F8C0",
 11371 => x"C0C0C0F9F9B0F8F9",
 11372 => x"C0C0C0F9F9B0F8A4",
 11373 => x"C0C0C0F9F9B0F8B0",
 11374 => x"C0C0C0F9F9B0F899",
 11375 => x"C0C0C0F9F9B0F892",
 11376 => x"C0C0C0F9F9B0F882",
 11377 => x"C0C0C0F9F9B0F8F8",
 11378 => x"C0C0C0F9F9B0F880",
 11379 => x"C0C0C0F9F9B0F890",
 11380 => x"C0C0C0F9F9B080C0",
 11381 => x"C0C0C0F9F9B080F9",
 11382 => x"C0C0C0F9F9B080A4",
 11383 => x"C0C0C0F9F9B080B0",
 11384 => x"C0C0C0F9F9B08099",
 11385 => x"C0C0C0F9F9B08092",
 11386 => x"C0C0C0F9F9B08082",
 11387 => x"C0C0C0F9F9B080F8",
 11388 => x"C0C0C0F9F9B08080",
 11389 => x"C0C0C0F9F9B08090",
 11390 => x"C0C0C0F9F9B090C0",
 11391 => x"C0C0C0F9F9B090F9",
 11392 => x"C0C0C0F9F9B090A4",
 11393 => x"C0C0C0F9F9B090B0",
 11394 => x"C0C0C0F9F9B09099",
 11395 => x"C0C0C0F9F9B09092",
 11396 => x"C0C0C0F9F9B09082",
 11397 => x"C0C0C0F9F9B090F8",
 11398 => x"C0C0C0F9F9B09080",
 11399 => x"C0C0C0F9F9B09090",
 11400 => x"C0C0C0F9F999C0C0",
 11401 => x"C0C0C0F9F999C0F9",
 11402 => x"C0C0C0F9F999C0A4",
 11403 => x"C0C0C0F9F999C0B0",
 11404 => x"C0C0C0F9F999C099",
 11405 => x"C0C0C0F9F999C092",
 11406 => x"C0C0C0F9F999C082",
 11407 => x"C0C0C0F9F999C0F8",
 11408 => x"C0C0C0F9F999C080",
 11409 => x"C0C0C0F9F999C090",
 11410 => x"C0C0C0F9F999F9C0",
 11411 => x"C0C0C0F9F999F9F9",
 11412 => x"C0C0C0F9F999F9A4",
 11413 => x"C0C0C0F9F999F9B0",
 11414 => x"C0C0C0F9F999F999",
 11415 => x"C0C0C0F9F999F992",
 11416 => x"C0C0C0F9F999F982",
 11417 => x"C0C0C0F9F999F9F8",
 11418 => x"C0C0C0F9F999F980",
 11419 => x"C0C0C0F9F999F990",
 11420 => x"C0C0C0F9F999A4C0",
 11421 => x"C0C0C0F9F999A4F9",
 11422 => x"C0C0C0F9F999A4A4",
 11423 => x"C0C0C0F9F999A4B0",
 11424 => x"C0C0C0F9F999A499",
 11425 => x"C0C0C0F9F999A492",
 11426 => x"C0C0C0F9F999A482",
 11427 => x"C0C0C0F9F999A4F8",
 11428 => x"C0C0C0F9F999A480",
 11429 => x"C0C0C0F9F999A490",
 11430 => x"C0C0C0F9F999B0C0",
 11431 => x"C0C0C0F9F999B0F9",
 11432 => x"C0C0C0F9F999B0A4",
 11433 => x"C0C0C0F9F999B0B0",
 11434 => x"C0C0C0F9F999B099",
 11435 => x"C0C0C0F9F999B092",
 11436 => x"C0C0C0F9F999B082",
 11437 => x"C0C0C0F9F999B0F8",
 11438 => x"C0C0C0F9F999B080",
 11439 => x"C0C0C0F9F999B090",
 11440 => x"C0C0C0F9F99999C0",
 11441 => x"C0C0C0F9F99999F9",
 11442 => x"C0C0C0F9F99999A4",
 11443 => x"C0C0C0F9F99999B0",
 11444 => x"C0C0C0F9F9999999",
 11445 => x"C0C0C0F9F9999992",
 11446 => x"C0C0C0F9F9999982",
 11447 => x"C0C0C0F9F99999F8",
 11448 => x"C0C0C0F9F9999980",
 11449 => x"C0C0C0F9F9999990",
 11450 => x"C0C0C0F9F99992C0",
 11451 => x"C0C0C0F9F99992F9",
 11452 => x"C0C0C0F9F99992A4",
 11453 => x"C0C0C0F9F99992B0",
 11454 => x"C0C0C0F9F9999299",
 11455 => x"C0C0C0F9F9999292",
 11456 => x"C0C0C0F9F9999282",
 11457 => x"C0C0C0F9F99992F8",
 11458 => x"C0C0C0F9F9999280",
 11459 => x"C0C0C0F9F9999290",
 11460 => x"C0C0C0F9F99982C0",
 11461 => x"C0C0C0F9F99982F9",
 11462 => x"C0C0C0F9F99982A4",
 11463 => x"C0C0C0F9F99982B0",
 11464 => x"C0C0C0F9F9998299",
 11465 => x"C0C0C0F9F9998292",
 11466 => x"C0C0C0F9F9998282",
 11467 => x"C0C0C0F9F99982F8",
 11468 => x"C0C0C0F9F9998280",
 11469 => x"C0C0C0F9F9998290",
 11470 => x"C0C0C0F9F999F8C0",
 11471 => x"C0C0C0F9F999F8F9",
 11472 => x"C0C0C0F9F999F8A4",
 11473 => x"C0C0C0F9F999F8B0",
 11474 => x"C0C0C0F9F999F899",
 11475 => x"C0C0C0F9F999F892",
 11476 => x"C0C0C0F9F999F882",
 11477 => x"C0C0C0F9F999F8F8",
 11478 => x"C0C0C0F9F999F880",
 11479 => x"C0C0C0F9F999F890",
 11480 => x"C0C0C0F9F99980C0",
 11481 => x"C0C0C0F9F99980F9",
 11482 => x"C0C0C0F9F99980A4",
 11483 => x"C0C0C0F9F99980B0",
 11484 => x"C0C0C0F9F9998099",
 11485 => x"C0C0C0F9F9998092",
 11486 => x"C0C0C0F9F9998082",
 11487 => x"C0C0C0F9F99980F8",
 11488 => x"C0C0C0F9F9998080",
 11489 => x"C0C0C0F9F9998090",
 11490 => x"C0C0C0F9F99990C0",
 11491 => x"C0C0C0F9F99990F9",
 11492 => x"C0C0C0F9F99990A4",
 11493 => x"C0C0C0F9F99990B0",
 11494 => x"C0C0C0F9F9999099",
 11495 => x"C0C0C0F9F9999092",
 11496 => x"C0C0C0F9F9999082",
 11497 => x"C0C0C0F9F99990F8",
 11498 => x"C0C0C0F9F9999080",
 11499 => x"C0C0C0F9F9999090",
 11500 => x"C0C0C0F9F992C0C0",
 11501 => x"C0C0C0F9F992C0F9",
 11502 => x"C0C0C0F9F992C0A4",
 11503 => x"C0C0C0F9F992C0B0",
 11504 => x"C0C0C0F9F992C099",
 11505 => x"C0C0C0F9F992C092",
 11506 => x"C0C0C0F9F992C082",
 11507 => x"C0C0C0F9F992C0F8",
 11508 => x"C0C0C0F9F992C080",
 11509 => x"C0C0C0F9F992C090",
 11510 => x"C0C0C0F9F992F9C0",
 11511 => x"C0C0C0F9F992F9F9",
 11512 => x"C0C0C0F9F992F9A4",
 11513 => x"C0C0C0F9F992F9B0",
 11514 => x"C0C0C0F9F992F999",
 11515 => x"C0C0C0F9F992F992",
 11516 => x"C0C0C0F9F992F982",
 11517 => x"C0C0C0F9F992F9F8",
 11518 => x"C0C0C0F9F992F980",
 11519 => x"C0C0C0F9F992F990",
 11520 => x"C0C0C0F9F992A4C0",
 11521 => x"C0C0C0F9F992A4F9",
 11522 => x"C0C0C0F9F992A4A4",
 11523 => x"C0C0C0F9F992A4B0",
 11524 => x"C0C0C0F9F992A499",
 11525 => x"C0C0C0F9F992A492",
 11526 => x"C0C0C0F9F992A482",
 11527 => x"C0C0C0F9F992A4F8",
 11528 => x"C0C0C0F9F992A480",
 11529 => x"C0C0C0F9F992A490",
 11530 => x"C0C0C0F9F992B0C0",
 11531 => x"C0C0C0F9F992B0F9",
 11532 => x"C0C0C0F9F992B0A4",
 11533 => x"C0C0C0F9F992B0B0",
 11534 => x"C0C0C0F9F992B099",
 11535 => x"C0C0C0F9F992B092",
 11536 => x"C0C0C0F9F992B082",
 11537 => x"C0C0C0F9F992B0F8",
 11538 => x"C0C0C0F9F992B080",
 11539 => x"C0C0C0F9F992B090",
 11540 => x"C0C0C0F9F99299C0",
 11541 => x"C0C0C0F9F99299F9",
 11542 => x"C0C0C0F9F99299A4",
 11543 => x"C0C0C0F9F99299B0",
 11544 => x"C0C0C0F9F9929999",
 11545 => x"C0C0C0F9F9929992",
 11546 => x"C0C0C0F9F9929982",
 11547 => x"C0C0C0F9F99299F8",
 11548 => x"C0C0C0F9F9929980",
 11549 => x"C0C0C0F9F9929990",
 11550 => x"C0C0C0F9F99292C0",
 11551 => x"C0C0C0F9F99292F9",
 11552 => x"C0C0C0F9F99292A4",
 11553 => x"C0C0C0F9F99292B0",
 11554 => x"C0C0C0F9F9929299",
 11555 => x"C0C0C0F9F9929292",
 11556 => x"C0C0C0F9F9929282",
 11557 => x"C0C0C0F9F99292F8",
 11558 => x"C0C0C0F9F9929280",
 11559 => x"C0C0C0F9F9929290",
 11560 => x"C0C0C0F9F99282C0",
 11561 => x"C0C0C0F9F99282F9",
 11562 => x"C0C0C0F9F99282A4",
 11563 => x"C0C0C0F9F99282B0",
 11564 => x"C0C0C0F9F9928299",
 11565 => x"C0C0C0F9F9928292",
 11566 => x"C0C0C0F9F9928282",
 11567 => x"C0C0C0F9F99282F8",
 11568 => x"C0C0C0F9F9928280",
 11569 => x"C0C0C0F9F9928290",
 11570 => x"C0C0C0F9F992F8C0",
 11571 => x"C0C0C0F9F992F8F9",
 11572 => x"C0C0C0F9F992F8A4",
 11573 => x"C0C0C0F9F992F8B0",
 11574 => x"C0C0C0F9F992F899",
 11575 => x"C0C0C0F9F992F892",
 11576 => x"C0C0C0F9F992F882",
 11577 => x"C0C0C0F9F992F8F8",
 11578 => x"C0C0C0F9F992F880",
 11579 => x"C0C0C0F9F992F890",
 11580 => x"C0C0C0F9F99280C0",
 11581 => x"C0C0C0F9F99280F9",
 11582 => x"C0C0C0F9F99280A4",
 11583 => x"C0C0C0F9F99280B0",
 11584 => x"C0C0C0F9F9928099",
 11585 => x"C0C0C0F9F9928092",
 11586 => x"C0C0C0F9F9928082",
 11587 => x"C0C0C0F9F99280F8",
 11588 => x"C0C0C0F9F9928080",
 11589 => x"C0C0C0F9F9928090",
 11590 => x"C0C0C0F9F99290C0",
 11591 => x"C0C0C0F9F99290F9",
 11592 => x"C0C0C0F9F99290A4",
 11593 => x"C0C0C0F9F99290B0",
 11594 => x"C0C0C0F9F9929099",
 11595 => x"C0C0C0F9F9929092",
 11596 => x"C0C0C0F9F9929082",
 11597 => x"C0C0C0F9F99290F8",
 11598 => x"C0C0C0F9F9929080",
 11599 => x"C0C0C0F9F9929090",
 11600 => x"C0C0C0F9F982C0C0",
 11601 => x"C0C0C0F9F982C0F9",
 11602 => x"C0C0C0F9F982C0A4",
 11603 => x"C0C0C0F9F982C0B0",
 11604 => x"C0C0C0F9F982C099",
 11605 => x"C0C0C0F9F982C092",
 11606 => x"C0C0C0F9F982C082",
 11607 => x"C0C0C0F9F982C0F8",
 11608 => x"C0C0C0F9F982C080",
 11609 => x"C0C0C0F9F982C090",
 11610 => x"C0C0C0F9F982F9C0",
 11611 => x"C0C0C0F9F982F9F9",
 11612 => x"C0C0C0F9F982F9A4",
 11613 => x"C0C0C0F9F982F9B0",
 11614 => x"C0C0C0F9F982F999",
 11615 => x"C0C0C0F9F982F992",
 11616 => x"C0C0C0F9F982F982",
 11617 => x"C0C0C0F9F982F9F8",
 11618 => x"C0C0C0F9F982F980",
 11619 => x"C0C0C0F9F982F990",
 11620 => x"C0C0C0F9F982A4C0",
 11621 => x"C0C0C0F9F982A4F9",
 11622 => x"C0C0C0F9F982A4A4",
 11623 => x"C0C0C0F9F982A4B0",
 11624 => x"C0C0C0F9F982A499",
 11625 => x"C0C0C0F9F982A492",
 11626 => x"C0C0C0F9F982A482",
 11627 => x"C0C0C0F9F982A4F8",
 11628 => x"C0C0C0F9F982A480",
 11629 => x"C0C0C0F9F982A490",
 11630 => x"C0C0C0F9F982B0C0",
 11631 => x"C0C0C0F9F982B0F9",
 11632 => x"C0C0C0F9F982B0A4",
 11633 => x"C0C0C0F9F982B0B0",
 11634 => x"C0C0C0F9F982B099",
 11635 => x"C0C0C0F9F982B092",
 11636 => x"C0C0C0F9F982B082",
 11637 => x"C0C0C0F9F982B0F8",
 11638 => x"C0C0C0F9F982B080",
 11639 => x"C0C0C0F9F982B090",
 11640 => x"C0C0C0F9F98299C0",
 11641 => x"C0C0C0F9F98299F9",
 11642 => x"C0C0C0F9F98299A4",
 11643 => x"C0C0C0F9F98299B0",
 11644 => x"C0C0C0F9F9829999",
 11645 => x"C0C0C0F9F9829992",
 11646 => x"C0C0C0F9F9829982",
 11647 => x"C0C0C0F9F98299F8",
 11648 => x"C0C0C0F9F9829980",
 11649 => x"C0C0C0F9F9829990",
 11650 => x"C0C0C0F9F98292C0",
 11651 => x"C0C0C0F9F98292F9",
 11652 => x"C0C0C0F9F98292A4",
 11653 => x"C0C0C0F9F98292B0",
 11654 => x"C0C0C0F9F9829299",
 11655 => x"C0C0C0F9F9829292",
 11656 => x"C0C0C0F9F9829282",
 11657 => x"C0C0C0F9F98292F8",
 11658 => x"C0C0C0F9F9829280",
 11659 => x"C0C0C0F9F9829290",
 11660 => x"C0C0C0F9F98282C0",
 11661 => x"C0C0C0F9F98282F9",
 11662 => x"C0C0C0F9F98282A4",
 11663 => x"C0C0C0F9F98282B0",
 11664 => x"C0C0C0F9F9828299",
 11665 => x"C0C0C0F9F9828292",
 11666 => x"C0C0C0F9F9828282",
 11667 => x"C0C0C0F9F98282F8",
 11668 => x"C0C0C0F9F9828280",
 11669 => x"C0C0C0F9F9828290",
 11670 => x"C0C0C0F9F982F8C0",
 11671 => x"C0C0C0F9F982F8F9",
 11672 => x"C0C0C0F9F982F8A4",
 11673 => x"C0C0C0F9F982F8B0",
 11674 => x"C0C0C0F9F982F899",
 11675 => x"C0C0C0F9F982F892",
 11676 => x"C0C0C0F9F982F882",
 11677 => x"C0C0C0F9F982F8F8",
 11678 => x"C0C0C0F9F982F880",
 11679 => x"C0C0C0F9F982F890",
 11680 => x"C0C0C0F9F98280C0",
 11681 => x"C0C0C0F9F98280F9",
 11682 => x"C0C0C0F9F98280A4",
 11683 => x"C0C0C0F9F98280B0",
 11684 => x"C0C0C0F9F9828099",
 11685 => x"C0C0C0F9F9828092",
 11686 => x"C0C0C0F9F9828082",
 11687 => x"C0C0C0F9F98280F8",
 11688 => x"C0C0C0F9F9828080",
 11689 => x"C0C0C0F9F9828090",
 11690 => x"C0C0C0F9F98290C0",
 11691 => x"C0C0C0F9F98290F9",
 11692 => x"C0C0C0F9F98290A4",
 11693 => x"C0C0C0F9F98290B0",
 11694 => x"C0C0C0F9F9829099",
 11695 => x"C0C0C0F9F9829092",
 11696 => x"C0C0C0F9F9829082",
 11697 => x"C0C0C0F9F98290F8",
 11698 => x"C0C0C0F9F9829080",
 11699 => x"C0C0C0F9F9829090",
 11700 => x"C0C0C0F9F9F8C0C0",
 11701 => x"C0C0C0F9F9F8C0F9",
 11702 => x"C0C0C0F9F9F8C0A4",
 11703 => x"C0C0C0F9F9F8C0B0",
 11704 => x"C0C0C0F9F9F8C099",
 11705 => x"C0C0C0F9F9F8C092",
 11706 => x"C0C0C0F9F9F8C082",
 11707 => x"C0C0C0F9F9F8C0F8",
 11708 => x"C0C0C0F9F9F8C080",
 11709 => x"C0C0C0F9F9F8C090",
 11710 => x"C0C0C0F9F9F8F9C0",
 11711 => x"C0C0C0F9F9F8F9F9",
 11712 => x"C0C0C0F9F9F8F9A4",
 11713 => x"C0C0C0F9F9F8F9B0",
 11714 => x"C0C0C0F9F9F8F999",
 11715 => x"C0C0C0F9F9F8F992",
 11716 => x"C0C0C0F9F9F8F982",
 11717 => x"C0C0C0F9F9F8F9F8",
 11718 => x"C0C0C0F9F9F8F980",
 11719 => x"C0C0C0F9F9F8F990",
 11720 => x"C0C0C0F9F9F8A4C0",
 11721 => x"C0C0C0F9F9F8A4F9",
 11722 => x"C0C0C0F9F9F8A4A4",
 11723 => x"C0C0C0F9F9F8A4B0",
 11724 => x"C0C0C0F9F9F8A499",
 11725 => x"C0C0C0F9F9F8A492",
 11726 => x"C0C0C0F9F9F8A482",
 11727 => x"C0C0C0F9F9F8A4F8",
 11728 => x"C0C0C0F9F9F8A480",
 11729 => x"C0C0C0F9F9F8A490",
 11730 => x"C0C0C0F9F9F8B0C0",
 11731 => x"C0C0C0F9F9F8B0F9",
 11732 => x"C0C0C0F9F9F8B0A4",
 11733 => x"C0C0C0F9F9F8B0B0",
 11734 => x"C0C0C0F9F9F8B099",
 11735 => x"C0C0C0F9F9F8B092",
 11736 => x"C0C0C0F9F9F8B082",
 11737 => x"C0C0C0F9F9F8B0F8",
 11738 => x"C0C0C0F9F9F8B080",
 11739 => x"C0C0C0F9F9F8B090",
 11740 => x"C0C0C0F9F9F899C0",
 11741 => x"C0C0C0F9F9F899F9",
 11742 => x"C0C0C0F9F9F899A4",
 11743 => x"C0C0C0F9F9F899B0",
 11744 => x"C0C0C0F9F9F89999",
 11745 => x"C0C0C0F9F9F89992",
 11746 => x"C0C0C0F9F9F89982",
 11747 => x"C0C0C0F9F9F899F8",
 11748 => x"C0C0C0F9F9F89980",
 11749 => x"C0C0C0F9F9F89990",
 11750 => x"C0C0C0F9F9F892C0",
 11751 => x"C0C0C0F9F9F892F9",
 11752 => x"C0C0C0F9F9F892A4",
 11753 => x"C0C0C0F9F9F892B0",
 11754 => x"C0C0C0F9F9F89299",
 11755 => x"C0C0C0F9F9F89292",
 11756 => x"C0C0C0F9F9F89282",
 11757 => x"C0C0C0F9F9F892F8",
 11758 => x"C0C0C0F9F9F89280",
 11759 => x"C0C0C0F9F9F89290",
 11760 => x"C0C0C0F9F9F882C0",
 11761 => x"C0C0C0F9F9F882F9",
 11762 => x"C0C0C0F9F9F882A4",
 11763 => x"C0C0C0F9F9F882B0",
 11764 => x"C0C0C0F9F9F88299",
 11765 => x"C0C0C0F9F9F88292",
 11766 => x"C0C0C0F9F9F88282",
 11767 => x"C0C0C0F9F9F882F8",
 11768 => x"C0C0C0F9F9F88280",
 11769 => x"C0C0C0F9F9F88290",
 11770 => x"C0C0C0F9F9F8F8C0",
 11771 => x"C0C0C0F9F9F8F8F9",
 11772 => x"C0C0C0F9F9F8F8A4",
 11773 => x"C0C0C0F9F9F8F8B0",
 11774 => x"C0C0C0F9F9F8F899",
 11775 => x"C0C0C0F9F9F8F892",
 11776 => x"C0C0C0F9F9F8F882",
 11777 => x"C0C0C0F9F9F8F8F8",
 11778 => x"C0C0C0F9F9F8F880",
 11779 => x"C0C0C0F9F9F8F890",
 11780 => x"C0C0C0F9F9F880C0",
 11781 => x"C0C0C0F9F9F880F9",
 11782 => x"C0C0C0F9F9F880A4",
 11783 => x"C0C0C0F9F9F880B0",
 11784 => x"C0C0C0F9F9F88099",
 11785 => x"C0C0C0F9F9F88092",
 11786 => x"C0C0C0F9F9F88082",
 11787 => x"C0C0C0F9F9F880F8",
 11788 => x"C0C0C0F9F9F88080",
 11789 => x"C0C0C0F9F9F88090",
 11790 => x"C0C0C0F9F9F890C0",
 11791 => x"C0C0C0F9F9F890F9",
 11792 => x"C0C0C0F9F9F890A4",
 11793 => x"C0C0C0F9F9F890B0",
 11794 => x"C0C0C0F9F9F89099",
 11795 => x"C0C0C0F9F9F89092",
 11796 => x"C0C0C0F9F9F89082",
 11797 => x"C0C0C0F9F9F890F8",
 11798 => x"C0C0C0F9F9F89080",
 11799 => x"C0C0C0F9F9F89090",
 11800 => x"C0C0C0F9F980C0C0",
 11801 => x"C0C0C0F9F980C0F9",
 11802 => x"C0C0C0F9F980C0A4",
 11803 => x"C0C0C0F9F980C0B0",
 11804 => x"C0C0C0F9F980C099",
 11805 => x"C0C0C0F9F980C092",
 11806 => x"C0C0C0F9F980C082",
 11807 => x"C0C0C0F9F980C0F8",
 11808 => x"C0C0C0F9F980C080",
 11809 => x"C0C0C0F9F980C090",
 11810 => x"C0C0C0F9F980F9C0",
 11811 => x"C0C0C0F9F980F9F9",
 11812 => x"C0C0C0F9F980F9A4",
 11813 => x"C0C0C0F9F980F9B0",
 11814 => x"C0C0C0F9F980F999",
 11815 => x"C0C0C0F9F980F992",
 11816 => x"C0C0C0F9F980F982",
 11817 => x"C0C0C0F9F980F9F8",
 11818 => x"C0C0C0F9F980F980",
 11819 => x"C0C0C0F9F980F990",
 11820 => x"C0C0C0F9F980A4C0",
 11821 => x"C0C0C0F9F980A4F9",
 11822 => x"C0C0C0F9F980A4A4",
 11823 => x"C0C0C0F9F980A4B0",
 11824 => x"C0C0C0F9F980A499",
 11825 => x"C0C0C0F9F980A492",
 11826 => x"C0C0C0F9F980A482",
 11827 => x"C0C0C0F9F980A4F8",
 11828 => x"C0C0C0F9F980A480",
 11829 => x"C0C0C0F9F980A490",
 11830 => x"C0C0C0F9F980B0C0",
 11831 => x"C0C0C0F9F980B0F9",
 11832 => x"C0C0C0F9F980B0A4",
 11833 => x"C0C0C0F9F980B0B0",
 11834 => x"C0C0C0F9F980B099",
 11835 => x"C0C0C0F9F980B092",
 11836 => x"C0C0C0F9F980B082",
 11837 => x"C0C0C0F9F980B0F8",
 11838 => x"C0C0C0F9F980B080",
 11839 => x"C0C0C0F9F980B090",
 11840 => x"C0C0C0F9F98099C0",
 11841 => x"C0C0C0F9F98099F9",
 11842 => x"C0C0C0F9F98099A4",
 11843 => x"C0C0C0F9F98099B0",
 11844 => x"C0C0C0F9F9809999",
 11845 => x"C0C0C0F9F9809992",
 11846 => x"C0C0C0F9F9809982",
 11847 => x"C0C0C0F9F98099F8",
 11848 => x"C0C0C0F9F9809980",
 11849 => x"C0C0C0F9F9809990",
 11850 => x"C0C0C0F9F98092C0",
 11851 => x"C0C0C0F9F98092F9",
 11852 => x"C0C0C0F9F98092A4",
 11853 => x"C0C0C0F9F98092B0",
 11854 => x"C0C0C0F9F9809299",
 11855 => x"C0C0C0F9F9809292",
 11856 => x"C0C0C0F9F9809282",
 11857 => x"C0C0C0F9F98092F8",
 11858 => x"C0C0C0F9F9809280",
 11859 => x"C0C0C0F9F9809290",
 11860 => x"C0C0C0F9F98082C0",
 11861 => x"C0C0C0F9F98082F9",
 11862 => x"C0C0C0F9F98082A4",
 11863 => x"C0C0C0F9F98082B0",
 11864 => x"C0C0C0F9F9808299",
 11865 => x"C0C0C0F9F9808292",
 11866 => x"C0C0C0F9F9808282",
 11867 => x"C0C0C0F9F98082F8",
 11868 => x"C0C0C0F9F9808280",
 11869 => x"C0C0C0F9F9808290",
 11870 => x"C0C0C0F9F980F8C0",
 11871 => x"C0C0C0F9F980F8F9",
 11872 => x"C0C0C0F9F980F8A4",
 11873 => x"C0C0C0F9F980F8B0",
 11874 => x"C0C0C0F9F980F899",
 11875 => x"C0C0C0F9F980F892",
 11876 => x"C0C0C0F9F980F882",
 11877 => x"C0C0C0F9F980F8F8",
 11878 => x"C0C0C0F9F980F880",
 11879 => x"C0C0C0F9F980F890",
 11880 => x"C0C0C0F9F98080C0",
 11881 => x"C0C0C0F9F98080F9",
 11882 => x"C0C0C0F9F98080A4",
 11883 => x"C0C0C0F9F98080B0",
 11884 => x"C0C0C0F9F9808099",
 11885 => x"C0C0C0F9F9808092",
 11886 => x"C0C0C0F9F9808082",
 11887 => x"C0C0C0F9F98080F8",
 11888 => x"C0C0C0F9F9808080",
 11889 => x"C0C0C0F9F9808090",
 11890 => x"C0C0C0F9F98090C0",
 11891 => x"C0C0C0F9F98090F9",
 11892 => x"C0C0C0F9F98090A4",
 11893 => x"C0C0C0F9F98090B0",
 11894 => x"C0C0C0F9F9809099",
 11895 => x"C0C0C0F9F9809092",
 11896 => x"C0C0C0F9F9809082",
 11897 => x"C0C0C0F9F98090F8",
 11898 => x"C0C0C0F9F9809080",
 11899 => x"C0C0C0F9F9809090",
 11900 => x"C0C0C0F9F990C0C0",
 11901 => x"C0C0C0F9F990C0F9",
 11902 => x"C0C0C0F9F990C0A4",
 11903 => x"C0C0C0F9F990C0B0",
 11904 => x"C0C0C0F9F990C099",
 11905 => x"C0C0C0F9F990C092",
 11906 => x"C0C0C0F9F990C082",
 11907 => x"C0C0C0F9F990C0F8",
 11908 => x"C0C0C0F9F990C080",
 11909 => x"C0C0C0F9F990C090",
 11910 => x"C0C0C0F9F990F9C0",
 11911 => x"C0C0C0F9F990F9F9",
 11912 => x"C0C0C0F9F990F9A4",
 11913 => x"C0C0C0F9F990F9B0",
 11914 => x"C0C0C0F9F990F999",
 11915 => x"C0C0C0F9F990F992",
 11916 => x"C0C0C0F9F990F982",
 11917 => x"C0C0C0F9F990F9F8",
 11918 => x"C0C0C0F9F990F980",
 11919 => x"C0C0C0F9F990F990",
 11920 => x"C0C0C0F9F990A4C0",
 11921 => x"C0C0C0F9F990A4F9",
 11922 => x"C0C0C0F9F990A4A4",
 11923 => x"C0C0C0F9F990A4B0",
 11924 => x"C0C0C0F9F990A499",
 11925 => x"C0C0C0F9F990A492",
 11926 => x"C0C0C0F9F990A482",
 11927 => x"C0C0C0F9F990A4F8",
 11928 => x"C0C0C0F9F990A480",
 11929 => x"C0C0C0F9F990A490",
 11930 => x"C0C0C0F9F990B0C0",
 11931 => x"C0C0C0F9F990B0F9",
 11932 => x"C0C0C0F9F990B0A4",
 11933 => x"C0C0C0F9F990B0B0",
 11934 => x"C0C0C0F9F990B099",
 11935 => x"C0C0C0F9F990B092",
 11936 => x"C0C0C0F9F990B082",
 11937 => x"C0C0C0F9F990B0F8",
 11938 => x"C0C0C0F9F990B080",
 11939 => x"C0C0C0F9F990B090",
 11940 => x"C0C0C0F9F99099C0",
 11941 => x"C0C0C0F9F99099F9",
 11942 => x"C0C0C0F9F99099A4",
 11943 => x"C0C0C0F9F99099B0",
 11944 => x"C0C0C0F9F9909999",
 11945 => x"C0C0C0F9F9909992",
 11946 => x"C0C0C0F9F9909982",
 11947 => x"C0C0C0F9F99099F8",
 11948 => x"C0C0C0F9F9909980",
 11949 => x"C0C0C0F9F9909990",
 11950 => x"C0C0C0F9F99092C0",
 11951 => x"C0C0C0F9F99092F9",
 11952 => x"C0C0C0F9F99092A4",
 11953 => x"C0C0C0F9F99092B0",
 11954 => x"C0C0C0F9F9909299",
 11955 => x"C0C0C0F9F9909292",
 11956 => x"C0C0C0F9F9909282",
 11957 => x"C0C0C0F9F99092F8",
 11958 => x"C0C0C0F9F9909280",
 11959 => x"C0C0C0F9F9909290",
 11960 => x"C0C0C0F9F99082C0",
 11961 => x"C0C0C0F9F99082F9",
 11962 => x"C0C0C0F9F99082A4",
 11963 => x"C0C0C0F9F99082B0",
 11964 => x"C0C0C0F9F9908299",
 11965 => x"C0C0C0F9F9908292",
 11966 => x"C0C0C0F9F9908282",
 11967 => x"C0C0C0F9F99082F8",
 11968 => x"C0C0C0F9F9908280",
 11969 => x"C0C0C0F9F9908290",
 11970 => x"C0C0C0F9F990F8C0",
 11971 => x"C0C0C0F9F990F8F9",
 11972 => x"C0C0C0F9F990F8A4",
 11973 => x"C0C0C0F9F990F8B0",
 11974 => x"C0C0C0F9F990F899",
 11975 => x"C0C0C0F9F990F892",
 11976 => x"C0C0C0F9F990F882",
 11977 => x"C0C0C0F9F990F8F8",
 11978 => x"C0C0C0F9F990F880",
 11979 => x"C0C0C0F9F990F890",
 11980 => x"C0C0C0F9F99080C0",
 11981 => x"C0C0C0F9F99080F9",
 11982 => x"C0C0C0F9F99080A4",
 11983 => x"C0C0C0F9F99080B0",
 11984 => x"C0C0C0F9F9908099",
 11985 => x"C0C0C0F9F9908092",
 11986 => x"C0C0C0F9F9908082",
 11987 => x"C0C0C0F9F99080F8",
 11988 => x"C0C0C0F9F9908080",
 11989 => x"C0C0C0F9F9908090",
 11990 => x"C0C0C0F9F99090C0",
 11991 => x"C0C0C0F9F99090F9",
 11992 => x"C0C0C0F9F99090A4",
 11993 => x"C0C0C0F9F99090B0",
 11994 => x"C0C0C0F9F9909099",
 11995 => x"C0C0C0F9F9909092",
 11996 => x"C0C0C0F9F9909082",
 11997 => x"C0C0C0F9F99090F8",
 11998 => x"C0C0C0F9F9909080",
 11999 => x"C0C0C0F9F9909090",
 12000 => x"C0C0C0F9A4C0C0C0",
 12001 => x"C0C0C0F9A4C0C0F9",
 12002 => x"C0C0C0F9A4C0C0A4",
 12003 => x"C0C0C0F9A4C0C0B0",
 12004 => x"C0C0C0F9A4C0C099",
 12005 => x"C0C0C0F9A4C0C092",
 12006 => x"C0C0C0F9A4C0C082",
 12007 => x"C0C0C0F9A4C0C0F8",
 12008 => x"C0C0C0F9A4C0C080",
 12009 => x"C0C0C0F9A4C0C090",
 12010 => x"C0C0C0F9A4C0F9C0",
 12011 => x"C0C0C0F9A4C0F9F9",
 12012 => x"C0C0C0F9A4C0F9A4",
 12013 => x"C0C0C0F9A4C0F9B0",
 12014 => x"C0C0C0F9A4C0F999",
 12015 => x"C0C0C0F9A4C0F992",
 12016 => x"C0C0C0F9A4C0F982",
 12017 => x"C0C0C0F9A4C0F9F8",
 12018 => x"C0C0C0F9A4C0F980",
 12019 => x"C0C0C0F9A4C0F990",
 12020 => x"C0C0C0F9A4C0A4C0",
 12021 => x"C0C0C0F9A4C0A4F9",
 12022 => x"C0C0C0F9A4C0A4A4",
 12023 => x"C0C0C0F9A4C0A4B0",
 12024 => x"C0C0C0F9A4C0A499",
 12025 => x"C0C0C0F9A4C0A492",
 12026 => x"C0C0C0F9A4C0A482",
 12027 => x"C0C0C0F9A4C0A4F8",
 12028 => x"C0C0C0F9A4C0A480",
 12029 => x"C0C0C0F9A4C0A490",
 12030 => x"C0C0C0F9A4C0B0C0",
 12031 => x"C0C0C0F9A4C0B0F9",
 12032 => x"C0C0C0F9A4C0B0A4",
 12033 => x"C0C0C0F9A4C0B0B0",
 12034 => x"C0C0C0F9A4C0B099",
 12035 => x"C0C0C0F9A4C0B092",
 12036 => x"C0C0C0F9A4C0B082",
 12037 => x"C0C0C0F9A4C0B0F8",
 12038 => x"C0C0C0F9A4C0B080",
 12039 => x"C0C0C0F9A4C0B090",
 12040 => x"C0C0C0F9A4C099C0",
 12041 => x"C0C0C0F9A4C099F9",
 12042 => x"C0C0C0F9A4C099A4",
 12043 => x"C0C0C0F9A4C099B0",
 12044 => x"C0C0C0F9A4C09999",
 12045 => x"C0C0C0F9A4C09992",
 12046 => x"C0C0C0F9A4C09982",
 12047 => x"C0C0C0F9A4C099F8",
 12048 => x"C0C0C0F9A4C09980",
 12049 => x"C0C0C0F9A4C09990",
 12050 => x"C0C0C0F9A4C092C0",
 12051 => x"C0C0C0F9A4C092F9",
 12052 => x"C0C0C0F9A4C092A4",
 12053 => x"C0C0C0F9A4C092B0",
 12054 => x"C0C0C0F9A4C09299",
 12055 => x"C0C0C0F9A4C09292",
 12056 => x"C0C0C0F9A4C09282",
 12057 => x"C0C0C0F9A4C092F8",
 12058 => x"C0C0C0F9A4C09280",
 12059 => x"C0C0C0F9A4C09290",
 12060 => x"C0C0C0F9A4C082C0",
 12061 => x"C0C0C0F9A4C082F9",
 12062 => x"C0C0C0F9A4C082A4",
 12063 => x"C0C0C0F9A4C082B0",
 12064 => x"C0C0C0F9A4C08299",
 12065 => x"C0C0C0F9A4C08292",
 12066 => x"C0C0C0F9A4C08282",
 12067 => x"C0C0C0F9A4C082F8",
 12068 => x"C0C0C0F9A4C08280",
 12069 => x"C0C0C0F9A4C08290",
 12070 => x"C0C0C0F9A4C0F8C0",
 12071 => x"C0C0C0F9A4C0F8F9",
 12072 => x"C0C0C0F9A4C0F8A4",
 12073 => x"C0C0C0F9A4C0F8B0",
 12074 => x"C0C0C0F9A4C0F899",
 12075 => x"C0C0C0F9A4C0F892",
 12076 => x"C0C0C0F9A4C0F882",
 12077 => x"C0C0C0F9A4C0F8F8",
 12078 => x"C0C0C0F9A4C0F880",
 12079 => x"C0C0C0F9A4C0F890",
 12080 => x"C0C0C0F9A4C080C0",
 12081 => x"C0C0C0F9A4C080F9",
 12082 => x"C0C0C0F9A4C080A4",
 12083 => x"C0C0C0F9A4C080B0",
 12084 => x"C0C0C0F9A4C08099",
 12085 => x"C0C0C0F9A4C08092",
 12086 => x"C0C0C0F9A4C08082",
 12087 => x"C0C0C0F9A4C080F8",
 12088 => x"C0C0C0F9A4C08080",
 12089 => x"C0C0C0F9A4C08090",
 12090 => x"C0C0C0F9A4C090C0",
 12091 => x"C0C0C0F9A4C090F9",
 12092 => x"C0C0C0F9A4C090A4",
 12093 => x"C0C0C0F9A4C090B0",
 12094 => x"C0C0C0F9A4C09099",
 12095 => x"C0C0C0F9A4C09092",
 12096 => x"C0C0C0F9A4C09082",
 12097 => x"C0C0C0F9A4C090F8",
 12098 => x"C0C0C0F9A4C09080",
 12099 => x"C0C0C0F9A4C09090",
 12100 => x"C0C0C0F9A4F9C0C0",
 12101 => x"C0C0C0F9A4F9C0F9",
 12102 => x"C0C0C0F9A4F9C0A4",
 12103 => x"C0C0C0F9A4F9C0B0",
 12104 => x"C0C0C0F9A4F9C099",
 12105 => x"C0C0C0F9A4F9C092",
 12106 => x"C0C0C0F9A4F9C082",
 12107 => x"C0C0C0F9A4F9C0F8",
 12108 => x"C0C0C0F9A4F9C080",
 12109 => x"C0C0C0F9A4F9C090",
 12110 => x"C0C0C0F9A4F9F9C0",
 12111 => x"C0C0C0F9A4F9F9F9",
 12112 => x"C0C0C0F9A4F9F9A4",
 12113 => x"C0C0C0F9A4F9F9B0",
 12114 => x"C0C0C0F9A4F9F999",
 12115 => x"C0C0C0F9A4F9F992",
 12116 => x"C0C0C0F9A4F9F982",
 12117 => x"C0C0C0F9A4F9F9F8",
 12118 => x"C0C0C0F9A4F9F980",
 12119 => x"C0C0C0F9A4F9F990",
 12120 => x"C0C0C0F9A4F9A4C0",
 12121 => x"C0C0C0F9A4F9A4F9",
 12122 => x"C0C0C0F9A4F9A4A4",
 12123 => x"C0C0C0F9A4F9A4B0",
 12124 => x"C0C0C0F9A4F9A499",
 12125 => x"C0C0C0F9A4F9A492",
 12126 => x"C0C0C0F9A4F9A482",
 12127 => x"C0C0C0F9A4F9A4F8",
 12128 => x"C0C0C0F9A4F9A480",
 12129 => x"C0C0C0F9A4F9A490",
 12130 => x"C0C0C0F9A4F9B0C0",
 12131 => x"C0C0C0F9A4F9B0F9",
 12132 => x"C0C0C0F9A4F9B0A4",
 12133 => x"C0C0C0F9A4F9B0B0",
 12134 => x"C0C0C0F9A4F9B099",
 12135 => x"C0C0C0F9A4F9B092",
 12136 => x"C0C0C0F9A4F9B082",
 12137 => x"C0C0C0F9A4F9B0F8",
 12138 => x"C0C0C0F9A4F9B080",
 12139 => x"C0C0C0F9A4F9B090",
 12140 => x"C0C0C0F9A4F999C0",
 12141 => x"C0C0C0F9A4F999F9",
 12142 => x"C0C0C0F9A4F999A4",
 12143 => x"C0C0C0F9A4F999B0",
 12144 => x"C0C0C0F9A4F99999",
 12145 => x"C0C0C0F9A4F99992",
 12146 => x"C0C0C0F9A4F99982",
 12147 => x"C0C0C0F9A4F999F8",
 12148 => x"C0C0C0F9A4F99980",
 12149 => x"C0C0C0F9A4F99990",
 12150 => x"C0C0C0F9A4F992C0",
 12151 => x"C0C0C0F9A4F992F9",
 12152 => x"C0C0C0F9A4F992A4",
 12153 => x"C0C0C0F9A4F992B0",
 12154 => x"C0C0C0F9A4F99299",
 12155 => x"C0C0C0F9A4F99292",
 12156 => x"C0C0C0F9A4F99282",
 12157 => x"C0C0C0F9A4F992F8",
 12158 => x"C0C0C0F9A4F99280",
 12159 => x"C0C0C0F9A4F99290",
 12160 => x"C0C0C0F9A4F982C0",
 12161 => x"C0C0C0F9A4F982F9",
 12162 => x"C0C0C0F9A4F982A4",
 12163 => x"C0C0C0F9A4F982B0",
 12164 => x"C0C0C0F9A4F98299",
 12165 => x"C0C0C0F9A4F98292",
 12166 => x"C0C0C0F9A4F98282",
 12167 => x"C0C0C0F9A4F982F8",
 12168 => x"C0C0C0F9A4F98280",
 12169 => x"C0C0C0F9A4F98290",
 12170 => x"C0C0C0F9A4F9F8C0",
 12171 => x"C0C0C0F9A4F9F8F9",
 12172 => x"C0C0C0F9A4F9F8A4",
 12173 => x"C0C0C0F9A4F9F8B0",
 12174 => x"C0C0C0F9A4F9F899",
 12175 => x"C0C0C0F9A4F9F892",
 12176 => x"C0C0C0F9A4F9F882",
 12177 => x"C0C0C0F9A4F9F8F8",
 12178 => x"C0C0C0F9A4F9F880",
 12179 => x"C0C0C0F9A4F9F890",
 12180 => x"C0C0C0F9A4F980C0",
 12181 => x"C0C0C0F9A4F980F9",
 12182 => x"C0C0C0F9A4F980A4",
 12183 => x"C0C0C0F9A4F980B0",
 12184 => x"C0C0C0F9A4F98099",
 12185 => x"C0C0C0F9A4F98092",
 12186 => x"C0C0C0F9A4F98082",
 12187 => x"C0C0C0F9A4F980F8",
 12188 => x"C0C0C0F9A4F98080",
 12189 => x"C0C0C0F9A4F98090",
 12190 => x"C0C0C0F9A4F990C0",
 12191 => x"C0C0C0F9A4F990F9",
 12192 => x"C0C0C0F9A4F990A4",
 12193 => x"C0C0C0F9A4F990B0",
 12194 => x"C0C0C0F9A4F99099",
 12195 => x"C0C0C0F9A4F99092",
 12196 => x"C0C0C0F9A4F99082",
 12197 => x"C0C0C0F9A4F990F8",
 12198 => x"C0C0C0F9A4F99080",
 12199 => x"C0C0C0F9A4F99090",
 12200 => x"C0C0C0F9A4A4C0C0",
 12201 => x"C0C0C0F9A4A4C0F9",
 12202 => x"C0C0C0F9A4A4C0A4",
 12203 => x"C0C0C0F9A4A4C0B0",
 12204 => x"C0C0C0F9A4A4C099",
 12205 => x"C0C0C0F9A4A4C092",
 12206 => x"C0C0C0F9A4A4C082",
 12207 => x"C0C0C0F9A4A4C0F8",
 12208 => x"C0C0C0F9A4A4C080",
 12209 => x"C0C0C0F9A4A4C090",
 12210 => x"C0C0C0F9A4A4F9C0",
 12211 => x"C0C0C0F9A4A4F9F9",
 12212 => x"C0C0C0F9A4A4F9A4",
 12213 => x"C0C0C0F9A4A4F9B0",
 12214 => x"C0C0C0F9A4A4F999",
 12215 => x"C0C0C0F9A4A4F992",
 12216 => x"C0C0C0F9A4A4F982",
 12217 => x"C0C0C0F9A4A4F9F8",
 12218 => x"C0C0C0F9A4A4F980",
 12219 => x"C0C0C0F9A4A4F990",
 12220 => x"C0C0C0F9A4A4A4C0",
 12221 => x"C0C0C0F9A4A4A4F9",
 12222 => x"C0C0C0F9A4A4A4A4",
 12223 => x"C0C0C0F9A4A4A4B0",
 12224 => x"C0C0C0F9A4A4A499",
 12225 => x"C0C0C0F9A4A4A492",
 12226 => x"C0C0C0F9A4A4A482",
 12227 => x"C0C0C0F9A4A4A4F8",
 12228 => x"C0C0C0F9A4A4A480",
 12229 => x"C0C0C0F9A4A4A490",
 12230 => x"C0C0C0F9A4A4B0C0",
 12231 => x"C0C0C0F9A4A4B0F9",
 12232 => x"C0C0C0F9A4A4B0A4",
 12233 => x"C0C0C0F9A4A4B0B0",
 12234 => x"C0C0C0F9A4A4B099",
 12235 => x"C0C0C0F9A4A4B092",
 12236 => x"C0C0C0F9A4A4B082",
 12237 => x"C0C0C0F9A4A4B0F8",
 12238 => x"C0C0C0F9A4A4B080",
 12239 => x"C0C0C0F9A4A4B090",
 12240 => x"C0C0C0F9A4A499C0",
 12241 => x"C0C0C0F9A4A499F9",
 12242 => x"C0C0C0F9A4A499A4",
 12243 => x"C0C0C0F9A4A499B0",
 12244 => x"C0C0C0F9A4A49999",
 12245 => x"C0C0C0F9A4A49992",
 12246 => x"C0C0C0F9A4A49982",
 12247 => x"C0C0C0F9A4A499F8",
 12248 => x"C0C0C0F9A4A49980",
 12249 => x"C0C0C0F9A4A49990",
 12250 => x"C0C0C0F9A4A492C0",
 12251 => x"C0C0C0F9A4A492F9",
 12252 => x"C0C0C0F9A4A492A4",
 12253 => x"C0C0C0F9A4A492B0",
 12254 => x"C0C0C0F9A4A49299",
 12255 => x"C0C0C0F9A4A49292",
 12256 => x"C0C0C0F9A4A49282",
 12257 => x"C0C0C0F9A4A492F8",
 12258 => x"C0C0C0F9A4A49280",
 12259 => x"C0C0C0F9A4A49290",
 12260 => x"C0C0C0F9A4A482C0",
 12261 => x"C0C0C0F9A4A482F9",
 12262 => x"C0C0C0F9A4A482A4",
 12263 => x"C0C0C0F9A4A482B0",
 12264 => x"C0C0C0F9A4A48299",
 12265 => x"C0C0C0F9A4A48292",
 12266 => x"C0C0C0F9A4A48282",
 12267 => x"C0C0C0F9A4A482F8",
 12268 => x"C0C0C0F9A4A48280",
 12269 => x"C0C0C0F9A4A48290",
 12270 => x"C0C0C0F9A4A4F8C0",
 12271 => x"C0C0C0F9A4A4F8F9",
 12272 => x"C0C0C0F9A4A4F8A4",
 12273 => x"C0C0C0F9A4A4F8B0",
 12274 => x"C0C0C0F9A4A4F899",
 12275 => x"C0C0C0F9A4A4F892",
 12276 => x"C0C0C0F9A4A4F882",
 12277 => x"C0C0C0F9A4A4F8F8",
 12278 => x"C0C0C0F9A4A4F880",
 12279 => x"C0C0C0F9A4A4F890",
 12280 => x"C0C0C0F9A4A480C0",
 12281 => x"C0C0C0F9A4A480F9",
 12282 => x"C0C0C0F9A4A480A4",
 12283 => x"C0C0C0F9A4A480B0",
 12284 => x"C0C0C0F9A4A48099",
 12285 => x"C0C0C0F9A4A48092",
 12286 => x"C0C0C0F9A4A48082",
 12287 => x"C0C0C0F9A4A480F8",
 12288 => x"C0C0C0F9A4A48080",
 12289 => x"C0C0C0F9A4A48090",
 12290 => x"C0C0C0F9A4A490C0",
 12291 => x"C0C0C0F9A4A490F9",
 12292 => x"C0C0C0F9A4A490A4",
 12293 => x"C0C0C0F9A4A490B0",
 12294 => x"C0C0C0F9A4A49099",
 12295 => x"C0C0C0F9A4A49092",
 12296 => x"C0C0C0F9A4A49082",
 12297 => x"C0C0C0F9A4A490F8",
 12298 => x"C0C0C0F9A4A49080",
 12299 => x"C0C0C0F9A4A49090",
 12300 => x"C0C0C0F9A4B0C0C0",
 12301 => x"C0C0C0F9A4B0C0F9",
 12302 => x"C0C0C0F9A4B0C0A4",
 12303 => x"C0C0C0F9A4B0C0B0",
 12304 => x"C0C0C0F9A4B0C099",
 12305 => x"C0C0C0F9A4B0C092",
 12306 => x"C0C0C0F9A4B0C082",
 12307 => x"C0C0C0F9A4B0C0F8",
 12308 => x"C0C0C0F9A4B0C080",
 12309 => x"C0C0C0F9A4B0C090",
 12310 => x"C0C0C0F9A4B0F9C0",
 12311 => x"C0C0C0F9A4B0F9F9",
 12312 => x"C0C0C0F9A4B0F9A4",
 12313 => x"C0C0C0F9A4B0F9B0",
 12314 => x"C0C0C0F9A4B0F999",
 12315 => x"C0C0C0F9A4B0F992",
 12316 => x"C0C0C0F9A4B0F982",
 12317 => x"C0C0C0F9A4B0F9F8",
 12318 => x"C0C0C0F9A4B0F980",
 12319 => x"C0C0C0F9A4B0F990",
 12320 => x"C0C0C0F9A4B0A4C0",
 12321 => x"C0C0C0F9A4B0A4F9",
 12322 => x"C0C0C0F9A4B0A4A4",
 12323 => x"C0C0C0F9A4B0A4B0",
 12324 => x"C0C0C0F9A4B0A499",
 12325 => x"C0C0C0F9A4B0A492",
 12326 => x"C0C0C0F9A4B0A482",
 12327 => x"C0C0C0F9A4B0A4F8",
 12328 => x"C0C0C0F9A4B0A480",
 12329 => x"C0C0C0F9A4B0A490",
 12330 => x"C0C0C0F9A4B0B0C0",
 12331 => x"C0C0C0F9A4B0B0F9",
 12332 => x"C0C0C0F9A4B0B0A4",
 12333 => x"C0C0C0F9A4B0B0B0",
 12334 => x"C0C0C0F9A4B0B099",
 12335 => x"C0C0C0F9A4B0B092",
 12336 => x"C0C0C0F9A4B0B082",
 12337 => x"C0C0C0F9A4B0B0F8",
 12338 => x"C0C0C0F9A4B0B080",
 12339 => x"C0C0C0F9A4B0B090",
 12340 => x"C0C0C0F9A4B099C0",
 12341 => x"C0C0C0F9A4B099F9",
 12342 => x"C0C0C0F9A4B099A4",
 12343 => x"C0C0C0F9A4B099B0",
 12344 => x"C0C0C0F9A4B09999",
 12345 => x"C0C0C0F9A4B09992",
 12346 => x"C0C0C0F9A4B09982",
 12347 => x"C0C0C0F9A4B099F8",
 12348 => x"C0C0C0F9A4B09980",
 12349 => x"C0C0C0F9A4B09990",
 12350 => x"C0C0C0F9A4B092C0",
 12351 => x"C0C0C0F9A4B092F9",
 12352 => x"C0C0C0F9A4B092A4",
 12353 => x"C0C0C0F9A4B092B0",
 12354 => x"C0C0C0F9A4B09299",
 12355 => x"C0C0C0F9A4B09292",
 12356 => x"C0C0C0F9A4B09282",
 12357 => x"C0C0C0F9A4B092F8",
 12358 => x"C0C0C0F9A4B09280",
 12359 => x"C0C0C0F9A4B09290",
 12360 => x"C0C0C0F9A4B082C0",
 12361 => x"C0C0C0F9A4B082F9",
 12362 => x"C0C0C0F9A4B082A4",
 12363 => x"C0C0C0F9A4B082B0",
 12364 => x"C0C0C0F9A4B08299",
 12365 => x"C0C0C0F9A4B08292",
 12366 => x"C0C0C0F9A4B08282",
 12367 => x"C0C0C0F9A4B082F8",
 12368 => x"C0C0C0F9A4B08280",
 12369 => x"C0C0C0F9A4B08290",
 12370 => x"C0C0C0F9A4B0F8C0",
 12371 => x"C0C0C0F9A4B0F8F9",
 12372 => x"C0C0C0F9A4B0F8A4",
 12373 => x"C0C0C0F9A4B0F8B0",
 12374 => x"C0C0C0F9A4B0F899",
 12375 => x"C0C0C0F9A4B0F892",
 12376 => x"C0C0C0F9A4B0F882",
 12377 => x"C0C0C0F9A4B0F8F8",
 12378 => x"C0C0C0F9A4B0F880",
 12379 => x"C0C0C0F9A4B0F890",
 12380 => x"C0C0C0F9A4B080C0",
 12381 => x"C0C0C0F9A4B080F9",
 12382 => x"C0C0C0F9A4B080A4",
 12383 => x"C0C0C0F9A4B080B0",
 12384 => x"C0C0C0F9A4B08099",
 12385 => x"C0C0C0F9A4B08092",
 12386 => x"C0C0C0F9A4B08082",
 12387 => x"C0C0C0F9A4B080F8",
 12388 => x"C0C0C0F9A4B08080",
 12389 => x"C0C0C0F9A4B08090",
 12390 => x"C0C0C0F9A4B090C0",
 12391 => x"C0C0C0F9A4B090F9",
 12392 => x"C0C0C0F9A4B090A4",
 12393 => x"C0C0C0F9A4B090B0",
 12394 => x"C0C0C0F9A4B09099",
 12395 => x"C0C0C0F9A4B09092",
 12396 => x"C0C0C0F9A4B09082",
 12397 => x"C0C0C0F9A4B090F8",
 12398 => x"C0C0C0F9A4B09080",
 12399 => x"C0C0C0F9A4B09090",
 12400 => x"C0C0C0F9A499C0C0",
 12401 => x"C0C0C0F9A499C0F9",
 12402 => x"C0C0C0F9A499C0A4",
 12403 => x"C0C0C0F9A499C0B0",
 12404 => x"C0C0C0F9A499C099",
 12405 => x"C0C0C0F9A499C092",
 12406 => x"C0C0C0F9A499C082",
 12407 => x"C0C0C0F9A499C0F8",
 12408 => x"C0C0C0F9A499C080",
 12409 => x"C0C0C0F9A499C090",
 12410 => x"C0C0C0F9A499F9C0",
 12411 => x"C0C0C0F9A499F9F9",
 12412 => x"C0C0C0F9A499F9A4",
 12413 => x"C0C0C0F9A499F9B0",
 12414 => x"C0C0C0F9A499F999",
 12415 => x"C0C0C0F9A499F992",
 12416 => x"C0C0C0F9A499F982",
 12417 => x"C0C0C0F9A499F9F8",
 12418 => x"C0C0C0F9A499F980",
 12419 => x"C0C0C0F9A499F990",
 12420 => x"C0C0C0F9A499A4C0",
 12421 => x"C0C0C0F9A499A4F9",
 12422 => x"C0C0C0F9A499A4A4",
 12423 => x"C0C0C0F9A499A4B0",
 12424 => x"C0C0C0F9A499A499",
 12425 => x"C0C0C0F9A499A492",
 12426 => x"C0C0C0F9A499A482",
 12427 => x"C0C0C0F9A499A4F8",
 12428 => x"C0C0C0F9A499A480",
 12429 => x"C0C0C0F9A499A490",
 12430 => x"C0C0C0F9A499B0C0",
 12431 => x"C0C0C0F9A499B0F9",
 12432 => x"C0C0C0F9A499B0A4",
 12433 => x"C0C0C0F9A499B0B0",
 12434 => x"C0C0C0F9A499B099",
 12435 => x"C0C0C0F9A499B092",
 12436 => x"C0C0C0F9A499B082",
 12437 => x"C0C0C0F9A499B0F8",
 12438 => x"C0C0C0F9A499B080",
 12439 => x"C0C0C0F9A499B090",
 12440 => x"C0C0C0F9A49999C0",
 12441 => x"C0C0C0F9A49999F9",
 12442 => x"C0C0C0F9A49999A4",
 12443 => x"C0C0C0F9A49999B0",
 12444 => x"C0C0C0F9A4999999",
 12445 => x"C0C0C0F9A4999992",
 12446 => x"C0C0C0F9A4999982",
 12447 => x"C0C0C0F9A49999F8",
 12448 => x"C0C0C0F9A4999980",
 12449 => x"C0C0C0F9A4999990",
 12450 => x"C0C0C0F9A49992C0",
 12451 => x"C0C0C0F9A49992F9",
 12452 => x"C0C0C0F9A49992A4",
 12453 => x"C0C0C0F9A49992B0",
 12454 => x"C0C0C0F9A4999299",
 12455 => x"C0C0C0F9A4999292",
 12456 => x"C0C0C0F9A4999282",
 12457 => x"C0C0C0F9A49992F8",
 12458 => x"C0C0C0F9A4999280",
 12459 => x"C0C0C0F9A4999290",
 12460 => x"C0C0C0F9A49982C0",
 12461 => x"C0C0C0F9A49982F9",
 12462 => x"C0C0C0F9A49982A4",
 12463 => x"C0C0C0F9A49982B0",
 12464 => x"C0C0C0F9A4998299",
 12465 => x"C0C0C0F9A4998292",
 12466 => x"C0C0C0F9A4998282",
 12467 => x"C0C0C0F9A49982F8",
 12468 => x"C0C0C0F9A4998280",
 12469 => x"C0C0C0F9A4998290",
 12470 => x"C0C0C0F9A499F8C0",
 12471 => x"C0C0C0F9A499F8F9",
 12472 => x"C0C0C0F9A499F8A4",
 12473 => x"C0C0C0F9A499F8B0",
 12474 => x"C0C0C0F9A499F899",
 12475 => x"C0C0C0F9A499F892",
 12476 => x"C0C0C0F9A499F882",
 12477 => x"C0C0C0F9A499F8F8",
 12478 => x"C0C0C0F9A499F880",
 12479 => x"C0C0C0F9A499F890",
 12480 => x"C0C0C0F9A49980C0",
 12481 => x"C0C0C0F9A49980F9",
 12482 => x"C0C0C0F9A49980A4",
 12483 => x"C0C0C0F9A49980B0",
 12484 => x"C0C0C0F9A4998099",
 12485 => x"C0C0C0F9A4998092",
 12486 => x"C0C0C0F9A4998082",
 12487 => x"C0C0C0F9A49980F8",
 12488 => x"C0C0C0F9A4998080",
 12489 => x"C0C0C0F9A4998090",
 12490 => x"C0C0C0F9A49990C0",
 12491 => x"C0C0C0F9A49990F9",
 12492 => x"C0C0C0F9A49990A4",
 12493 => x"C0C0C0F9A49990B0",
 12494 => x"C0C0C0F9A4999099",
 12495 => x"C0C0C0F9A4999092",
 12496 => x"C0C0C0F9A4999082",
 12497 => x"C0C0C0F9A49990F8",
 12498 => x"C0C0C0F9A4999080",
 12499 => x"C0C0C0F9A4999090",
 12500 => x"C0C0C0F9A492C0C0",
 12501 => x"C0C0C0F9A492C0F9",
 12502 => x"C0C0C0F9A492C0A4",
 12503 => x"C0C0C0F9A492C0B0",
 12504 => x"C0C0C0F9A492C099",
 12505 => x"C0C0C0F9A492C092",
 12506 => x"C0C0C0F9A492C082",
 12507 => x"C0C0C0F9A492C0F8",
 12508 => x"C0C0C0F9A492C080",
 12509 => x"C0C0C0F9A492C090",
 12510 => x"C0C0C0F9A492F9C0",
 12511 => x"C0C0C0F9A492F9F9",
 12512 => x"C0C0C0F9A492F9A4",
 12513 => x"C0C0C0F9A492F9B0",
 12514 => x"C0C0C0F9A492F999",
 12515 => x"C0C0C0F9A492F992",
 12516 => x"C0C0C0F9A492F982",
 12517 => x"C0C0C0F9A492F9F8",
 12518 => x"C0C0C0F9A492F980",
 12519 => x"C0C0C0F9A492F990",
 12520 => x"C0C0C0F9A492A4C0",
 12521 => x"C0C0C0F9A492A4F9",
 12522 => x"C0C0C0F9A492A4A4",
 12523 => x"C0C0C0F9A492A4B0",
 12524 => x"C0C0C0F9A492A499",
 12525 => x"C0C0C0F9A492A492",
 12526 => x"C0C0C0F9A492A482",
 12527 => x"C0C0C0F9A492A4F8",
 12528 => x"C0C0C0F9A492A480",
 12529 => x"C0C0C0F9A492A490",
 12530 => x"C0C0C0F9A492B0C0",
 12531 => x"C0C0C0F9A492B0F9",
 12532 => x"C0C0C0F9A492B0A4",
 12533 => x"C0C0C0F9A492B0B0",
 12534 => x"C0C0C0F9A492B099",
 12535 => x"C0C0C0F9A492B092",
 12536 => x"C0C0C0F9A492B082",
 12537 => x"C0C0C0F9A492B0F8",
 12538 => x"C0C0C0F9A492B080",
 12539 => x"C0C0C0F9A492B090",
 12540 => x"C0C0C0F9A49299C0",
 12541 => x"C0C0C0F9A49299F9",
 12542 => x"C0C0C0F9A49299A4",
 12543 => x"C0C0C0F9A49299B0",
 12544 => x"C0C0C0F9A4929999",
 12545 => x"C0C0C0F9A4929992",
 12546 => x"C0C0C0F9A4929982",
 12547 => x"C0C0C0F9A49299F8",
 12548 => x"C0C0C0F9A4929980",
 12549 => x"C0C0C0F9A4929990",
 12550 => x"C0C0C0F9A49292C0",
 12551 => x"C0C0C0F9A49292F9",
 12552 => x"C0C0C0F9A49292A4",
 12553 => x"C0C0C0F9A49292B0",
 12554 => x"C0C0C0F9A4929299",
 12555 => x"C0C0C0F9A4929292",
 12556 => x"C0C0C0F9A4929282",
 12557 => x"C0C0C0F9A49292F8",
 12558 => x"C0C0C0F9A4929280",
 12559 => x"C0C0C0F9A4929290",
 12560 => x"C0C0C0F9A49282C0",
 12561 => x"C0C0C0F9A49282F9",
 12562 => x"C0C0C0F9A49282A4",
 12563 => x"C0C0C0F9A49282B0",
 12564 => x"C0C0C0F9A4928299",
 12565 => x"C0C0C0F9A4928292",
 12566 => x"C0C0C0F9A4928282",
 12567 => x"C0C0C0F9A49282F8",
 12568 => x"C0C0C0F9A4928280",
 12569 => x"C0C0C0F9A4928290",
 12570 => x"C0C0C0F9A492F8C0",
 12571 => x"C0C0C0F9A492F8F9",
 12572 => x"C0C0C0F9A492F8A4",
 12573 => x"C0C0C0F9A492F8B0",
 12574 => x"C0C0C0F9A492F899",
 12575 => x"C0C0C0F9A492F892",
 12576 => x"C0C0C0F9A492F882",
 12577 => x"C0C0C0F9A492F8F8",
 12578 => x"C0C0C0F9A492F880",
 12579 => x"C0C0C0F9A492F890",
 12580 => x"C0C0C0F9A49280C0",
 12581 => x"C0C0C0F9A49280F9",
 12582 => x"C0C0C0F9A49280A4",
 12583 => x"C0C0C0F9A49280B0",
 12584 => x"C0C0C0F9A4928099",
 12585 => x"C0C0C0F9A4928092",
 12586 => x"C0C0C0F9A4928082",
 12587 => x"C0C0C0F9A49280F8",
 12588 => x"C0C0C0F9A4928080",
 12589 => x"C0C0C0F9A4928090",
 12590 => x"C0C0C0F9A49290C0",
 12591 => x"C0C0C0F9A49290F9",
 12592 => x"C0C0C0F9A49290A4",
 12593 => x"C0C0C0F9A49290B0",
 12594 => x"C0C0C0F9A4929099",
 12595 => x"C0C0C0F9A4929092",
 12596 => x"C0C0C0F9A4929082",
 12597 => x"C0C0C0F9A49290F8",
 12598 => x"C0C0C0F9A4929080",
 12599 => x"C0C0C0F9A4929090",
 12600 => x"C0C0C0F9A482C0C0",
 12601 => x"C0C0C0F9A482C0F9",
 12602 => x"C0C0C0F9A482C0A4",
 12603 => x"C0C0C0F9A482C0B0",
 12604 => x"C0C0C0F9A482C099",
 12605 => x"C0C0C0F9A482C092",
 12606 => x"C0C0C0F9A482C082",
 12607 => x"C0C0C0F9A482C0F8",
 12608 => x"C0C0C0F9A482C080",
 12609 => x"C0C0C0F9A482C090",
 12610 => x"C0C0C0F9A482F9C0",
 12611 => x"C0C0C0F9A482F9F9",
 12612 => x"C0C0C0F9A482F9A4",
 12613 => x"C0C0C0F9A482F9B0",
 12614 => x"C0C0C0F9A482F999",
 12615 => x"C0C0C0F9A482F992",
 12616 => x"C0C0C0F9A482F982",
 12617 => x"C0C0C0F9A482F9F8",
 12618 => x"C0C0C0F9A482F980",
 12619 => x"C0C0C0F9A482F990",
 12620 => x"C0C0C0F9A482A4C0",
 12621 => x"C0C0C0F9A482A4F9",
 12622 => x"C0C0C0F9A482A4A4",
 12623 => x"C0C0C0F9A482A4B0",
 12624 => x"C0C0C0F9A482A499",
 12625 => x"C0C0C0F9A482A492",
 12626 => x"C0C0C0F9A482A482",
 12627 => x"C0C0C0F9A482A4F8",
 12628 => x"C0C0C0F9A482A480",
 12629 => x"C0C0C0F9A482A490",
 12630 => x"C0C0C0F9A482B0C0",
 12631 => x"C0C0C0F9A482B0F9",
 12632 => x"C0C0C0F9A482B0A4",
 12633 => x"C0C0C0F9A482B0B0",
 12634 => x"C0C0C0F9A482B099",
 12635 => x"C0C0C0F9A482B092",
 12636 => x"C0C0C0F9A482B082",
 12637 => x"C0C0C0F9A482B0F8",
 12638 => x"C0C0C0F9A482B080",
 12639 => x"C0C0C0F9A482B090",
 12640 => x"C0C0C0F9A48299C0",
 12641 => x"C0C0C0F9A48299F9",
 12642 => x"C0C0C0F9A48299A4",
 12643 => x"C0C0C0F9A48299B0",
 12644 => x"C0C0C0F9A4829999",
 12645 => x"C0C0C0F9A4829992",
 12646 => x"C0C0C0F9A4829982",
 12647 => x"C0C0C0F9A48299F8",
 12648 => x"C0C0C0F9A4829980",
 12649 => x"C0C0C0F9A4829990",
 12650 => x"C0C0C0F9A48292C0",
 12651 => x"C0C0C0F9A48292F9",
 12652 => x"C0C0C0F9A48292A4",
 12653 => x"C0C0C0F9A48292B0",
 12654 => x"C0C0C0F9A4829299",
 12655 => x"C0C0C0F9A4829292",
 12656 => x"C0C0C0F9A4829282",
 12657 => x"C0C0C0F9A48292F8",
 12658 => x"C0C0C0F9A4829280",
 12659 => x"C0C0C0F9A4829290",
 12660 => x"C0C0C0F9A48282C0",
 12661 => x"C0C0C0F9A48282F9",
 12662 => x"C0C0C0F9A48282A4",
 12663 => x"C0C0C0F9A48282B0",
 12664 => x"C0C0C0F9A4828299",
 12665 => x"C0C0C0F9A4828292",
 12666 => x"C0C0C0F9A4828282",
 12667 => x"C0C0C0F9A48282F8",
 12668 => x"C0C0C0F9A4828280",
 12669 => x"C0C0C0F9A4828290",
 12670 => x"C0C0C0F9A482F8C0",
 12671 => x"C0C0C0F9A482F8F9",
 12672 => x"C0C0C0F9A482F8A4",
 12673 => x"C0C0C0F9A482F8B0",
 12674 => x"C0C0C0F9A482F899",
 12675 => x"C0C0C0F9A482F892",
 12676 => x"C0C0C0F9A482F882",
 12677 => x"C0C0C0F9A482F8F8",
 12678 => x"C0C0C0F9A482F880",
 12679 => x"C0C0C0F9A482F890",
 12680 => x"C0C0C0F9A48280C0",
 12681 => x"C0C0C0F9A48280F9",
 12682 => x"C0C0C0F9A48280A4",
 12683 => x"C0C0C0F9A48280B0",
 12684 => x"C0C0C0F9A4828099",
 12685 => x"C0C0C0F9A4828092",
 12686 => x"C0C0C0F9A4828082",
 12687 => x"C0C0C0F9A48280F8",
 12688 => x"C0C0C0F9A4828080",
 12689 => x"C0C0C0F9A4828090",
 12690 => x"C0C0C0F9A48290C0",
 12691 => x"C0C0C0F9A48290F9",
 12692 => x"C0C0C0F9A48290A4",
 12693 => x"C0C0C0F9A48290B0",
 12694 => x"C0C0C0F9A4829099",
 12695 => x"C0C0C0F9A4829092",
 12696 => x"C0C0C0F9A4829082",
 12697 => x"C0C0C0F9A48290F8",
 12698 => x"C0C0C0F9A4829080",
 12699 => x"C0C0C0F9A4829090",
 12700 => x"C0C0C0F9A4F8C0C0",
 12701 => x"C0C0C0F9A4F8C0F9",
 12702 => x"C0C0C0F9A4F8C0A4",
 12703 => x"C0C0C0F9A4F8C0B0",
 12704 => x"C0C0C0F9A4F8C099",
 12705 => x"C0C0C0F9A4F8C092",
 12706 => x"C0C0C0F9A4F8C082",
 12707 => x"C0C0C0F9A4F8C0F8",
 12708 => x"C0C0C0F9A4F8C080",
 12709 => x"C0C0C0F9A4F8C090",
 12710 => x"C0C0C0F9A4F8F9C0",
 12711 => x"C0C0C0F9A4F8F9F9",
 12712 => x"C0C0C0F9A4F8F9A4",
 12713 => x"C0C0C0F9A4F8F9B0",
 12714 => x"C0C0C0F9A4F8F999",
 12715 => x"C0C0C0F9A4F8F992",
 12716 => x"C0C0C0F9A4F8F982",
 12717 => x"C0C0C0F9A4F8F9F8",
 12718 => x"C0C0C0F9A4F8F980",
 12719 => x"C0C0C0F9A4F8F990",
 12720 => x"C0C0C0F9A4F8A4C0",
 12721 => x"C0C0C0F9A4F8A4F9",
 12722 => x"C0C0C0F9A4F8A4A4",
 12723 => x"C0C0C0F9A4F8A4B0",
 12724 => x"C0C0C0F9A4F8A499",
 12725 => x"C0C0C0F9A4F8A492",
 12726 => x"C0C0C0F9A4F8A482",
 12727 => x"C0C0C0F9A4F8A4F8",
 12728 => x"C0C0C0F9A4F8A480",
 12729 => x"C0C0C0F9A4F8A490",
 12730 => x"C0C0C0F9A4F8B0C0",
 12731 => x"C0C0C0F9A4F8B0F9",
 12732 => x"C0C0C0F9A4F8B0A4",
 12733 => x"C0C0C0F9A4F8B0B0",
 12734 => x"C0C0C0F9A4F8B099",
 12735 => x"C0C0C0F9A4F8B092",
 12736 => x"C0C0C0F9A4F8B082",
 12737 => x"C0C0C0F9A4F8B0F8",
 12738 => x"C0C0C0F9A4F8B080",
 12739 => x"C0C0C0F9A4F8B090",
 12740 => x"C0C0C0F9A4F899C0",
 12741 => x"C0C0C0F9A4F899F9",
 12742 => x"C0C0C0F9A4F899A4",
 12743 => x"C0C0C0F9A4F899B0",
 12744 => x"C0C0C0F9A4F89999",
 12745 => x"C0C0C0F9A4F89992",
 12746 => x"C0C0C0F9A4F89982",
 12747 => x"C0C0C0F9A4F899F8",
 12748 => x"C0C0C0F9A4F89980",
 12749 => x"C0C0C0F9A4F89990",
 12750 => x"C0C0C0F9A4F892C0",
 12751 => x"C0C0C0F9A4F892F9",
 12752 => x"C0C0C0F9A4F892A4",
 12753 => x"C0C0C0F9A4F892B0",
 12754 => x"C0C0C0F9A4F89299",
 12755 => x"C0C0C0F9A4F89292",
 12756 => x"C0C0C0F9A4F89282",
 12757 => x"C0C0C0F9A4F892F8",
 12758 => x"C0C0C0F9A4F89280",
 12759 => x"C0C0C0F9A4F89290",
 12760 => x"C0C0C0F9A4F882C0",
 12761 => x"C0C0C0F9A4F882F9",
 12762 => x"C0C0C0F9A4F882A4",
 12763 => x"C0C0C0F9A4F882B0",
 12764 => x"C0C0C0F9A4F88299",
 12765 => x"C0C0C0F9A4F88292",
 12766 => x"C0C0C0F9A4F88282",
 12767 => x"C0C0C0F9A4F882F8",
 12768 => x"C0C0C0F9A4F88280",
 12769 => x"C0C0C0F9A4F88290",
 12770 => x"C0C0C0F9A4F8F8C0",
 12771 => x"C0C0C0F9A4F8F8F9",
 12772 => x"C0C0C0F9A4F8F8A4",
 12773 => x"C0C0C0F9A4F8F8B0",
 12774 => x"C0C0C0F9A4F8F899",
 12775 => x"C0C0C0F9A4F8F892",
 12776 => x"C0C0C0F9A4F8F882",
 12777 => x"C0C0C0F9A4F8F8F8",
 12778 => x"C0C0C0F9A4F8F880",
 12779 => x"C0C0C0F9A4F8F890",
 12780 => x"C0C0C0F9A4F880C0",
 12781 => x"C0C0C0F9A4F880F9",
 12782 => x"C0C0C0F9A4F880A4",
 12783 => x"C0C0C0F9A4F880B0",
 12784 => x"C0C0C0F9A4F88099",
 12785 => x"C0C0C0F9A4F88092",
 12786 => x"C0C0C0F9A4F88082",
 12787 => x"C0C0C0F9A4F880F8",
 12788 => x"C0C0C0F9A4F88080",
 12789 => x"C0C0C0F9A4F88090",
 12790 => x"C0C0C0F9A4F890C0",
 12791 => x"C0C0C0F9A4F890F9",
 12792 => x"C0C0C0F9A4F890A4",
 12793 => x"C0C0C0F9A4F890B0",
 12794 => x"C0C0C0F9A4F89099",
 12795 => x"C0C0C0F9A4F89092",
 12796 => x"C0C0C0F9A4F89082",
 12797 => x"C0C0C0F9A4F890F8",
 12798 => x"C0C0C0F9A4F89080",
 12799 => x"C0C0C0F9A4F89090",
 12800 => x"C0C0C0F9A480C0C0",
 12801 => x"C0C0C0F9A480C0F9",
 12802 => x"C0C0C0F9A480C0A4",
 12803 => x"C0C0C0F9A480C0B0",
 12804 => x"C0C0C0F9A480C099",
 12805 => x"C0C0C0F9A480C092",
 12806 => x"C0C0C0F9A480C082",
 12807 => x"C0C0C0F9A480C0F8",
 12808 => x"C0C0C0F9A480C080",
 12809 => x"C0C0C0F9A480C090",
 12810 => x"C0C0C0F9A480F9C0",
 12811 => x"C0C0C0F9A480F9F9",
 12812 => x"C0C0C0F9A480F9A4",
 12813 => x"C0C0C0F9A480F9B0",
 12814 => x"C0C0C0F9A480F999",
 12815 => x"C0C0C0F9A480F992",
 12816 => x"C0C0C0F9A480F982",
 12817 => x"C0C0C0F9A480F9F8",
 12818 => x"C0C0C0F9A480F980",
 12819 => x"C0C0C0F9A480F990",
 12820 => x"C0C0C0F9A480A4C0",
 12821 => x"C0C0C0F9A480A4F9",
 12822 => x"C0C0C0F9A480A4A4",
 12823 => x"C0C0C0F9A480A4B0",
 12824 => x"C0C0C0F9A480A499",
 12825 => x"C0C0C0F9A480A492",
 12826 => x"C0C0C0F9A480A482",
 12827 => x"C0C0C0F9A480A4F8",
 12828 => x"C0C0C0F9A480A480",
 12829 => x"C0C0C0F9A480A490",
 12830 => x"C0C0C0F9A480B0C0",
 12831 => x"C0C0C0F9A480B0F9",
 12832 => x"C0C0C0F9A480B0A4",
 12833 => x"C0C0C0F9A480B0B0",
 12834 => x"C0C0C0F9A480B099",
 12835 => x"C0C0C0F9A480B092",
 12836 => x"C0C0C0F9A480B082",
 12837 => x"C0C0C0F9A480B0F8",
 12838 => x"C0C0C0F9A480B080",
 12839 => x"C0C0C0F9A480B090",
 12840 => x"C0C0C0F9A48099C0",
 12841 => x"C0C0C0F9A48099F9",
 12842 => x"C0C0C0F9A48099A4",
 12843 => x"C0C0C0F9A48099B0",
 12844 => x"C0C0C0F9A4809999",
 12845 => x"C0C0C0F9A4809992",
 12846 => x"C0C0C0F9A4809982",
 12847 => x"C0C0C0F9A48099F8",
 12848 => x"C0C0C0F9A4809980",
 12849 => x"C0C0C0F9A4809990",
 12850 => x"C0C0C0F9A48092C0",
 12851 => x"C0C0C0F9A48092F9",
 12852 => x"C0C0C0F9A48092A4",
 12853 => x"C0C0C0F9A48092B0",
 12854 => x"C0C0C0F9A4809299",
 12855 => x"C0C0C0F9A4809292",
 12856 => x"C0C0C0F9A4809282",
 12857 => x"C0C0C0F9A48092F8",
 12858 => x"C0C0C0F9A4809280",
 12859 => x"C0C0C0F9A4809290",
 12860 => x"C0C0C0F9A48082C0",
 12861 => x"C0C0C0F9A48082F9",
 12862 => x"C0C0C0F9A48082A4",
 12863 => x"C0C0C0F9A48082B0",
 12864 => x"C0C0C0F9A4808299",
 12865 => x"C0C0C0F9A4808292",
 12866 => x"C0C0C0F9A4808282",
 12867 => x"C0C0C0F9A48082F8",
 12868 => x"C0C0C0F9A4808280",
 12869 => x"C0C0C0F9A4808290",
 12870 => x"C0C0C0F9A480F8C0",
 12871 => x"C0C0C0F9A480F8F9",
 12872 => x"C0C0C0F9A480F8A4",
 12873 => x"C0C0C0F9A480F8B0",
 12874 => x"C0C0C0F9A480F899",
 12875 => x"C0C0C0F9A480F892",
 12876 => x"C0C0C0F9A480F882",
 12877 => x"C0C0C0F9A480F8F8",
 12878 => x"C0C0C0F9A480F880",
 12879 => x"C0C0C0F9A480F890",
 12880 => x"C0C0C0F9A48080C0",
 12881 => x"C0C0C0F9A48080F9",
 12882 => x"C0C0C0F9A48080A4",
 12883 => x"C0C0C0F9A48080B0",
 12884 => x"C0C0C0F9A4808099",
 12885 => x"C0C0C0F9A4808092",
 12886 => x"C0C0C0F9A4808082",
 12887 => x"C0C0C0F9A48080F8",
 12888 => x"C0C0C0F9A4808080",
 12889 => x"C0C0C0F9A4808090",
 12890 => x"C0C0C0F9A48090C0",
 12891 => x"C0C0C0F9A48090F9",
 12892 => x"C0C0C0F9A48090A4",
 12893 => x"C0C0C0F9A48090B0",
 12894 => x"C0C0C0F9A4809099",
 12895 => x"C0C0C0F9A4809092",
 12896 => x"C0C0C0F9A4809082",
 12897 => x"C0C0C0F9A48090F8",
 12898 => x"C0C0C0F9A4809080",
 12899 => x"C0C0C0F9A4809090",
 12900 => x"C0C0C0F9A490C0C0",
 12901 => x"C0C0C0F9A490C0F9",
 12902 => x"C0C0C0F9A490C0A4",
 12903 => x"C0C0C0F9A490C0B0",
 12904 => x"C0C0C0F9A490C099",
 12905 => x"C0C0C0F9A490C092",
 12906 => x"C0C0C0F9A490C082",
 12907 => x"C0C0C0F9A490C0F8",
 12908 => x"C0C0C0F9A490C080",
 12909 => x"C0C0C0F9A490C090",
 12910 => x"C0C0C0F9A490F9C0",
 12911 => x"C0C0C0F9A490F9F9",
 12912 => x"C0C0C0F9A490F9A4",
 12913 => x"C0C0C0F9A490F9B0",
 12914 => x"C0C0C0F9A490F999",
 12915 => x"C0C0C0F9A490F992",
 12916 => x"C0C0C0F9A490F982",
 12917 => x"C0C0C0F9A490F9F8",
 12918 => x"C0C0C0F9A490F980",
 12919 => x"C0C0C0F9A490F990",
 12920 => x"C0C0C0F9A490A4C0",
 12921 => x"C0C0C0F9A490A4F9",
 12922 => x"C0C0C0F9A490A4A4",
 12923 => x"C0C0C0F9A490A4B0",
 12924 => x"C0C0C0F9A490A499",
 12925 => x"C0C0C0F9A490A492",
 12926 => x"C0C0C0F9A490A482",
 12927 => x"C0C0C0F9A490A4F8",
 12928 => x"C0C0C0F9A490A480",
 12929 => x"C0C0C0F9A490A490",
 12930 => x"C0C0C0F9A490B0C0",
 12931 => x"C0C0C0F9A490B0F9",
 12932 => x"C0C0C0F9A490B0A4",
 12933 => x"C0C0C0F9A490B0B0",
 12934 => x"C0C0C0F9A490B099",
 12935 => x"C0C0C0F9A490B092",
 12936 => x"C0C0C0F9A490B082",
 12937 => x"C0C0C0F9A490B0F8",
 12938 => x"C0C0C0F9A490B080",
 12939 => x"C0C0C0F9A490B090",
 12940 => x"C0C0C0F9A49099C0",
 12941 => x"C0C0C0F9A49099F9",
 12942 => x"C0C0C0F9A49099A4",
 12943 => x"C0C0C0F9A49099B0",
 12944 => x"C0C0C0F9A4909999",
 12945 => x"C0C0C0F9A4909992",
 12946 => x"C0C0C0F9A4909982",
 12947 => x"C0C0C0F9A49099F8",
 12948 => x"C0C0C0F9A4909980",
 12949 => x"C0C0C0F9A4909990",
 12950 => x"C0C0C0F9A49092C0",
 12951 => x"C0C0C0F9A49092F9",
 12952 => x"C0C0C0F9A49092A4",
 12953 => x"C0C0C0F9A49092B0",
 12954 => x"C0C0C0F9A4909299",
 12955 => x"C0C0C0F9A4909292",
 12956 => x"C0C0C0F9A4909282",
 12957 => x"C0C0C0F9A49092F8",
 12958 => x"C0C0C0F9A4909280",
 12959 => x"C0C0C0F9A4909290",
 12960 => x"C0C0C0F9A49082C0",
 12961 => x"C0C0C0F9A49082F9",
 12962 => x"C0C0C0F9A49082A4",
 12963 => x"C0C0C0F9A49082B0",
 12964 => x"C0C0C0F9A4908299",
 12965 => x"C0C0C0F9A4908292",
 12966 => x"C0C0C0F9A4908282",
 12967 => x"C0C0C0F9A49082F8",
 12968 => x"C0C0C0F9A4908280",
 12969 => x"C0C0C0F9A4908290",
 12970 => x"C0C0C0F9A490F8C0",
 12971 => x"C0C0C0F9A490F8F9",
 12972 => x"C0C0C0F9A490F8A4",
 12973 => x"C0C0C0F9A490F8B0",
 12974 => x"C0C0C0F9A490F899",
 12975 => x"C0C0C0F9A490F892",
 12976 => x"C0C0C0F9A490F882",
 12977 => x"C0C0C0F9A490F8F8",
 12978 => x"C0C0C0F9A490F880",
 12979 => x"C0C0C0F9A490F890",
 12980 => x"C0C0C0F9A49080C0",
 12981 => x"C0C0C0F9A49080F9",
 12982 => x"C0C0C0F9A49080A4",
 12983 => x"C0C0C0F9A49080B0",
 12984 => x"C0C0C0F9A4908099",
 12985 => x"C0C0C0F9A4908092",
 12986 => x"C0C0C0F9A4908082",
 12987 => x"C0C0C0F9A49080F8",
 12988 => x"C0C0C0F9A4908080",
 12989 => x"C0C0C0F9A4908090",
 12990 => x"C0C0C0F9A49090C0",
 12991 => x"C0C0C0F9A49090F9",
 12992 => x"C0C0C0F9A49090A4",
 12993 => x"C0C0C0F9A49090B0",
 12994 => x"C0C0C0F9A4909099",
 12995 => x"C0C0C0F9A4909092",
 12996 => x"C0C0C0F9A4909082",
 12997 => x"C0C0C0F9A49090F8",
 12998 => x"C0C0C0F9A4909080",
 12999 => x"C0C0C0F9A4909090",
 13000 => x"C0C0C0F9B0C0C0C0",
 13001 => x"C0C0C0F9B0C0C0F9",
 13002 => x"C0C0C0F9B0C0C0A4",
 13003 => x"C0C0C0F9B0C0C0B0",
 13004 => x"C0C0C0F9B0C0C099",
 13005 => x"C0C0C0F9B0C0C092",
 13006 => x"C0C0C0F9B0C0C082",
 13007 => x"C0C0C0F9B0C0C0F8",
 13008 => x"C0C0C0F9B0C0C080",
 13009 => x"C0C0C0F9B0C0C090",
 13010 => x"C0C0C0F9B0C0F9C0",
 13011 => x"C0C0C0F9B0C0F9F9",
 13012 => x"C0C0C0F9B0C0F9A4",
 13013 => x"C0C0C0F9B0C0F9B0",
 13014 => x"C0C0C0F9B0C0F999",
 13015 => x"C0C0C0F9B0C0F992",
 13016 => x"C0C0C0F9B0C0F982",
 13017 => x"C0C0C0F9B0C0F9F8",
 13018 => x"C0C0C0F9B0C0F980",
 13019 => x"C0C0C0F9B0C0F990",
 13020 => x"C0C0C0F9B0C0A4C0",
 13021 => x"C0C0C0F9B0C0A4F9",
 13022 => x"C0C0C0F9B0C0A4A4",
 13023 => x"C0C0C0F9B0C0A4B0",
 13024 => x"C0C0C0F9B0C0A499",
 13025 => x"C0C0C0F9B0C0A492",
 13026 => x"C0C0C0F9B0C0A482",
 13027 => x"C0C0C0F9B0C0A4F8",
 13028 => x"C0C0C0F9B0C0A480",
 13029 => x"C0C0C0F9B0C0A490",
 13030 => x"C0C0C0F9B0C0B0C0",
 13031 => x"C0C0C0F9B0C0B0F9",
 13032 => x"C0C0C0F9B0C0B0A4",
 13033 => x"C0C0C0F9B0C0B0B0",
 13034 => x"C0C0C0F9B0C0B099",
 13035 => x"C0C0C0F9B0C0B092",
 13036 => x"C0C0C0F9B0C0B082",
 13037 => x"C0C0C0F9B0C0B0F8",
 13038 => x"C0C0C0F9B0C0B080",
 13039 => x"C0C0C0F9B0C0B090",
 13040 => x"C0C0C0F9B0C099C0",
 13041 => x"C0C0C0F9B0C099F9",
 13042 => x"C0C0C0F9B0C099A4",
 13043 => x"C0C0C0F9B0C099B0",
 13044 => x"C0C0C0F9B0C09999",
 13045 => x"C0C0C0F9B0C09992",
 13046 => x"C0C0C0F9B0C09982",
 13047 => x"C0C0C0F9B0C099F8",
 13048 => x"C0C0C0F9B0C09980",
 13049 => x"C0C0C0F9B0C09990",
 13050 => x"C0C0C0F9B0C092C0",
 13051 => x"C0C0C0F9B0C092F9",
 13052 => x"C0C0C0F9B0C092A4",
 13053 => x"C0C0C0F9B0C092B0",
 13054 => x"C0C0C0F9B0C09299",
 13055 => x"C0C0C0F9B0C09292",
 13056 => x"C0C0C0F9B0C09282",
 13057 => x"C0C0C0F9B0C092F8",
 13058 => x"C0C0C0F9B0C09280",
 13059 => x"C0C0C0F9B0C09290",
 13060 => x"C0C0C0F9B0C082C0",
 13061 => x"C0C0C0F9B0C082F9",
 13062 => x"C0C0C0F9B0C082A4",
 13063 => x"C0C0C0F9B0C082B0",
 13064 => x"C0C0C0F9B0C08299",
 13065 => x"C0C0C0F9B0C08292",
 13066 => x"C0C0C0F9B0C08282",
 13067 => x"C0C0C0F9B0C082F8",
 13068 => x"C0C0C0F9B0C08280",
 13069 => x"C0C0C0F9B0C08290",
 13070 => x"C0C0C0F9B0C0F8C0",
 13071 => x"C0C0C0F9B0C0F8F9",
 13072 => x"C0C0C0F9B0C0F8A4",
 13073 => x"C0C0C0F9B0C0F8B0",
 13074 => x"C0C0C0F9B0C0F899",
 13075 => x"C0C0C0F9B0C0F892",
 13076 => x"C0C0C0F9B0C0F882",
 13077 => x"C0C0C0F9B0C0F8F8",
 13078 => x"C0C0C0F9B0C0F880",
 13079 => x"C0C0C0F9B0C0F890",
 13080 => x"C0C0C0F9B0C080C0",
 13081 => x"C0C0C0F9B0C080F9",
 13082 => x"C0C0C0F9B0C080A4",
 13083 => x"C0C0C0F9B0C080B0",
 13084 => x"C0C0C0F9B0C08099",
 13085 => x"C0C0C0F9B0C08092",
 13086 => x"C0C0C0F9B0C08082",
 13087 => x"C0C0C0F9B0C080F8",
 13088 => x"C0C0C0F9B0C08080",
 13089 => x"C0C0C0F9B0C08090",
 13090 => x"C0C0C0F9B0C090C0",
 13091 => x"C0C0C0F9B0C090F9",
 13092 => x"C0C0C0F9B0C090A4",
 13093 => x"C0C0C0F9B0C090B0",
 13094 => x"C0C0C0F9B0C09099",
 13095 => x"C0C0C0F9B0C09092",
 13096 => x"C0C0C0F9B0C09082",
 13097 => x"C0C0C0F9B0C090F8",
 13098 => x"C0C0C0F9B0C09080",
 13099 => x"C0C0C0F9B0C09090",
 13100 => x"C0C0C0F9B0F9C0C0",
 13101 => x"C0C0C0F9B0F9C0F9",
 13102 => x"C0C0C0F9B0F9C0A4",
 13103 => x"C0C0C0F9B0F9C0B0",
 13104 => x"C0C0C0F9B0F9C099",
 13105 => x"C0C0C0F9B0F9C092",
 13106 => x"C0C0C0F9B0F9C082",
 13107 => x"C0C0C0F9B0F9C0F8",
 13108 => x"C0C0C0F9B0F9C080",
 13109 => x"C0C0C0F9B0F9C090",
 13110 => x"C0C0C0F9B0F9F9C0",
 13111 => x"C0C0C0F9B0F9F9F9",
 13112 => x"C0C0C0F9B0F9F9A4",
 13113 => x"C0C0C0F9B0F9F9B0",
 13114 => x"C0C0C0F9B0F9F999",
 13115 => x"C0C0C0F9B0F9F992",
 13116 => x"C0C0C0F9B0F9F982",
 13117 => x"C0C0C0F9B0F9F9F8",
 13118 => x"C0C0C0F9B0F9F980",
 13119 => x"C0C0C0F9B0F9F990",
 13120 => x"C0C0C0F9B0F9A4C0",
 13121 => x"C0C0C0F9B0F9A4F9",
 13122 => x"C0C0C0F9B0F9A4A4",
 13123 => x"C0C0C0F9B0F9A4B0",
 13124 => x"C0C0C0F9B0F9A499",
 13125 => x"C0C0C0F9B0F9A492",
 13126 => x"C0C0C0F9B0F9A482",
 13127 => x"C0C0C0F9B0F9A4F8",
 13128 => x"C0C0C0F9B0F9A480",
 13129 => x"C0C0C0F9B0F9A490",
 13130 => x"C0C0C0F9B0F9B0C0",
 13131 => x"C0C0C0F9B0F9B0F9",
 13132 => x"C0C0C0F9B0F9B0A4",
 13133 => x"C0C0C0F9B0F9B0B0",
 13134 => x"C0C0C0F9B0F9B099",
 13135 => x"C0C0C0F9B0F9B092",
 13136 => x"C0C0C0F9B0F9B082",
 13137 => x"C0C0C0F9B0F9B0F8",
 13138 => x"C0C0C0F9B0F9B080",
 13139 => x"C0C0C0F9B0F9B090",
 13140 => x"C0C0C0F9B0F999C0",
 13141 => x"C0C0C0F9B0F999F9",
 13142 => x"C0C0C0F9B0F999A4",
 13143 => x"C0C0C0F9B0F999B0",
 13144 => x"C0C0C0F9B0F99999",
 13145 => x"C0C0C0F9B0F99992",
 13146 => x"C0C0C0F9B0F99982",
 13147 => x"C0C0C0F9B0F999F8",
 13148 => x"C0C0C0F9B0F99980",
 13149 => x"C0C0C0F9B0F99990",
 13150 => x"C0C0C0F9B0F992C0",
 13151 => x"C0C0C0F9B0F992F9",
 13152 => x"C0C0C0F9B0F992A4",
 13153 => x"C0C0C0F9B0F992B0",
 13154 => x"C0C0C0F9B0F99299",
 13155 => x"C0C0C0F9B0F99292",
 13156 => x"C0C0C0F9B0F99282",
 13157 => x"C0C0C0F9B0F992F8",
 13158 => x"C0C0C0F9B0F99280",
 13159 => x"C0C0C0F9B0F99290",
 13160 => x"C0C0C0F9B0F982C0",
 13161 => x"C0C0C0F9B0F982F9",
 13162 => x"C0C0C0F9B0F982A4",
 13163 => x"C0C0C0F9B0F982B0",
 13164 => x"C0C0C0F9B0F98299",
 13165 => x"C0C0C0F9B0F98292",
 13166 => x"C0C0C0F9B0F98282",
 13167 => x"C0C0C0F9B0F982F8",
 13168 => x"C0C0C0F9B0F98280",
 13169 => x"C0C0C0F9B0F98290",
 13170 => x"C0C0C0F9B0F9F8C0",
 13171 => x"C0C0C0F9B0F9F8F9",
 13172 => x"C0C0C0F9B0F9F8A4",
 13173 => x"C0C0C0F9B0F9F8B0",
 13174 => x"C0C0C0F9B0F9F899",
 13175 => x"C0C0C0F9B0F9F892",
 13176 => x"C0C0C0F9B0F9F882",
 13177 => x"C0C0C0F9B0F9F8F8",
 13178 => x"C0C0C0F9B0F9F880",
 13179 => x"C0C0C0F9B0F9F890",
 13180 => x"C0C0C0F9B0F980C0",
 13181 => x"C0C0C0F9B0F980F9",
 13182 => x"C0C0C0F9B0F980A4",
 13183 => x"C0C0C0F9B0F980B0",
 13184 => x"C0C0C0F9B0F98099",
 13185 => x"C0C0C0F9B0F98092",
 13186 => x"C0C0C0F9B0F98082",
 13187 => x"C0C0C0F9B0F980F8",
 13188 => x"C0C0C0F9B0F98080",
 13189 => x"C0C0C0F9B0F98090",
 13190 => x"C0C0C0F9B0F990C0",
 13191 => x"C0C0C0F9B0F990F9",
 13192 => x"C0C0C0F9B0F990A4",
 13193 => x"C0C0C0F9B0F990B0",
 13194 => x"C0C0C0F9B0F99099",
 13195 => x"C0C0C0F9B0F99092",
 13196 => x"C0C0C0F9B0F99082",
 13197 => x"C0C0C0F9B0F990F8",
 13198 => x"C0C0C0F9B0F99080",
 13199 => x"C0C0C0F9B0F99090",
 13200 => x"C0C0C0F9B0A4C0C0",
 13201 => x"C0C0C0F9B0A4C0F9",
 13202 => x"C0C0C0F9B0A4C0A4",
 13203 => x"C0C0C0F9B0A4C0B0",
 13204 => x"C0C0C0F9B0A4C099",
 13205 => x"C0C0C0F9B0A4C092",
 13206 => x"C0C0C0F9B0A4C082",
 13207 => x"C0C0C0F9B0A4C0F8",
 13208 => x"C0C0C0F9B0A4C080",
 13209 => x"C0C0C0F9B0A4C090",
 13210 => x"C0C0C0F9B0A4F9C0",
 13211 => x"C0C0C0F9B0A4F9F9",
 13212 => x"C0C0C0F9B0A4F9A4",
 13213 => x"C0C0C0F9B0A4F9B0",
 13214 => x"C0C0C0F9B0A4F999",
 13215 => x"C0C0C0F9B0A4F992",
 13216 => x"C0C0C0F9B0A4F982",
 13217 => x"C0C0C0F9B0A4F9F8",
 13218 => x"C0C0C0F9B0A4F980",
 13219 => x"C0C0C0F9B0A4F990",
 13220 => x"C0C0C0F9B0A4A4C0",
 13221 => x"C0C0C0F9B0A4A4F9",
 13222 => x"C0C0C0F9B0A4A4A4",
 13223 => x"C0C0C0F9B0A4A4B0",
 13224 => x"C0C0C0F9B0A4A499",
 13225 => x"C0C0C0F9B0A4A492",
 13226 => x"C0C0C0F9B0A4A482",
 13227 => x"C0C0C0F9B0A4A4F8",
 13228 => x"C0C0C0F9B0A4A480",
 13229 => x"C0C0C0F9B0A4A490",
 13230 => x"C0C0C0F9B0A4B0C0",
 13231 => x"C0C0C0F9B0A4B0F9",
 13232 => x"C0C0C0F9B0A4B0A4",
 13233 => x"C0C0C0F9B0A4B0B0",
 13234 => x"C0C0C0F9B0A4B099",
 13235 => x"C0C0C0F9B0A4B092",
 13236 => x"C0C0C0F9B0A4B082",
 13237 => x"C0C0C0F9B0A4B0F8",
 13238 => x"C0C0C0F9B0A4B080",
 13239 => x"C0C0C0F9B0A4B090",
 13240 => x"C0C0C0F9B0A499C0",
 13241 => x"C0C0C0F9B0A499F9",
 13242 => x"C0C0C0F9B0A499A4",
 13243 => x"C0C0C0F9B0A499B0",
 13244 => x"C0C0C0F9B0A49999",
 13245 => x"C0C0C0F9B0A49992",
 13246 => x"C0C0C0F9B0A49982",
 13247 => x"C0C0C0F9B0A499F8",
 13248 => x"C0C0C0F9B0A49980",
 13249 => x"C0C0C0F9B0A49990",
 13250 => x"C0C0C0F9B0A492C0",
 13251 => x"C0C0C0F9B0A492F9",
 13252 => x"C0C0C0F9B0A492A4",
 13253 => x"C0C0C0F9B0A492B0",
 13254 => x"C0C0C0F9B0A49299",
 13255 => x"C0C0C0F9B0A49292",
 13256 => x"C0C0C0F9B0A49282",
 13257 => x"C0C0C0F9B0A492F8",
 13258 => x"C0C0C0F9B0A49280",
 13259 => x"C0C0C0F9B0A49290",
 13260 => x"C0C0C0F9B0A482C0",
 13261 => x"C0C0C0F9B0A482F9",
 13262 => x"C0C0C0F9B0A482A4",
 13263 => x"C0C0C0F9B0A482B0",
 13264 => x"C0C0C0F9B0A48299",
 13265 => x"C0C0C0F9B0A48292",
 13266 => x"C0C0C0F9B0A48282",
 13267 => x"C0C0C0F9B0A482F8",
 13268 => x"C0C0C0F9B0A48280",
 13269 => x"C0C0C0F9B0A48290",
 13270 => x"C0C0C0F9B0A4F8C0",
 13271 => x"C0C0C0F9B0A4F8F9",
 13272 => x"C0C0C0F9B0A4F8A4",
 13273 => x"C0C0C0F9B0A4F8B0",
 13274 => x"C0C0C0F9B0A4F899",
 13275 => x"C0C0C0F9B0A4F892",
 13276 => x"C0C0C0F9B0A4F882",
 13277 => x"C0C0C0F9B0A4F8F8",
 13278 => x"C0C0C0F9B0A4F880",
 13279 => x"C0C0C0F9B0A4F890",
 13280 => x"C0C0C0F9B0A480C0",
 13281 => x"C0C0C0F9B0A480F9",
 13282 => x"C0C0C0F9B0A480A4",
 13283 => x"C0C0C0F9B0A480B0",
 13284 => x"C0C0C0F9B0A48099",
 13285 => x"C0C0C0F9B0A48092",
 13286 => x"C0C0C0F9B0A48082",
 13287 => x"C0C0C0F9B0A480F8",
 13288 => x"C0C0C0F9B0A48080",
 13289 => x"C0C0C0F9B0A48090",
 13290 => x"C0C0C0F9B0A490C0",
 13291 => x"C0C0C0F9B0A490F9",
 13292 => x"C0C0C0F9B0A490A4",
 13293 => x"C0C0C0F9B0A490B0",
 13294 => x"C0C0C0F9B0A49099",
 13295 => x"C0C0C0F9B0A49092",
 13296 => x"C0C0C0F9B0A49082",
 13297 => x"C0C0C0F9B0A490F8",
 13298 => x"C0C0C0F9B0A49080",
 13299 => x"C0C0C0F9B0A49090",
 13300 => x"C0C0C0F9B0B0C0C0",
 13301 => x"C0C0C0F9B0B0C0F9",
 13302 => x"C0C0C0F9B0B0C0A4",
 13303 => x"C0C0C0F9B0B0C0B0",
 13304 => x"C0C0C0F9B0B0C099",
 13305 => x"C0C0C0F9B0B0C092",
 13306 => x"C0C0C0F9B0B0C082",
 13307 => x"C0C0C0F9B0B0C0F8",
 13308 => x"C0C0C0F9B0B0C080",
 13309 => x"C0C0C0F9B0B0C090",
 13310 => x"C0C0C0F9B0B0F9C0",
 13311 => x"C0C0C0F9B0B0F9F9",
 13312 => x"C0C0C0F9B0B0F9A4",
 13313 => x"C0C0C0F9B0B0F9B0",
 13314 => x"C0C0C0F9B0B0F999",
 13315 => x"C0C0C0F9B0B0F992",
 13316 => x"C0C0C0F9B0B0F982",
 13317 => x"C0C0C0F9B0B0F9F8",
 13318 => x"C0C0C0F9B0B0F980",
 13319 => x"C0C0C0F9B0B0F990",
 13320 => x"C0C0C0F9B0B0A4C0",
 13321 => x"C0C0C0F9B0B0A4F9",
 13322 => x"C0C0C0F9B0B0A4A4",
 13323 => x"C0C0C0F9B0B0A4B0",
 13324 => x"C0C0C0F9B0B0A499",
 13325 => x"C0C0C0F9B0B0A492",
 13326 => x"C0C0C0F9B0B0A482",
 13327 => x"C0C0C0F9B0B0A4F8",
 13328 => x"C0C0C0F9B0B0A480",
 13329 => x"C0C0C0F9B0B0A490",
 13330 => x"C0C0C0F9B0B0B0C0",
 13331 => x"C0C0C0F9B0B0B0F9",
 13332 => x"C0C0C0F9B0B0B0A4",
 13333 => x"C0C0C0F9B0B0B0B0",
 13334 => x"C0C0C0F9B0B0B099",
 13335 => x"C0C0C0F9B0B0B092",
 13336 => x"C0C0C0F9B0B0B082",
 13337 => x"C0C0C0F9B0B0B0F8",
 13338 => x"C0C0C0F9B0B0B080",
 13339 => x"C0C0C0F9B0B0B090",
 13340 => x"C0C0C0F9B0B099C0",
 13341 => x"C0C0C0F9B0B099F9",
 13342 => x"C0C0C0F9B0B099A4",
 13343 => x"C0C0C0F9B0B099B0",
 13344 => x"C0C0C0F9B0B09999",
 13345 => x"C0C0C0F9B0B09992",
 13346 => x"C0C0C0F9B0B09982",
 13347 => x"C0C0C0F9B0B099F8",
 13348 => x"C0C0C0F9B0B09980",
 13349 => x"C0C0C0F9B0B09990",
 13350 => x"C0C0C0F9B0B092C0",
 13351 => x"C0C0C0F9B0B092F9",
 13352 => x"C0C0C0F9B0B092A4",
 13353 => x"C0C0C0F9B0B092B0",
 13354 => x"C0C0C0F9B0B09299",
 13355 => x"C0C0C0F9B0B09292",
 13356 => x"C0C0C0F9B0B09282",
 13357 => x"C0C0C0F9B0B092F8",
 13358 => x"C0C0C0F9B0B09280",
 13359 => x"C0C0C0F9B0B09290",
 13360 => x"C0C0C0F9B0B082C0",
 13361 => x"C0C0C0F9B0B082F9",
 13362 => x"C0C0C0F9B0B082A4",
 13363 => x"C0C0C0F9B0B082B0",
 13364 => x"C0C0C0F9B0B08299",
 13365 => x"C0C0C0F9B0B08292",
 13366 => x"C0C0C0F9B0B08282",
 13367 => x"C0C0C0F9B0B082F8",
 13368 => x"C0C0C0F9B0B08280",
 13369 => x"C0C0C0F9B0B08290",
 13370 => x"C0C0C0F9B0B0F8C0",
 13371 => x"C0C0C0F9B0B0F8F9",
 13372 => x"C0C0C0F9B0B0F8A4",
 13373 => x"C0C0C0F9B0B0F8B0",
 13374 => x"C0C0C0F9B0B0F899",
 13375 => x"C0C0C0F9B0B0F892",
 13376 => x"C0C0C0F9B0B0F882",
 13377 => x"C0C0C0F9B0B0F8F8",
 13378 => x"C0C0C0F9B0B0F880",
 13379 => x"C0C0C0F9B0B0F890",
 13380 => x"C0C0C0F9B0B080C0",
 13381 => x"C0C0C0F9B0B080F9",
 13382 => x"C0C0C0F9B0B080A4",
 13383 => x"C0C0C0F9B0B080B0",
 13384 => x"C0C0C0F9B0B08099",
 13385 => x"C0C0C0F9B0B08092",
 13386 => x"C0C0C0F9B0B08082",
 13387 => x"C0C0C0F9B0B080F8",
 13388 => x"C0C0C0F9B0B08080",
 13389 => x"C0C0C0F9B0B08090",
 13390 => x"C0C0C0F9B0B090C0",
 13391 => x"C0C0C0F9B0B090F9",
 13392 => x"C0C0C0F9B0B090A4",
 13393 => x"C0C0C0F9B0B090B0",
 13394 => x"C0C0C0F9B0B09099",
 13395 => x"C0C0C0F9B0B09092",
 13396 => x"C0C0C0F9B0B09082",
 13397 => x"C0C0C0F9B0B090F8",
 13398 => x"C0C0C0F9B0B09080",
 13399 => x"C0C0C0F9B0B09090",
 13400 => x"C0C0C0F9B099C0C0",
 13401 => x"C0C0C0F9B099C0F9",
 13402 => x"C0C0C0F9B099C0A4",
 13403 => x"C0C0C0F9B099C0B0",
 13404 => x"C0C0C0F9B099C099",
 13405 => x"C0C0C0F9B099C092",
 13406 => x"C0C0C0F9B099C082",
 13407 => x"C0C0C0F9B099C0F8",
 13408 => x"C0C0C0F9B099C080",
 13409 => x"C0C0C0F9B099C090",
 13410 => x"C0C0C0F9B099F9C0",
 13411 => x"C0C0C0F9B099F9F9",
 13412 => x"C0C0C0F9B099F9A4",
 13413 => x"C0C0C0F9B099F9B0",
 13414 => x"C0C0C0F9B099F999",
 13415 => x"C0C0C0F9B099F992",
 13416 => x"C0C0C0F9B099F982",
 13417 => x"C0C0C0F9B099F9F8",
 13418 => x"C0C0C0F9B099F980",
 13419 => x"C0C0C0F9B099F990",
 13420 => x"C0C0C0F9B099A4C0",
 13421 => x"C0C0C0F9B099A4F9",
 13422 => x"C0C0C0F9B099A4A4",
 13423 => x"C0C0C0F9B099A4B0",
 13424 => x"C0C0C0F9B099A499",
 13425 => x"C0C0C0F9B099A492",
 13426 => x"C0C0C0F9B099A482",
 13427 => x"C0C0C0F9B099A4F8",
 13428 => x"C0C0C0F9B099A480",
 13429 => x"C0C0C0F9B099A490",
 13430 => x"C0C0C0F9B099B0C0",
 13431 => x"C0C0C0F9B099B0F9",
 13432 => x"C0C0C0F9B099B0A4",
 13433 => x"C0C0C0F9B099B0B0",
 13434 => x"C0C0C0F9B099B099",
 13435 => x"C0C0C0F9B099B092",
 13436 => x"C0C0C0F9B099B082",
 13437 => x"C0C0C0F9B099B0F8",
 13438 => x"C0C0C0F9B099B080",
 13439 => x"C0C0C0F9B099B090",
 13440 => x"C0C0C0F9B09999C0",
 13441 => x"C0C0C0F9B09999F9",
 13442 => x"C0C0C0F9B09999A4",
 13443 => x"C0C0C0F9B09999B0",
 13444 => x"C0C0C0F9B0999999",
 13445 => x"C0C0C0F9B0999992",
 13446 => x"C0C0C0F9B0999982",
 13447 => x"C0C0C0F9B09999F8",
 13448 => x"C0C0C0F9B0999980",
 13449 => x"C0C0C0F9B0999990",
 13450 => x"C0C0C0F9B09992C0",
 13451 => x"C0C0C0F9B09992F9",
 13452 => x"C0C0C0F9B09992A4",
 13453 => x"C0C0C0F9B09992B0",
 13454 => x"C0C0C0F9B0999299",
 13455 => x"C0C0C0F9B0999292",
 13456 => x"C0C0C0F9B0999282",
 13457 => x"C0C0C0F9B09992F8",
 13458 => x"C0C0C0F9B0999280",
 13459 => x"C0C0C0F9B0999290",
 13460 => x"C0C0C0F9B09982C0",
 13461 => x"C0C0C0F9B09982F9",
 13462 => x"C0C0C0F9B09982A4",
 13463 => x"C0C0C0F9B09982B0",
 13464 => x"C0C0C0F9B0998299",
 13465 => x"C0C0C0F9B0998292",
 13466 => x"C0C0C0F9B0998282",
 13467 => x"C0C0C0F9B09982F8",
 13468 => x"C0C0C0F9B0998280",
 13469 => x"C0C0C0F9B0998290",
 13470 => x"C0C0C0F9B099F8C0",
 13471 => x"C0C0C0F9B099F8F9",
 13472 => x"C0C0C0F9B099F8A4",
 13473 => x"C0C0C0F9B099F8B0",
 13474 => x"C0C0C0F9B099F899",
 13475 => x"C0C0C0F9B099F892",
 13476 => x"C0C0C0F9B099F882",
 13477 => x"C0C0C0F9B099F8F8",
 13478 => x"C0C0C0F9B099F880",
 13479 => x"C0C0C0F9B099F890",
 13480 => x"C0C0C0F9B09980C0",
 13481 => x"C0C0C0F9B09980F9",
 13482 => x"C0C0C0F9B09980A4",
 13483 => x"C0C0C0F9B09980B0",
 13484 => x"C0C0C0F9B0998099",
 13485 => x"C0C0C0F9B0998092",
 13486 => x"C0C0C0F9B0998082",
 13487 => x"C0C0C0F9B09980F8",
 13488 => x"C0C0C0F9B0998080",
 13489 => x"C0C0C0F9B0998090",
 13490 => x"C0C0C0F9B09990C0",
 13491 => x"C0C0C0F9B09990F9",
 13492 => x"C0C0C0F9B09990A4",
 13493 => x"C0C0C0F9B09990B0",
 13494 => x"C0C0C0F9B0999099",
 13495 => x"C0C0C0F9B0999092",
 13496 => x"C0C0C0F9B0999082",
 13497 => x"C0C0C0F9B09990F8",
 13498 => x"C0C0C0F9B0999080",
 13499 => x"C0C0C0F9B0999090",
 13500 => x"C0C0C0F9B092C0C0",
 13501 => x"C0C0C0F9B092C0F9",
 13502 => x"C0C0C0F9B092C0A4",
 13503 => x"C0C0C0F9B092C0B0",
 13504 => x"C0C0C0F9B092C099",
 13505 => x"C0C0C0F9B092C092",
 13506 => x"C0C0C0F9B092C082",
 13507 => x"C0C0C0F9B092C0F8",
 13508 => x"C0C0C0F9B092C080",
 13509 => x"C0C0C0F9B092C090",
 13510 => x"C0C0C0F9B092F9C0",
 13511 => x"C0C0C0F9B092F9F9",
 13512 => x"C0C0C0F9B092F9A4",
 13513 => x"C0C0C0F9B092F9B0",
 13514 => x"C0C0C0F9B092F999",
 13515 => x"C0C0C0F9B092F992",
 13516 => x"C0C0C0F9B092F982",
 13517 => x"C0C0C0F9B092F9F8",
 13518 => x"C0C0C0F9B092F980",
 13519 => x"C0C0C0F9B092F990",
 13520 => x"C0C0C0F9B092A4C0",
 13521 => x"C0C0C0F9B092A4F9",
 13522 => x"C0C0C0F9B092A4A4",
 13523 => x"C0C0C0F9B092A4B0",
 13524 => x"C0C0C0F9B092A499",
 13525 => x"C0C0C0F9B092A492",
 13526 => x"C0C0C0F9B092A482",
 13527 => x"C0C0C0F9B092A4F8",
 13528 => x"C0C0C0F9B092A480",
 13529 => x"C0C0C0F9B092A490",
 13530 => x"C0C0C0F9B092B0C0",
 13531 => x"C0C0C0F9B092B0F9",
 13532 => x"C0C0C0F9B092B0A4",
 13533 => x"C0C0C0F9B092B0B0",
 13534 => x"C0C0C0F9B092B099",
 13535 => x"C0C0C0F9B092B092",
 13536 => x"C0C0C0F9B092B082",
 13537 => x"C0C0C0F9B092B0F8",
 13538 => x"C0C0C0F9B092B080",
 13539 => x"C0C0C0F9B092B090",
 13540 => x"C0C0C0F9B09299C0",
 13541 => x"C0C0C0F9B09299F9",
 13542 => x"C0C0C0F9B09299A4",
 13543 => x"C0C0C0F9B09299B0",
 13544 => x"C0C0C0F9B0929999",
 13545 => x"C0C0C0F9B0929992",
 13546 => x"C0C0C0F9B0929982",
 13547 => x"C0C0C0F9B09299F8",
 13548 => x"C0C0C0F9B0929980",
 13549 => x"C0C0C0F9B0929990",
 13550 => x"C0C0C0F9B09292C0",
 13551 => x"C0C0C0F9B09292F9",
 13552 => x"C0C0C0F9B09292A4",
 13553 => x"C0C0C0F9B09292B0",
 13554 => x"C0C0C0F9B0929299",
 13555 => x"C0C0C0F9B0929292",
 13556 => x"C0C0C0F9B0929282",
 13557 => x"C0C0C0F9B09292F8",
 13558 => x"C0C0C0F9B0929280",
 13559 => x"C0C0C0F9B0929290",
 13560 => x"C0C0C0F9B09282C0",
 13561 => x"C0C0C0F9B09282F9",
 13562 => x"C0C0C0F9B09282A4",
 13563 => x"C0C0C0F9B09282B0",
 13564 => x"C0C0C0F9B0928299",
 13565 => x"C0C0C0F9B0928292",
 13566 => x"C0C0C0F9B0928282",
 13567 => x"C0C0C0F9B09282F8",
 13568 => x"C0C0C0F9B0928280",
 13569 => x"C0C0C0F9B0928290",
 13570 => x"C0C0C0F9B092F8C0",
 13571 => x"C0C0C0F9B092F8F9",
 13572 => x"C0C0C0F9B092F8A4",
 13573 => x"C0C0C0F9B092F8B0",
 13574 => x"C0C0C0F9B092F899",
 13575 => x"C0C0C0F9B092F892",
 13576 => x"C0C0C0F9B092F882",
 13577 => x"C0C0C0F9B092F8F8",
 13578 => x"C0C0C0F9B092F880",
 13579 => x"C0C0C0F9B092F890",
 13580 => x"C0C0C0F9B09280C0",
 13581 => x"C0C0C0F9B09280F9",
 13582 => x"C0C0C0F9B09280A4",
 13583 => x"C0C0C0F9B09280B0",
 13584 => x"C0C0C0F9B0928099",
 13585 => x"C0C0C0F9B0928092",
 13586 => x"C0C0C0F9B0928082",
 13587 => x"C0C0C0F9B09280F8",
 13588 => x"C0C0C0F9B0928080",
 13589 => x"C0C0C0F9B0928090",
 13590 => x"C0C0C0F9B09290C0",
 13591 => x"C0C0C0F9B09290F9",
 13592 => x"C0C0C0F9B09290A4",
 13593 => x"C0C0C0F9B09290B0",
 13594 => x"C0C0C0F9B0929099",
 13595 => x"C0C0C0F9B0929092",
 13596 => x"C0C0C0F9B0929082",
 13597 => x"C0C0C0F9B09290F8",
 13598 => x"C0C0C0F9B0929080",
 13599 => x"C0C0C0F9B0929090",
 13600 => x"C0C0C0F9B082C0C0",
 13601 => x"C0C0C0F9B082C0F9",
 13602 => x"C0C0C0F9B082C0A4",
 13603 => x"C0C0C0F9B082C0B0",
 13604 => x"C0C0C0F9B082C099",
 13605 => x"C0C0C0F9B082C092",
 13606 => x"C0C0C0F9B082C082",
 13607 => x"C0C0C0F9B082C0F8",
 13608 => x"C0C0C0F9B082C080",
 13609 => x"C0C0C0F9B082C090",
 13610 => x"C0C0C0F9B082F9C0",
 13611 => x"C0C0C0F9B082F9F9",
 13612 => x"C0C0C0F9B082F9A4",
 13613 => x"C0C0C0F9B082F9B0",
 13614 => x"C0C0C0F9B082F999",
 13615 => x"C0C0C0F9B082F992",
 13616 => x"C0C0C0F9B082F982",
 13617 => x"C0C0C0F9B082F9F8",
 13618 => x"C0C0C0F9B082F980",
 13619 => x"C0C0C0F9B082F990",
 13620 => x"C0C0C0F9B082A4C0",
 13621 => x"C0C0C0F9B082A4F9",
 13622 => x"C0C0C0F9B082A4A4",
 13623 => x"C0C0C0F9B082A4B0",
 13624 => x"C0C0C0F9B082A499",
 13625 => x"C0C0C0F9B082A492",
 13626 => x"C0C0C0F9B082A482",
 13627 => x"C0C0C0F9B082A4F8",
 13628 => x"C0C0C0F9B082A480",
 13629 => x"C0C0C0F9B082A490",
 13630 => x"C0C0C0F9B082B0C0",
 13631 => x"C0C0C0F9B082B0F9",
 13632 => x"C0C0C0F9B082B0A4",
 13633 => x"C0C0C0F9B082B0B0",
 13634 => x"C0C0C0F9B082B099",
 13635 => x"C0C0C0F9B082B092",
 13636 => x"C0C0C0F9B082B082",
 13637 => x"C0C0C0F9B082B0F8",
 13638 => x"C0C0C0F9B082B080",
 13639 => x"C0C0C0F9B082B090",
 13640 => x"C0C0C0F9B08299C0",
 13641 => x"C0C0C0F9B08299F9",
 13642 => x"C0C0C0F9B08299A4",
 13643 => x"C0C0C0F9B08299B0",
 13644 => x"C0C0C0F9B0829999",
 13645 => x"C0C0C0F9B0829992",
 13646 => x"C0C0C0F9B0829982",
 13647 => x"C0C0C0F9B08299F8",
 13648 => x"C0C0C0F9B0829980",
 13649 => x"C0C0C0F9B0829990",
 13650 => x"C0C0C0F9B08292C0",
 13651 => x"C0C0C0F9B08292F9",
 13652 => x"C0C0C0F9B08292A4",
 13653 => x"C0C0C0F9B08292B0",
 13654 => x"C0C0C0F9B0829299",
 13655 => x"C0C0C0F9B0829292",
 13656 => x"C0C0C0F9B0829282",
 13657 => x"C0C0C0F9B08292F8",
 13658 => x"C0C0C0F9B0829280",
 13659 => x"C0C0C0F9B0829290",
 13660 => x"C0C0C0F9B08282C0",
 13661 => x"C0C0C0F9B08282F9",
 13662 => x"C0C0C0F9B08282A4",
 13663 => x"C0C0C0F9B08282B0",
 13664 => x"C0C0C0F9B0828299",
 13665 => x"C0C0C0F9B0828292",
 13666 => x"C0C0C0F9B0828282",
 13667 => x"C0C0C0F9B08282F8",
 13668 => x"C0C0C0F9B0828280",
 13669 => x"C0C0C0F9B0828290",
 13670 => x"C0C0C0F9B082F8C0",
 13671 => x"C0C0C0F9B082F8F9",
 13672 => x"C0C0C0F9B082F8A4",
 13673 => x"C0C0C0F9B082F8B0",
 13674 => x"C0C0C0F9B082F899",
 13675 => x"C0C0C0F9B082F892",
 13676 => x"C0C0C0F9B082F882",
 13677 => x"C0C0C0F9B082F8F8",
 13678 => x"C0C0C0F9B082F880",
 13679 => x"C0C0C0F9B082F890",
 13680 => x"C0C0C0F9B08280C0",
 13681 => x"C0C0C0F9B08280F9",
 13682 => x"C0C0C0F9B08280A4",
 13683 => x"C0C0C0F9B08280B0",
 13684 => x"C0C0C0F9B0828099",
 13685 => x"C0C0C0F9B0828092",
 13686 => x"C0C0C0F9B0828082",
 13687 => x"C0C0C0F9B08280F8",
 13688 => x"C0C0C0F9B0828080",
 13689 => x"C0C0C0F9B0828090",
 13690 => x"C0C0C0F9B08290C0",
 13691 => x"C0C0C0F9B08290F9",
 13692 => x"C0C0C0F9B08290A4",
 13693 => x"C0C0C0F9B08290B0",
 13694 => x"C0C0C0F9B0829099",
 13695 => x"C0C0C0F9B0829092",
 13696 => x"C0C0C0F9B0829082",
 13697 => x"C0C0C0F9B08290F8",
 13698 => x"C0C0C0F9B0829080",
 13699 => x"C0C0C0F9B0829090",
 13700 => x"C0C0C0F9B0F8C0C0",
 13701 => x"C0C0C0F9B0F8C0F9",
 13702 => x"C0C0C0F9B0F8C0A4",
 13703 => x"C0C0C0F9B0F8C0B0",
 13704 => x"C0C0C0F9B0F8C099",
 13705 => x"C0C0C0F9B0F8C092",
 13706 => x"C0C0C0F9B0F8C082",
 13707 => x"C0C0C0F9B0F8C0F8",
 13708 => x"C0C0C0F9B0F8C080",
 13709 => x"C0C0C0F9B0F8C090",
 13710 => x"C0C0C0F9B0F8F9C0",
 13711 => x"C0C0C0F9B0F8F9F9",
 13712 => x"C0C0C0F9B0F8F9A4",
 13713 => x"C0C0C0F9B0F8F9B0",
 13714 => x"C0C0C0F9B0F8F999",
 13715 => x"C0C0C0F9B0F8F992",
 13716 => x"C0C0C0F9B0F8F982",
 13717 => x"C0C0C0F9B0F8F9F8",
 13718 => x"C0C0C0F9B0F8F980",
 13719 => x"C0C0C0F9B0F8F990",
 13720 => x"C0C0C0F9B0F8A4C0",
 13721 => x"C0C0C0F9B0F8A4F9",
 13722 => x"C0C0C0F9B0F8A4A4",
 13723 => x"C0C0C0F9B0F8A4B0",
 13724 => x"C0C0C0F9B0F8A499",
 13725 => x"C0C0C0F9B0F8A492",
 13726 => x"C0C0C0F9B0F8A482",
 13727 => x"C0C0C0F9B0F8A4F8",
 13728 => x"C0C0C0F9B0F8A480",
 13729 => x"C0C0C0F9B0F8A490",
 13730 => x"C0C0C0F9B0F8B0C0",
 13731 => x"C0C0C0F9B0F8B0F9",
 13732 => x"C0C0C0F9B0F8B0A4",
 13733 => x"C0C0C0F9B0F8B0B0",
 13734 => x"C0C0C0F9B0F8B099",
 13735 => x"C0C0C0F9B0F8B092",
 13736 => x"C0C0C0F9B0F8B082",
 13737 => x"C0C0C0F9B0F8B0F8",
 13738 => x"C0C0C0F9B0F8B080",
 13739 => x"C0C0C0F9B0F8B090",
 13740 => x"C0C0C0F9B0F899C0",
 13741 => x"C0C0C0F9B0F899F9",
 13742 => x"C0C0C0F9B0F899A4",
 13743 => x"C0C0C0F9B0F899B0",
 13744 => x"C0C0C0F9B0F89999",
 13745 => x"C0C0C0F9B0F89992",
 13746 => x"C0C0C0F9B0F89982",
 13747 => x"C0C0C0F9B0F899F8",
 13748 => x"C0C0C0F9B0F89980",
 13749 => x"C0C0C0F9B0F89990",
 13750 => x"C0C0C0F9B0F892C0",
 13751 => x"C0C0C0F9B0F892F9",
 13752 => x"C0C0C0F9B0F892A4",
 13753 => x"C0C0C0F9B0F892B0",
 13754 => x"C0C0C0F9B0F89299",
 13755 => x"C0C0C0F9B0F89292",
 13756 => x"C0C0C0F9B0F89282",
 13757 => x"C0C0C0F9B0F892F8",
 13758 => x"C0C0C0F9B0F89280",
 13759 => x"C0C0C0F9B0F89290",
 13760 => x"C0C0C0F9B0F882C0",
 13761 => x"C0C0C0F9B0F882F9",
 13762 => x"C0C0C0F9B0F882A4",
 13763 => x"C0C0C0F9B0F882B0",
 13764 => x"C0C0C0F9B0F88299",
 13765 => x"C0C0C0F9B0F88292",
 13766 => x"C0C0C0F9B0F88282",
 13767 => x"C0C0C0F9B0F882F8",
 13768 => x"C0C0C0F9B0F88280",
 13769 => x"C0C0C0F9B0F88290",
 13770 => x"C0C0C0F9B0F8F8C0",
 13771 => x"C0C0C0F9B0F8F8F9",
 13772 => x"C0C0C0F9B0F8F8A4",
 13773 => x"C0C0C0F9B0F8F8B0",
 13774 => x"C0C0C0F9B0F8F899",
 13775 => x"C0C0C0F9B0F8F892",
 13776 => x"C0C0C0F9B0F8F882",
 13777 => x"C0C0C0F9B0F8F8F8",
 13778 => x"C0C0C0F9B0F8F880",
 13779 => x"C0C0C0F9B0F8F890",
 13780 => x"C0C0C0F9B0F880C0",
 13781 => x"C0C0C0F9B0F880F9",
 13782 => x"C0C0C0F9B0F880A4",
 13783 => x"C0C0C0F9B0F880B0",
 13784 => x"C0C0C0F9B0F88099",
 13785 => x"C0C0C0F9B0F88092",
 13786 => x"C0C0C0F9B0F88082",
 13787 => x"C0C0C0F9B0F880F8",
 13788 => x"C0C0C0F9B0F88080",
 13789 => x"C0C0C0F9B0F88090",
 13790 => x"C0C0C0F9B0F890C0",
 13791 => x"C0C0C0F9B0F890F9",
 13792 => x"C0C0C0F9B0F890A4",
 13793 => x"C0C0C0F9B0F890B0",
 13794 => x"C0C0C0F9B0F89099",
 13795 => x"C0C0C0F9B0F89092",
 13796 => x"C0C0C0F9B0F89082",
 13797 => x"C0C0C0F9B0F890F8",
 13798 => x"C0C0C0F9B0F89080",
 13799 => x"C0C0C0F9B0F89090",
 13800 => x"C0C0C0F9B080C0C0",
 13801 => x"C0C0C0F9B080C0F9",
 13802 => x"C0C0C0F9B080C0A4",
 13803 => x"C0C0C0F9B080C0B0",
 13804 => x"C0C0C0F9B080C099",
 13805 => x"C0C0C0F9B080C092",
 13806 => x"C0C0C0F9B080C082",
 13807 => x"C0C0C0F9B080C0F8",
 13808 => x"C0C0C0F9B080C080",
 13809 => x"C0C0C0F9B080C090",
 13810 => x"C0C0C0F9B080F9C0",
 13811 => x"C0C0C0F9B080F9F9",
 13812 => x"C0C0C0F9B080F9A4",
 13813 => x"C0C0C0F9B080F9B0",
 13814 => x"C0C0C0F9B080F999",
 13815 => x"C0C0C0F9B080F992",
 13816 => x"C0C0C0F9B080F982",
 13817 => x"C0C0C0F9B080F9F8",
 13818 => x"C0C0C0F9B080F980",
 13819 => x"C0C0C0F9B080F990",
 13820 => x"C0C0C0F9B080A4C0",
 13821 => x"C0C0C0F9B080A4F9",
 13822 => x"C0C0C0F9B080A4A4",
 13823 => x"C0C0C0F9B080A4B0",
 13824 => x"C0C0C0F9B080A499",
 13825 => x"C0C0C0F9B080A492",
 13826 => x"C0C0C0F9B080A482",
 13827 => x"C0C0C0F9B080A4F8",
 13828 => x"C0C0C0F9B080A480",
 13829 => x"C0C0C0F9B080A490",
 13830 => x"C0C0C0F9B080B0C0",
 13831 => x"C0C0C0F9B080B0F9",
 13832 => x"C0C0C0F9B080B0A4",
 13833 => x"C0C0C0F9B080B0B0",
 13834 => x"C0C0C0F9B080B099",
 13835 => x"C0C0C0F9B080B092",
 13836 => x"C0C0C0F9B080B082",
 13837 => x"C0C0C0F9B080B0F8",
 13838 => x"C0C0C0F9B080B080",
 13839 => x"C0C0C0F9B080B090",
 13840 => x"C0C0C0F9B08099C0",
 13841 => x"C0C0C0F9B08099F9",
 13842 => x"C0C0C0F9B08099A4",
 13843 => x"C0C0C0F9B08099B0",
 13844 => x"C0C0C0F9B0809999",
 13845 => x"C0C0C0F9B0809992",
 13846 => x"C0C0C0F9B0809982",
 13847 => x"C0C0C0F9B08099F8",
 13848 => x"C0C0C0F9B0809980",
 13849 => x"C0C0C0F9B0809990",
 13850 => x"C0C0C0F9B08092C0",
 13851 => x"C0C0C0F9B08092F9",
 13852 => x"C0C0C0F9B08092A4",
 13853 => x"C0C0C0F9B08092B0",
 13854 => x"C0C0C0F9B0809299",
 13855 => x"C0C0C0F9B0809292",
 13856 => x"C0C0C0F9B0809282",
 13857 => x"C0C0C0F9B08092F8",
 13858 => x"C0C0C0F9B0809280",
 13859 => x"C0C0C0F9B0809290",
 13860 => x"C0C0C0F9B08082C0",
 13861 => x"C0C0C0F9B08082F9",
 13862 => x"C0C0C0F9B08082A4",
 13863 => x"C0C0C0F9B08082B0",
 13864 => x"C0C0C0F9B0808299",
 13865 => x"C0C0C0F9B0808292",
 13866 => x"C0C0C0F9B0808282",
 13867 => x"C0C0C0F9B08082F8",
 13868 => x"C0C0C0F9B0808280",
 13869 => x"C0C0C0F9B0808290",
 13870 => x"C0C0C0F9B080F8C0",
 13871 => x"C0C0C0F9B080F8F9",
 13872 => x"C0C0C0F9B080F8A4",
 13873 => x"C0C0C0F9B080F8B0",
 13874 => x"C0C0C0F9B080F899",
 13875 => x"C0C0C0F9B080F892",
 13876 => x"C0C0C0F9B080F882",
 13877 => x"C0C0C0F9B080F8F8",
 13878 => x"C0C0C0F9B080F880",
 13879 => x"C0C0C0F9B080F890",
 13880 => x"C0C0C0F9B08080C0",
 13881 => x"C0C0C0F9B08080F9",
 13882 => x"C0C0C0F9B08080A4",
 13883 => x"C0C0C0F9B08080B0",
 13884 => x"C0C0C0F9B0808099",
 13885 => x"C0C0C0F9B0808092",
 13886 => x"C0C0C0F9B0808082",
 13887 => x"C0C0C0F9B08080F8",
 13888 => x"C0C0C0F9B0808080",
 13889 => x"C0C0C0F9B0808090",
 13890 => x"C0C0C0F9B08090C0",
 13891 => x"C0C0C0F9B08090F9",
 13892 => x"C0C0C0F9B08090A4",
 13893 => x"C0C0C0F9B08090B0",
 13894 => x"C0C0C0F9B0809099",
 13895 => x"C0C0C0F9B0809092",
 13896 => x"C0C0C0F9B0809082",
 13897 => x"C0C0C0F9B08090F8",
 13898 => x"C0C0C0F9B0809080",
 13899 => x"C0C0C0F9B0809090",
 13900 => x"C0C0C0F9B090C0C0",
 13901 => x"C0C0C0F9B090C0F9",
 13902 => x"C0C0C0F9B090C0A4",
 13903 => x"C0C0C0F9B090C0B0",
 13904 => x"C0C0C0F9B090C099",
 13905 => x"C0C0C0F9B090C092",
 13906 => x"C0C0C0F9B090C082",
 13907 => x"C0C0C0F9B090C0F8",
 13908 => x"C0C0C0F9B090C080",
 13909 => x"C0C0C0F9B090C090",
 13910 => x"C0C0C0F9B090F9C0",
 13911 => x"C0C0C0F9B090F9F9",
 13912 => x"C0C0C0F9B090F9A4",
 13913 => x"C0C0C0F9B090F9B0",
 13914 => x"C0C0C0F9B090F999",
 13915 => x"C0C0C0F9B090F992",
 13916 => x"C0C0C0F9B090F982",
 13917 => x"C0C0C0F9B090F9F8",
 13918 => x"C0C0C0F9B090F980",
 13919 => x"C0C0C0F9B090F990",
 13920 => x"C0C0C0F9B090A4C0",
 13921 => x"C0C0C0F9B090A4F9",
 13922 => x"C0C0C0F9B090A4A4",
 13923 => x"C0C0C0F9B090A4B0",
 13924 => x"C0C0C0F9B090A499",
 13925 => x"C0C0C0F9B090A492",
 13926 => x"C0C0C0F9B090A482",
 13927 => x"C0C0C0F9B090A4F8",
 13928 => x"C0C0C0F9B090A480",
 13929 => x"C0C0C0F9B090A490",
 13930 => x"C0C0C0F9B090B0C0",
 13931 => x"C0C0C0F9B090B0F9",
 13932 => x"C0C0C0F9B090B0A4",
 13933 => x"C0C0C0F9B090B0B0",
 13934 => x"C0C0C0F9B090B099",
 13935 => x"C0C0C0F9B090B092",
 13936 => x"C0C0C0F9B090B082",
 13937 => x"C0C0C0F9B090B0F8",
 13938 => x"C0C0C0F9B090B080",
 13939 => x"C0C0C0F9B090B090",
 13940 => x"C0C0C0F9B09099C0",
 13941 => x"C0C0C0F9B09099F9",
 13942 => x"C0C0C0F9B09099A4",
 13943 => x"C0C0C0F9B09099B0",
 13944 => x"C0C0C0F9B0909999",
 13945 => x"C0C0C0F9B0909992",
 13946 => x"C0C0C0F9B0909982",
 13947 => x"C0C0C0F9B09099F8",
 13948 => x"C0C0C0F9B0909980",
 13949 => x"C0C0C0F9B0909990",
 13950 => x"C0C0C0F9B09092C0",
 13951 => x"C0C0C0F9B09092F9",
 13952 => x"C0C0C0F9B09092A4",
 13953 => x"C0C0C0F9B09092B0",
 13954 => x"C0C0C0F9B0909299",
 13955 => x"C0C0C0F9B0909292",
 13956 => x"C0C0C0F9B0909282",
 13957 => x"C0C0C0F9B09092F8",
 13958 => x"C0C0C0F9B0909280",
 13959 => x"C0C0C0F9B0909290",
 13960 => x"C0C0C0F9B09082C0",
 13961 => x"C0C0C0F9B09082F9",
 13962 => x"C0C0C0F9B09082A4",
 13963 => x"C0C0C0F9B09082B0",
 13964 => x"C0C0C0F9B0908299",
 13965 => x"C0C0C0F9B0908292",
 13966 => x"C0C0C0F9B0908282",
 13967 => x"C0C0C0F9B09082F8",
 13968 => x"C0C0C0F9B0908280",
 13969 => x"C0C0C0F9B0908290",
 13970 => x"C0C0C0F9B090F8C0",
 13971 => x"C0C0C0F9B090F8F9",
 13972 => x"C0C0C0F9B090F8A4",
 13973 => x"C0C0C0F9B090F8B0",
 13974 => x"C0C0C0F9B090F899",
 13975 => x"C0C0C0F9B090F892",
 13976 => x"C0C0C0F9B090F882",
 13977 => x"C0C0C0F9B090F8F8",
 13978 => x"C0C0C0F9B090F880",
 13979 => x"C0C0C0F9B090F890",
 13980 => x"C0C0C0F9B09080C0",
 13981 => x"C0C0C0F9B09080F9",
 13982 => x"C0C0C0F9B09080A4",
 13983 => x"C0C0C0F9B09080B0",
 13984 => x"C0C0C0F9B0908099",
 13985 => x"C0C0C0F9B0908092",
 13986 => x"C0C0C0F9B0908082",
 13987 => x"C0C0C0F9B09080F8",
 13988 => x"C0C0C0F9B0908080",
 13989 => x"C0C0C0F9B0908090",
 13990 => x"C0C0C0F9B09090C0",
 13991 => x"C0C0C0F9B09090F9",
 13992 => x"C0C0C0F9B09090A4",
 13993 => x"C0C0C0F9B09090B0",
 13994 => x"C0C0C0F9B0909099",
 13995 => x"C0C0C0F9B0909092",
 13996 => x"C0C0C0F9B0909082",
 13997 => x"C0C0C0F9B09090F8",
 13998 => x"C0C0C0F9B0909080",
 13999 => x"C0C0C0F9B0909090",
 14000 => x"C0C0C0F999C0C0C0",
 14001 => x"C0C0C0F999C0C0F9",
 14002 => x"C0C0C0F999C0C0A4",
 14003 => x"C0C0C0F999C0C0B0",
 14004 => x"C0C0C0F999C0C099",
 14005 => x"C0C0C0F999C0C092",
 14006 => x"C0C0C0F999C0C082",
 14007 => x"C0C0C0F999C0C0F8",
 14008 => x"C0C0C0F999C0C080",
 14009 => x"C0C0C0F999C0C090",
 14010 => x"C0C0C0F999C0F9C0",
 14011 => x"C0C0C0F999C0F9F9",
 14012 => x"C0C0C0F999C0F9A4",
 14013 => x"C0C0C0F999C0F9B0",
 14014 => x"C0C0C0F999C0F999",
 14015 => x"C0C0C0F999C0F992",
 14016 => x"C0C0C0F999C0F982",
 14017 => x"C0C0C0F999C0F9F8",
 14018 => x"C0C0C0F999C0F980",
 14019 => x"C0C0C0F999C0F990",
 14020 => x"C0C0C0F999C0A4C0",
 14021 => x"C0C0C0F999C0A4F9",
 14022 => x"C0C0C0F999C0A4A4",
 14023 => x"C0C0C0F999C0A4B0",
 14024 => x"C0C0C0F999C0A499",
 14025 => x"C0C0C0F999C0A492",
 14026 => x"C0C0C0F999C0A482",
 14027 => x"C0C0C0F999C0A4F8",
 14028 => x"C0C0C0F999C0A480",
 14029 => x"C0C0C0F999C0A490",
 14030 => x"C0C0C0F999C0B0C0",
 14031 => x"C0C0C0F999C0B0F9",
 14032 => x"C0C0C0F999C0B0A4",
 14033 => x"C0C0C0F999C0B0B0",
 14034 => x"C0C0C0F999C0B099",
 14035 => x"C0C0C0F999C0B092",
 14036 => x"C0C0C0F999C0B082",
 14037 => x"C0C0C0F999C0B0F8",
 14038 => x"C0C0C0F999C0B080",
 14039 => x"C0C0C0F999C0B090",
 14040 => x"C0C0C0F999C099C0",
 14041 => x"C0C0C0F999C099F9",
 14042 => x"C0C0C0F999C099A4",
 14043 => x"C0C0C0F999C099B0",
 14044 => x"C0C0C0F999C09999",
 14045 => x"C0C0C0F999C09992",
 14046 => x"C0C0C0F999C09982",
 14047 => x"C0C0C0F999C099F8",
 14048 => x"C0C0C0F999C09980",
 14049 => x"C0C0C0F999C09990",
 14050 => x"C0C0C0F999C092C0",
 14051 => x"C0C0C0F999C092F9",
 14052 => x"C0C0C0F999C092A4",
 14053 => x"C0C0C0F999C092B0",
 14054 => x"C0C0C0F999C09299",
 14055 => x"C0C0C0F999C09292",
 14056 => x"C0C0C0F999C09282",
 14057 => x"C0C0C0F999C092F8",
 14058 => x"C0C0C0F999C09280",
 14059 => x"C0C0C0F999C09290",
 14060 => x"C0C0C0F999C082C0",
 14061 => x"C0C0C0F999C082F9",
 14062 => x"C0C0C0F999C082A4",
 14063 => x"C0C0C0F999C082B0",
 14064 => x"C0C0C0F999C08299",
 14065 => x"C0C0C0F999C08292",
 14066 => x"C0C0C0F999C08282",
 14067 => x"C0C0C0F999C082F8",
 14068 => x"C0C0C0F999C08280",
 14069 => x"C0C0C0F999C08290",
 14070 => x"C0C0C0F999C0F8C0",
 14071 => x"C0C0C0F999C0F8F9",
 14072 => x"C0C0C0F999C0F8A4",
 14073 => x"C0C0C0F999C0F8B0",
 14074 => x"C0C0C0F999C0F899",
 14075 => x"C0C0C0F999C0F892",
 14076 => x"C0C0C0F999C0F882",
 14077 => x"C0C0C0F999C0F8F8",
 14078 => x"C0C0C0F999C0F880",
 14079 => x"C0C0C0F999C0F890",
 14080 => x"C0C0C0F999C080C0",
 14081 => x"C0C0C0F999C080F9",
 14082 => x"C0C0C0F999C080A4",
 14083 => x"C0C0C0F999C080B0",
 14084 => x"C0C0C0F999C08099",
 14085 => x"C0C0C0F999C08092",
 14086 => x"C0C0C0F999C08082",
 14087 => x"C0C0C0F999C080F8",
 14088 => x"C0C0C0F999C08080",
 14089 => x"C0C0C0F999C08090",
 14090 => x"C0C0C0F999C090C0",
 14091 => x"C0C0C0F999C090F9",
 14092 => x"C0C0C0F999C090A4",
 14093 => x"C0C0C0F999C090B0",
 14094 => x"C0C0C0F999C09099",
 14095 => x"C0C0C0F999C09092",
 14096 => x"C0C0C0F999C09082",
 14097 => x"C0C0C0F999C090F8",
 14098 => x"C0C0C0F999C09080",
 14099 => x"C0C0C0F999C09090",
 14100 => x"C0C0C0F999F9C0C0",
 14101 => x"C0C0C0F999F9C0F9",
 14102 => x"C0C0C0F999F9C0A4",
 14103 => x"C0C0C0F999F9C0B0",
 14104 => x"C0C0C0F999F9C099",
 14105 => x"C0C0C0F999F9C092",
 14106 => x"C0C0C0F999F9C082",
 14107 => x"C0C0C0F999F9C0F8",
 14108 => x"C0C0C0F999F9C080",
 14109 => x"C0C0C0F999F9C090",
 14110 => x"C0C0C0F999F9F9C0",
 14111 => x"C0C0C0F999F9F9F9",
 14112 => x"C0C0C0F999F9F9A4",
 14113 => x"C0C0C0F999F9F9B0",
 14114 => x"C0C0C0F999F9F999",
 14115 => x"C0C0C0F999F9F992",
 14116 => x"C0C0C0F999F9F982",
 14117 => x"C0C0C0F999F9F9F8",
 14118 => x"C0C0C0F999F9F980",
 14119 => x"C0C0C0F999F9F990",
 14120 => x"C0C0C0F999F9A4C0",
 14121 => x"C0C0C0F999F9A4F9",
 14122 => x"C0C0C0F999F9A4A4",
 14123 => x"C0C0C0F999F9A4B0",
 14124 => x"C0C0C0F999F9A499",
 14125 => x"C0C0C0F999F9A492",
 14126 => x"C0C0C0F999F9A482",
 14127 => x"C0C0C0F999F9A4F8",
 14128 => x"C0C0C0F999F9A480",
 14129 => x"C0C0C0F999F9A490",
 14130 => x"C0C0C0F999F9B0C0",
 14131 => x"C0C0C0F999F9B0F9",
 14132 => x"C0C0C0F999F9B0A4",
 14133 => x"C0C0C0F999F9B0B0",
 14134 => x"C0C0C0F999F9B099",
 14135 => x"C0C0C0F999F9B092",
 14136 => x"C0C0C0F999F9B082",
 14137 => x"C0C0C0F999F9B0F8",
 14138 => x"C0C0C0F999F9B080",
 14139 => x"C0C0C0F999F9B090",
 14140 => x"C0C0C0F999F999C0",
 14141 => x"C0C0C0F999F999F9",
 14142 => x"C0C0C0F999F999A4",
 14143 => x"C0C0C0F999F999B0",
 14144 => x"C0C0C0F999F99999",
 14145 => x"C0C0C0F999F99992",
 14146 => x"C0C0C0F999F99982",
 14147 => x"C0C0C0F999F999F8",
 14148 => x"C0C0C0F999F99980",
 14149 => x"C0C0C0F999F99990",
 14150 => x"C0C0C0F999F992C0",
 14151 => x"C0C0C0F999F992F9",
 14152 => x"C0C0C0F999F992A4",
 14153 => x"C0C0C0F999F992B0",
 14154 => x"C0C0C0F999F99299",
 14155 => x"C0C0C0F999F99292",
 14156 => x"C0C0C0F999F99282",
 14157 => x"C0C0C0F999F992F8",
 14158 => x"C0C0C0F999F99280",
 14159 => x"C0C0C0F999F99290",
 14160 => x"C0C0C0F999F982C0",
 14161 => x"C0C0C0F999F982F9",
 14162 => x"C0C0C0F999F982A4",
 14163 => x"C0C0C0F999F982B0",
 14164 => x"C0C0C0F999F98299",
 14165 => x"C0C0C0F999F98292",
 14166 => x"C0C0C0F999F98282",
 14167 => x"C0C0C0F999F982F8",
 14168 => x"C0C0C0F999F98280",
 14169 => x"C0C0C0F999F98290",
 14170 => x"C0C0C0F999F9F8C0",
 14171 => x"C0C0C0F999F9F8F9",
 14172 => x"C0C0C0F999F9F8A4",
 14173 => x"C0C0C0F999F9F8B0",
 14174 => x"C0C0C0F999F9F899",
 14175 => x"C0C0C0F999F9F892",
 14176 => x"C0C0C0F999F9F882",
 14177 => x"C0C0C0F999F9F8F8",
 14178 => x"C0C0C0F999F9F880",
 14179 => x"C0C0C0F999F9F890",
 14180 => x"C0C0C0F999F980C0",
 14181 => x"C0C0C0F999F980F9",
 14182 => x"C0C0C0F999F980A4",
 14183 => x"C0C0C0F999F980B0",
 14184 => x"C0C0C0F999F98099",
 14185 => x"C0C0C0F999F98092",
 14186 => x"C0C0C0F999F98082",
 14187 => x"C0C0C0F999F980F8",
 14188 => x"C0C0C0F999F98080",
 14189 => x"C0C0C0F999F98090",
 14190 => x"C0C0C0F999F990C0",
 14191 => x"C0C0C0F999F990F9",
 14192 => x"C0C0C0F999F990A4",
 14193 => x"C0C0C0F999F990B0",
 14194 => x"C0C0C0F999F99099",
 14195 => x"C0C0C0F999F99092",
 14196 => x"C0C0C0F999F99082",
 14197 => x"C0C0C0F999F990F8",
 14198 => x"C0C0C0F999F99080",
 14199 => x"C0C0C0F999F99090",
 14200 => x"C0C0C0F999A4C0C0",
 14201 => x"C0C0C0F999A4C0F9",
 14202 => x"C0C0C0F999A4C0A4",
 14203 => x"C0C0C0F999A4C0B0",
 14204 => x"C0C0C0F999A4C099",
 14205 => x"C0C0C0F999A4C092",
 14206 => x"C0C0C0F999A4C082",
 14207 => x"C0C0C0F999A4C0F8",
 14208 => x"C0C0C0F999A4C080",
 14209 => x"C0C0C0F999A4C090",
 14210 => x"C0C0C0F999A4F9C0",
 14211 => x"C0C0C0F999A4F9F9",
 14212 => x"C0C0C0F999A4F9A4",
 14213 => x"C0C0C0F999A4F9B0",
 14214 => x"C0C0C0F999A4F999",
 14215 => x"C0C0C0F999A4F992",
 14216 => x"C0C0C0F999A4F982",
 14217 => x"C0C0C0F999A4F9F8",
 14218 => x"C0C0C0F999A4F980",
 14219 => x"C0C0C0F999A4F990",
 14220 => x"C0C0C0F999A4A4C0",
 14221 => x"C0C0C0F999A4A4F9",
 14222 => x"C0C0C0F999A4A4A4",
 14223 => x"C0C0C0F999A4A4B0",
 14224 => x"C0C0C0F999A4A499",
 14225 => x"C0C0C0F999A4A492",
 14226 => x"C0C0C0F999A4A482",
 14227 => x"C0C0C0F999A4A4F8",
 14228 => x"C0C0C0F999A4A480",
 14229 => x"C0C0C0F999A4A490",
 14230 => x"C0C0C0F999A4B0C0",
 14231 => x"C0C0C0F999A4B0F9",
 14232 => x"C0C0C0F999A4B0A4",
 14233 => x"C0C0C0F999A4B0B0",
 14234 => x"C0C0C0F999A4B099",
 14235 => x"C0C0C0F999A4B092",
 14236 => x"C0C0C0F999A4B082",
 14237 => x"C0C0C0F999A4B0F8",
 14238 => x"C0C0C0F999A4B080",
 14239 => x"C0C0C0F999A4B090",
 14240 => x"C0C0C0F999A499C0",
 14241 => x"C0C0C0F999A499F9",
 14242 => x"C0C0C0F999A499A4",
 14243 => x"C0C0C0F999A499B0",
 14244 => x"C0C0C0F999A49999",
 14245 => x"C0C0C0F999A49992",
 14246 => x"C0C0C0F999A49982",
 14247 => x"C0C0C0F999A499F8",
 14248 => x"C0C0C0F999A49980",
 14249 => x"C0C0C0F999A49990",
 14250 => x"C0C0C0F999A492C0",
 14251 => x"C0C0C0F999A492F9",
 14252 => x"C0C0C0F999A492A4",
 14253 => x"C0C0C0F999A492B0",
 14254 => x"C0C0C0F999A49299",
 14255 => x"C0C0C0F999A49292",
 14256 => x"C0C0C0F999A49282",
 14257 => x"C0C0C0F999A492F8",
 14258 => x"C0C0C0F999A49280",
 14259 => x"C0C0C0F999A49290",
 14260 => x"C0C0C0F999A482C0",
 14261 => x"C0C0C0F999A482F9",
 14262 => x"C0C0C0F999A482A4",
 14263 => x"C0C0C0F999A482B0",
 14264 => x"C0C0C0F999A48299",
 14265 => x"C0C0C0F999A48292",
 14266 => x"C0C0C0F999A48282",
 14267 => x"C0C0C0F999A482F8",
 14268 => x"C0C0C0F999A48280",
 14269 => x"C0C0C0F999A48290",
 14270 => x"C0C0C0F999A4F8C0",
 14271 => x"C0C0C0F999A4F8F9",
 14272 => x"C0C0C0F999A4F8A4",
 14273 => x"C0C0C0F999A4F8B0",
 14274 => x"C0C0C0F999A4F899",
 14275 => x"C0C0C0F999A4F892",
 14276 => x"C0C0C0F999A4F882",
 14277 => x"C0C0C0F999A4F8F8",
 14278 => x"C0C0C0F999A4F880",
 14279 => x"C0C0C0F999A4F890",
 14280 => x"C0C0C0F999A480C0",
 14281 => x"C0C0C0F999A480F9",
 14282 => x"C0C0C0F999A480A4",
 14283 => x"C0C0C0F999A480B0",
 14284 => x"C0C0C0F999A48099",
 14285 => x"C0C0C0F999A48092",
 14286 => x"C0C0C0F999A48082",
 14287 => x"C0C0C0F999A480F8",
 14288 => x"C0C0C0F999A48080",
 14289 => x"C0C0C0F999A48090",
 14290 => x"C0C0C0F999A490C0",
 14291 => x"C0C0C0F999A490F9",
 14292 => x"C0C0C0F999A490A4",
 14293 => x"C0C0C0F999A490B0",
 14294 => x"C0C0C0F999A49099",
 14295 => x"C0C0C0F999A49092",
 14296 => x"C0C0C0F999A49082",
 14297 => x"C0C0C0F999A490F8",
 14298 => x"C0C0C0F999A49080",
 14299 => x"C0C0C0F999A49090",
 14300 => x"C0C0C0F999B0C0C0",
 14301 => x"C0C0C0F999B0C0F9",
 14302 => x"C0C0C0F999B0C0A4",
 14303 => x"C0C0C0F999B0C0B0",
 14304 => x"C0C0C0F999B0C099",
 14305 => x"C0C0C0F999B0C092",
 14306 => x"C0C0C0F999B0C082",
 14307 => x"C0C0C0F999B0C0F8",
 14308 => x"C0C0C0F999B0C080",
 14309 => x"C0C0C0F999B0C090",
 14310 => x"C0C0C0F999B0F9C0",
 14311 => x"C0C0C0F999B0F9F9",
 14312 => x"C0C0C0F999B0F9A4",
 14313 => x"C0C0C0F999B0F9B0",
 14314 => x"C0C0C0F999B0F999",
 14315 => x"C0C0C0F999B0F992",
 14316 => x"C0C0C0F999B0F982",
 14317 => x"C0C0C0F999B0F9F8",
 14318 => x"C0C0C0F999B0F980",
 14319 => x"C0C0C0F999B0F990",
 14320 => x"C0C0C0F999B0A4C0",
 14321 => x"C0C0C0F999B0A4F9",
 14322 => x"C0C0C0F999B0A4A4",
 14323 => x"C0C0C0F999B0A4B0",
 14324 => x"C0C0C0F999B0A499",
 14325 => x"C0C0C0F999B0A492",
 14326 => x"C0C0C0F999B0A482",
 14327 => x"C0C0C0F999B0A4F8",
 14328 => x"C0C0C0F999B0A480",
 14329 => x"C0C0C0F999B0A490",
 14330 => x"C0C0C0F999B0B0C0",
 14331 => x"C0C0C0F999B0B0F9",
 14332 => x"C0C0C0F999B0B0A4",
 14333 => x"C0C0C0F999B0B0B0",
 14334 => x"C0C0C0F999B0B099",
 14335 => x"C0C0C0F999B0B092",
 14336 => x"C0C0C0F999B0B082",
 14337 => x"C0C0C0F999B0B0F8",
 14338 => x"C0C0C0F999B0B080",
 14339 => x"C0C0C0F999B0B090",
 14340 => x"C0C0C0F999B099C0",
 14341 => x"C0C0C0F999B099F9",
 14342 => x"C0C0C0F999B099A4",
 14343 => x"C0C0C0F999B099B0",
 14344 => x"C0C0C0F999B09999",
 14345 => x"C0C0C0F999B09992",
 14346 => x"C0C0C0F999B09982",
 14347 => x"C0C0C0F999B099F8",
 14348 => x"C0C0C0F999B09980",
 14349 => x"C0C0C0F999B09990",
 14350 => x"C0C0C0F999B092C0",
 14351 => x"C0C0C0F999B092F9",
 14352 => x"C0C0C0F999B092A4",
 14353 => x"C0C0C0F999B092B0",
 14354 => x"C0C0C0F999B09299",
 14355 => x"C0C0C0F999B09292",
 14356 => x"C0C0C0F999B09282",
 14357 => x"C0C0C0F999B092F8",
 14358 => x"C0C0C0F999B09280",
 14359 => x"C0C0C0F999B09290",
 14360 => x"C0C0C0F999B082C0",
 14361 => x"C0C0C0F999B082F9",
 14362 => x"C0C0C0F999B082A4",
 14363 => x"C0C0C0F999B082B0",
 14364 => x"C0C0C0F999B08299",
 14365 => x"C0C0C0F999B08292",
 14366 => x"C0C0C0F999B08282",
 14367 => x"C0C0C0F999B082F8",
 14368 => x"C0C0C0F999B08280",
 14369 => x"C0C0C0F999B08290",
 14370 => x"C0C0C0F999B0F8C0",
 14371 => x"C0C0C0F999B0F8F9",
 14372 => x"C0C0C0F999B0F8A4",
 14373 => x"C0C0C0F999B0F8B0",
 14374 => x"C0C0C0F999B0F899",
 14375 => x"C0C0C0F999B0F892",
 14376 => x"C0C0C0F999B0F882",
 14377 => x"C0C0C0F999B0F8F8",
 14378 => x"C0C0C0F999B0F880",
 14379 => x"C0C0C0F999B0F890",
 14380 => x"C0C0C0F999B080C0",
 14381 => x"C0C0C0F999B080F9",
 14382 => x"C0C0C0F999B080A4",
 14383 => x"C0C0C0F999B080B0",
 14384 => x"C0C0C0F999B08099",
 14385 => x"C0C0C0F999B08092",
 14386 => x"C0C0C0F999B08082",
 14387 => x"C0C0C0F999B080F8",
 14388 => x"C0C0C0F999B08080",
 14389 => x"C0C0C0F999B08090",
 14390 => x"C0C0C0F999B090C0",
 14391 => x"C0C0C0F999B090F9",
 14392 => x"C0C0C0F999B090A4",
 14393 => x"C0C0C0F999B090B0",
 14394 => x"C0C0C0F999B09099",
 14395 => x"C0C0C0F999B09092",
 14396 => x"C0C0C0F999B09082",
 14397 => x"C0C0C0F999B090F8",
 14398 => x"C0C0C0F999B09080",
 14399 => x"C0C0C0F999B09090",
 14400 => x"C0C0C0F99999C0C0",
 14401 => x"C0C0C0F99999C0F9",
 14402 => x"C0C0C0F99999C0A4",
 14403 => x"C0C0C0F99999C0B0",
 14404 => x"C0C0C0F99999C099",
 14405 => x"C0C0C0F99999C092",
 14406 => x"C0C0C0F99999C082",
 14407 => x"C0C0C0F99999C0F8",
 14408 => x"C0C0C0F99999C080",
 14409 => x"C0C0C0F99999C090",
 14410 => x"C0C0C0F99999F9C0",
 14411 => x"C0C0C0F99999F9F9",
 14412 => x"C0C0C0F99999F9A4",
 14413 => x"C0C0C0F99999F9B0",
 14414 => x"C0C0C0F99999F999",
 14415 => x"C0C0C0F99999F992",
 14416 => x"C0C0C0F99999F982",
 14417 => x"C0C0C0F99999F9F8",
 14418 => x"C0C0C0F99999F980",
 14419 => x"C0C0C0F99999F990",
 14420 => x"C0C0C0F99999A4C0",
 14421 => x"C0C0C0F99999A4F9",
 14422 => x"C0C0C0F99999A4A4",
 14423 => x"C0C0C0F99999A4B0",
 14424 => x"C0C0C0F99999A499",
 14425 => x"C0C0C0F99999A492",
 14426 => x"C0C0C0F99999A482",
 14427 => x"C0C0C0F99999A4F8",
 14428 => x"C0C0C0F99999A480",
 14429 => x"C0C0C0F99999A490",
 14430 => x"C0C0C0F99999B0C0",
 14431 => x"C0C0C0F99999B0F9",
 14432 => x"C0C0C0F99999B0A4",
 14433 => x"C0C0C0F99999B0B0",
 14434 => x"C0C0C0F99999B099",
 14435 => x"C0C0C0F99999B092",
 14436 => x"C0C0C0F99999B082",
 14437 => x"C0C0C0F99999B0F8",
 14438 => x"C0C0C0F99999B080",
 14439 => x"C0C0C0F99999B090",
 14440 => x"C0C0C0F9999999C0",
 14441 => x"C0C0C0F9999999F9",
 14442 => x"C0C0C0F9999999A4",
 14443 => x"C0C0C0F9999999B0",
 14444 => x"C0C0C0F999999999",
 14445 => x"C0C0C0F999999992",
 14446 => x"C0C0C0F999999982",
 14447 => x"C0C0C0F9999999F8",
 14448 => x"C0C0C0F999999980",
 14449 => x"C0C0C0F999999990",
 14450 => x"C0C0C0F9999992C0",
 14451 => x"C0C0C0F9999992F9",
 14452 => x"C0C0C0F9999992A4",
 14453 => x"C0C0C0F9999992B0",
 14454 => x"C0C0C0F999999299",
 14455 => x"C0C0C0F999999292",
 14456 => x"C0C0C0F999999282",
 14457 => x"C0C0C0F9999992F8",
 14458 => x"C0C0C0F999999280",
 14459 => x"C0C0C0F999999290",
 14460 => x"C0C0C0F9999982C0",
 14461 => x"C0C0C0F9999982F9",
 14462 => x"C0C0C0F9999982A4",
 14463 => x"C0C0C0F9999982B0",
 14464 => x"C0C0C0F999998299",
 14465 => x"C0C0C0F999998292",
 14466 => x"C0C0C0F999998282",
 14467 => x"C0C0C0F9999982F8",
 14468 => x"C0C0C0F999998280",
 14469 => x"C0C0C0F999998290",
 14470 => x"C0C0C0F99999F8C0",
 14471 => x"C0C0C0F99999F8F9",
 14472 => x"C0C0C0F99999F8A4",
 14473 => x"C0C0C0F99999F8B0",
 14474 => x"C0C0C0F99999F899",
 14475 => x"C0C0C0F99999F892",
 14476 => x"C0C0C0F99999F882",
 14477 => x"C0C0C0F99999F8F8",
 14478 => x"C0C0C0F99999F880",
 14479 => x"C0C0C0F99999F890",
 14480 => x"C0C0C0F9999980C0",
 14481 => x"C0C0C0F9999980F9",
 14482 => x"C0C0C0F9999980A4",
 14483 => x"C0C0C0F9999980B0",
 14484 => x"C0C0C0F999998099",
 14485 => x"C0C0C0F999998092",
 14486 => x"C0C0C0F999998082",
 14487 => x"C0C0C0F9999980F8",
 14488 => x"C0C0C0F999998080",
 14489 => x"C0C0C0F999998090",
 14490 => x"C0C0C0F9999990C0",
 14491 => x"C0C0C0F9999990F9",
 14492 => x"C0C0C0F9999990A4",
 14493 => x"C0C0C0F9999990B0",
 14494 => x"C0C0C0F999999099",
 14495 => x"C0C0C0F999999092",
 14496 => x"C0C0C0F999999082",
 14497 => x"C0C0C0F9999990F8",
 14498 => x"C0C0C0F999999080",
 14499 => x"C0C0C0F999999090",
 14500 => x"C0C0C0F99992C0C0",
 14501 => x"C0C0C0F99992C0F9",
 14502 => x"C0C0C0F99992C0A4",
 14503 => x"C0C0C0F99992C0B0",
 14504 => x"C0C0C0F99992C099",
 14505 => x"C0C0C0F99992C092",
 14506 => x"C0C0C0F99992C082",
 14507 => x"C0C0C0F99992C0F8",
 14508 => x"C0C0C0F99992C080",
 14509 => x"C0C0C0F99992C090",
 14510 => x"C0C0C0F99992F9C0",
 14511 => x"C0C0C0F99992F9F9",
 14512 => x"C0C0C0F99992F9A4",
 14513 => x"C0C0C0F99992F9B0",
 14514 => x"C0C0C0F99992F999",
 14515 => x"C0C0C0F99992F992",
 14516 => x"C0C0C0F99992F982",
 14517 => x"C0C0C0F99992F9F8",
 14518 => x"C0C0C0F99992F980",
 14519 => x"C0C0C0F99992F990",
 14520 => x"C0C0C0F99992A4C0",
 14521 => x"C0C0C0F99992A4F9",
 14522 => x"C0C0C0F99992A4A4",
 14523 => x"C0C0C0F99992A4B0",
 14524 => x"C0C0C0F99992A499",
 14525 => x"C0C0C0F99992A492",
 14526 => x"C0C0C0F99992A482",
 14527 => x"C0C0C0F99992A4F8",
 14528 => x"C0C0C0F99992A480",
 14529 => x"C0C0C0F99992A490",
 14530 => x"C0C0C0F99992B0C0",
 14531 => x"C0C0C0F99992B0F9",
 14532 => x"C0C0C0F99992B0A4",
 14533 => x"C0C0C0F99992B0B0",
 14534 => x"C0C0C0F99992B099",
 14535 => x"C0C0C0F99992B092",
 14536 => x"C0C0C0F99992B082",
 14537 => x"C0C0C0F99992B0F8",
 14538 => x"C0C0C0F99992B080",
 14539 => x"C0C0C0F99992B090",
 14540 => x"C0C0C0F9999299C0",
 14541 => x"C0C0C0F9999299F9",
 14542 => x"C0C0C0F9999299A4",
 14543 => x"C0C0C0F9999299B0",
 14544 => x"C0C0C0F999929999",
 14545 => x"C0C0C0F999929992",
 14546 => x"C0C0C0F999929982",
 14547 => x"C0C0C0F9999299F8",
 14548 => x"C0C0C0F999929980",
 14549 => x"C0C0C0F999929990",
 14550 => x"C0C0C0F9999292C0",
 14551 => x"C0C0C0F9999292F9",
 14552 => x"C0C0C0F9999292A4",
 14553 => x"C0C0C0F9999292B0",
 14554 => x"C0C0C0F999929299",
 14555 => x"C0C0C0F999929292",
 14556 => x"C0C0C0F999929282",
 14557 => x"C0C0C0F9999292F8",
 14558 => x"C0C0C0F999929280",
 14559 => x"C0C0C0F999929290",
 14560 => x"C0C0C0F9999282C0",
 14561 => x"C0C0C0F9999282F9",
 14562 => x"C0C0C0F9999282A4",
 14563 => x"C0C0C0F9999282B0",
 14564 => x"C0C0C0F999928299",
 14565 => x"C0C0C0F999928292",
 14566 => x"C0C0C0F999928282",
 14567 => x"C0C0C0F9999282F8",
 14568 => x"C0C0C0F999928280",
 14569 => x"C0C0C0F999928290",
 14570 => x"C0C0C0F99992F8C0",
 14571 => x"C0C0C0F99992F8F9",
 14572 => x"C0C0C0F99992F8A4",
 14573 => x"C0C0C0F99992F8B0",
 14574 => x"C0C0C0F99992F899",
 14575 => x"C0C0C0F99992F892",
 14576 => x"C0C0C0F99992F882",
 14577 => x"C0C0C0F99992F8F8",
 14578 => x"C0C0C0F99992F880",
 14579 => x"C0C0C0F99992F890",
 14580 => x"C0C0C0F9999280C0",
 14581 => x"C0C0C0F9999280F9",
 14582 => x"C0C0C0F9999280A4",
 14583 => x"C0C0C0F9999280B0",
 14584 => x"C0C0C0F999928099",
 14585 => x"C0C0C0F999928092",
 14586 => x"C0C0C0F999928082",
 14587 => x"C0C0C0F9999280F8",
 14588 => x"C0C0C0F999928080",
 14589 => x"C0C0C0F999928090",
 14590 => x"C0C0C0F9999290C0",
 14591 => x"C0C0C0F9999290F9",
 14592 => x"C0C0C0F9999290A4",
 14593 => x"C0C0C0F9999290B0",
 14594 => x"C0C0C0F999929099",
 14595 => x"C0C0C0F999929092",
 14596 => x"C0C0C0F999929082",
 14597 => x"C0C0C0F9999290F8",
 14598 => x"C0C0C0F999929080",
 14599 => x"C0C0C0F999929090",
 14600 => x"C0C0C0F99982C0C0",
 14601 => x"C0C0C0F99982C0F9",
 14602 => x"C0C0C0F99982C0A4",
 14603 => x"C0C0C0F99982C0B0",
 14604 => x"C0C0C0F99982C099",
 14605 => x"C0C0C0F99982C092",
 14606 => x"C0C0C0F99982C082",
 14607 => x"C0C0C0F99982C0F8",
 14608 => x"C0C0C0F99982C080",
 14609 => x"C0C0C0F99982C090",
 14610 => x"C0C0C0F99982F9C0",
 14611 => x"C0C0C0F99982F9F9",
 14612 => x"C0C0C0F99982F9A4",
 14613 => x"C0C0C0F99982F9B0",
 14614 => x"C0C0C0F99982F999",
 14615 => x"C0C0C0F99982F992",
 14616 => x"C0C0C0F99982F982",
 14617 => x"C0C0C0F99982F9F8",
 14618 => x"C0C0C0F99982F980",
 14619 => x"C0C0C0F99982F990",
 14620 => x"C0C0C0F99982A4C0",
 14621 => x"C0C0C0F99982A4F9",
 14622 => x"C0C0C0F99982A4A4",
 14623 => x"C0C0C0F99982A4B0",
 14624 => x"C0C0C0F99982A499",
 14625 => x"C0C0C0F99982A492",
 14626 => x"C0C0C0F99982A482",
 14627 => x"C0C0C0F99982A4F8",
 14628 => x"C0C0C0F99982A480",
 14629 => x"C0C0C0F99982A490",
 14630 => x"C0C0C0F99982B0C0",
 14631 => x"C0C0C0F99982B0F9",
 14632 => x"C0C0C0F99982B0A4",
 14633 => x"C0C0C0F99982B0B0",
 14634 => x"C0C0C0F99982B099",
 14635 => x"C0C0C0F99982B092",
 14636 => x"C0C0C0F99982B082",
 14637 => x"C0C0C0F99982B0F8",
 14638 => x"C0C0C0F99982B080",
 14639 => x"C0C0C0F99982B090",
 14640 => x"C0C0C0F9998299C0",
 14641 => x"C0C0C0F9998299F9",
 14642 => x"C0C0C0F9998299A4",
 14643 => x"C0C0C0F9998299B0",
 14644 => x"C0C0C0F999829999",
 14645 => x"C0C0C0F999829992",
 14646 => x"C0C0C0F999829982",
 14647 => x"C0C0C0F9998299F8",
 14648 => x"C0C0C0F999829980",
 14649 => x"C0C0C0F999829990",
 14650 => x"C0C0C0F9998292C0",
 14651 => x"C0C0C0F9998292F9",
 14652 => x"C0C0C0F9998292A4",
 14653 => x"C0C0C0F9998292B0",
 14654 => x"C0C0C0F999829299",
 14655 => x"C0C0C0F999829292",
 14656 => x"C0C0C0F999829282",
 14657 => x"C0C0C0F9998292F8",
 14658 => x"C0C0C0F999829280",
 14659 => x"C0C0C0F999829290",
 14660 => x"C0C0C0F9998282C0",
 14661 => x"C0C0C0F9998282F9",
 14662 => x"C0C0C0F9998282A4",
 14663 => x"C0C0C0F9998282B0",
 14664 => x"C0C0C0F999828299",
 14665 => x"C0C0C0F999828292",
 14666 => x"C0C0C0F999828282",
 14667 => x"C0C0C0F9998282F8",
 14668 => x"C0C0C0F999828280",
 14669 => x"C0C0C0F999828290",
 14670 => x"C0C0C0F99982F8C0",
 14671 => x"C0C0C0F99982F8F9",
 14672 => x"C0C0C0F99982F8A4",
 14673 => x"C0C0C0F99982F8B0",
 14674 => x"C0C0C0F99982F899",
 14675 => x"C0C0C0F99982F892",
 14676 => x"C0C0C0F99982F882",
 14677 => x"C0C0C0F99982F8F8",
 14678 => x"C0C0C0F99982F880",
 14679 => x"C0C0C0F99982F890",
 14680 => x"C0C0C0F9998280C0",
 14681 => x"C0C0C0F9998280F9",
 14682 => x"C0C0C0F9998280A4",
 14683 => x"C0C0C0F9998280B0",
 14684 => x"C0C0C0F999828099",
 14685 => x"C0C0C0F999828092",
 14686 => x"C0C0C0F999828082",
 14687 => x"C0C0C0F9998280F8",
 14688 => x"C0C0C0F999828080",
 14689 => x"C0C0C0F999828090",
 14690 => x"C0C0C0F9998290C0",
 14691 => x"C0C0C0F9998290F9",
 14692 => x"C0C0C0F9998290A4",
 14693 => x"C0C0C0F9998290B0",
 14694 => x"C0C0C0F999829099",
 14695 => x"C0C0C0F999829092",
 14696 => x"C0C0C0F999829082",
 14697 => x"C0C0C0F9998290F8",
 14698 => x"C0C0C0F999829080",
 14699 => x"C0C0C0F999829090",
 14700 => x"C0C0C0F999F8C0C0",
 14701 => x"C0C0C0F999F8C0F9",
 14702 => x"C0C0C0F999F8C0A4",
 14703 => x"C0C0C0F999F8C0B0",
 14704 => x"C0C0C0F999F8C099",
 14705 => x"C0C0C0F999F8C092",
 14706 => x"C0C0C0F999F8C082",
 14707 => x"C0C0C0F999F8C0F8",
 14708 => x"C0C0C0F999F8C080",
 14709 => x"C0C0C0F999F8C090",
 14710 => x"C0C0C0F999F8F9C0",
 14711 => x"C0C0C0F999F8F9F9",
 14712 => x"C0C0C0F999F8F9A4",
 14713 => x"C0C0C0F999F8F9B0",
 14714 => x"C0C0C0F999F8F999",
 14715 => x"C0C0C0F999F8F992",
 14716 => x"C0C0C0F999F8F982",
 14717 => x"C0C0C0F999F8F9F8",
 14718 => x"C0C0C0F999F8F980",
 14719 => x"C0C0C0F999F8F990",
 14720 => x"C0C0C0F999F8A4C0",
 14721 => x"C0C0C0F999F8A4F9",
 14722 => x"C0C0C0F999F8A4A4",
 14723 => x"C0C0C0F999F8A4B0",
 14724 => x"C0C0C0F999F8A499",
 14725 => x"C0C0C0F999F8A492",
 14726 => x"C0C0C0F999F8A482",
 14727 => x"C0C0C0F999F8A4F8",
 14728 => x"C0C0C0F999F8A480",
 14729 => x"C0C0C0F999F8A490",
 14730 => x"C0C0C0F999F8B0C0",
 14731 => x"C0C0C0F999F8B0F9",
 14732 => x"C0C0C0F999F8B0A4",
 14733 => x"C0C0C0F999F8B0B0",
 14734 => x"C0C0C0F999F8B099",
 14735 => x"C0C0C0F999F8B092",
 14736 => x"C0C0C0F999F8B082",
 14737 => x"C0C0C0F999F8B0F8",
 14738 => x"C0C0C0F999F8B080",
 14739 => x"C0C0C0F999F8B090",
 14740 => x"C0C0C0F999F899C0",
 14741 => x"C0C0C0F999F899F9",
 14742 => x"C0C0C0F999F899A4",
 14743 => x"C0C0C0F999F899B0",
 14744 => x"C0C0C0F999F89999",
 14745 => x"C0C0C0F999F89992",
 14746 => x"C0C0C0F999F89982",
 14747 => x"C0C0C0F999F899F8",
 14748 => x"C0C0C0F999F89980",
 14749 => x"C0C0C0F999F89990",
 14750 => x"C0C0C0F999F892C0",
 14751 => x"C0C0C0F999F892F9",
 14752 => x"C0C0C0F999F892A4",
 14753 => x"C0C0C0F999F892B0",
 14754 => x"C0C0C0F999F89299",
 14755 => x"C0C0C0F999F89292",
 14756 => x"C0C0C0F999F89282",
 14757 => x"C0C0C0F999F892F8",
 14758 => x"C0C0C0F999F89280",
 14759 => x"C0C0C0F999F89290",
 14760 => x"C0C0C0F999F882C0",
 14761 => x"C0C0C0F999F882F9",
 14762 => x"C0C0C0F999F882A4",
 14763 => x"C0C0C0F999F882B0",
 14764 => x"C0C0C0F999F88299",
 14765 => x"C0C0C0F999F88292",
 14766 => x"C0C0C0F999F88282",
 14767 => x"C0C0C0F999F882F8",
 14768 => x"C0C0C0F999F88280",
 14769 => x"C0C0C0F999F88290",
 14770 => x"C0C0C0F999F8F8C0",
 14771 => x"C0C0C0F999F8F8F9",
 14772 => x"C0C0C0F999F8F8A4",
 14773 => x"C0C0C0F999F8F8B0",
 14774 => x"C0C0C0F999F8F899",
 14775 => x"C0C0C0F999F8F892",
 14776 => x"C0C0C0F999F8F882",
 14777 => x"C0C0C0F999F8F8F8",
 14778 => x"C0C0C0F999F8F880",
 14779 => x"C0C0C0F999F8F890",
 14780 => x"C0C0C0F999F880C0",
 14781 => x"C0C0C0F999F880F9",
 14782 => x"C0C0C0F999F880A4",
 14783 => x"C0C0C0F999F880B0",
 14784 => x"C0C0C0F999F88099",
 14785 => x"C0C0C0F999F88092",
 14786 => x"C0C0C0F999F88082",
 14787 => x"C0C0C0F999F880F8",
 14788 => x"C0C0C0F999F88080",
 14789 => x"C0C0C0F999F88090",
 14790 => x"C0C0C0F999F890C0",
 14791 => x"C0C0C0F999F890F9",
 14792 => x"C0C0C0F999F890A4",
 14793 => x"C0C0C0F999F890B0",
 14794 => x"C0C0C0F999F89099",
 14795 => x"C0C0C0F999F89092",
 14796 => x"C0C0C0F999F89082",
 14797 => x"C0C0C0F999F890F8",
 14798 => x"C0C0C0F999F89080",
 14799 => x"C0C0C0F999F89090",
 14800 => x"C0C0C0F99980C0C0",
 14801 => x"C0C0C0F99980C0F9",
 14802 => x"C0C0C0F99980C0A4",
 14803 => x"C0C0C0F99980C0B0",
 14804 => x"C0C0C0F99980C099",
 14805 => x"C0C0C0F99980C092",
 14806 => x"C0C0C0F99980C082",
 14807 => x"C0C0C0F99980C0F8",
 14808 => x"C0C0C0F99980C080",
 14809 => x"C0C0C0F99980C090",
 14810 => x"C0C0C0F99980F9C0",
 14811 => x"C0C0C0F99980F9F9",
 14812 => x"C0C0C0F99980F9A4",
 14813 => x"C0C0C0F99980F9B0",
 14814 => x"C0C0C0F99980F999",
 14815 => x"C0C0C0F99980F992",
 14816 => x"C0C0C0F99980F982",
 14817 => x"C0C0C0F99980F9F8",
 14818 => x"C0C0C0F99980F980",
 14819 => x"C0C0C0F99980F990",
 14820 => x"C0C0C0F99980A4C0",
 14821 => x"C0C0C0F99980A4F9",
 14822 => x"C0C0C0F99980A4A4",
 14823 => x"C0C0C0F99980A4B0",
 14824 => x"C0C0C0F99980A499",
 14825 => x"C0C0C0F99980A492",
 14826 => x"C0C0C0F99980A482",
 14827 => x"C0C0C0F99980A4F8",
 14828 => x"C0C0C0F99980A480",
 14829 => x"C0C0C0F99980A490",
 14830 => x"C0C0C0F99980B0C0",
 14831 => x"C0C0C0F99980B0F9",
 14832 => x"C0C0C0F99980B0A4",
 14833 => x"C0C0C0F99980B0B0",
 14834 => x"C0C0C0F99980B099",
 14835 => x"C0C0C0F99980B092",
 14836 => x"C0C0C0F99980B082",
 14837 => x"C0C0C0F99980B0F8",
 14838 => x"C0C0C0F99980B080",
 14839 => x"C0C0C0F99980B090",
 14840 => x"C0C0C0F9998099C0",
 14841 => x"C0C0C0F9998099F9",
 14842 => x"C0C0C0F9998099A4",
 14843 => x"C0C0C0F9998099B0",
 14844 => x"C0C0C0F999809999",
 14845 => x"C0C0C0F999809992",
 14846 => x"C0C0C0F999809982",
 14847 => x"C0C0C0F9998099F8",
 14848 => x"C0C0C0F999809980",
 14849 => x"C0C0C0F999809990",
 14850 => x"C0C0C0F9998092C0",
 14851 => x"C0C0C0F9998092F9",
 14852 => x"C0C0C0F9998092A4",
 14853 => x"C0C0C0F9998092B0",
 14854 => x"C0C0C0F999809299",
 14855 => x"C0C0C0F999809292",
 14856 => x"C0C0C0F999809282",
 14857 => x"C0C0C0F9998092F8",
 14858 => x"C0C0C0F999809280",
 14859 => x"C0C0C0F999809290",
 14860 => x"C0C0C0F9998082C0",
 14861 => x"C0C0C0F9998082F9",
 14862 => x"C0C0C0F9998082A4",
 14863 => x"C0C0C0F9998082B0",
 14864 => x"C0C0C0F999808299",
 14865 => x"C0C0C0F999808292",
 14866 => x"C0C0C0F999808282",
 14867 => x"C0C0C0F9998082F8",
 14868 => x"C0C0C0F999808280",
 14869 => x"C0C0C0F999808290",
 14870 => x"C0C0C0F99980F8C0",
 14871 => x"C0C0C0F99980F8F9",
 14872 => x"C0C0C0F99980F8A4",
 14873 => x"C0C0C0F99980F8B0",
 14874 => x"C0C0C0F99980F899",
 14875 => x"C0C0C0F99980F892",
 14876 => x"C0C0C0F99980F882",
 14877 => x"C0C0C0F99980F8F8",
 14878 => x"C0C0C0F99980F880",
 14879 => x"C0C0C0F99980F890",
 14880 => x"C0C0C0F9998080C0",
 14881 => x"C0C0C0F9998080F9",
 14882 => x"C0C0C0F9998080A4",
 14883 => x"C0C0C0F9998080B0",
 14884 => x"C0C0C0F999808099",
 14885 => x"C0C0C0F999808092",
 14886 => x"C0C0C0F999808082",
 14887 => x"C0C0C0F9998080F8",
 14888 => x"C0C0C0F999808080",
 14889 => x"C0C0C0F999808090",
 14890 => x"C0C0C0F9998090C0",
 14891 => x"C0C0C0F9998090F9",
 14892 => x"C0C0C0F9998090A4",
 14893 => x"C0C0C0F9998090B0",
 14894 => x"C0C0C0F999809099",
 14895 => x"C0C0C0F999809092",
 14896 => x"C0C0C0F999809082",
 14897 => x"C0C0C0F9998090F8",
 14898 => x"C0C0C0F999809080",
 14899 => x"C0C0C0F999809090",
 14900 => x"C0C0C0F99990C0C0",
 14901 => x"C0C0C0F99990C0F9",
 14902 => x"C0C0C0F99990C0A4",
 14903 => x"C0C0C0F99990C0B0",
 14904 => x"C0C0C0F99990C099",
 14905 => x"C0C0C0F99990C092",
 14906 => x"C0C0C0F99990C082",
 14907 => x"C0C0C0F99990C0F8",
 14908 => x"C0C0C0F99990C080",
 14909 => x"C0C0C0F99990C090",
 14910 => x"C0C0C0F99990F9C0",
 14911 => x"C0C0C0F99990F9F9",
 14912 => x"C0C0C0F99990F9A4",
 14913 => x"C0C0C0F99990F9B0",
 14914 => x"C0C0C0F99990F999",
 14915 => x"C0C0C0F99990F992",
 14916 => x"C0C0C0F99990F982",
 14917 => x"C0C0C0F99990F9F8",
 14918 => x"C0C0C0F99990F980",
 14919 => x"C0C0C0F99990F990",
 14920 => x"C0C0C0F99990A4C0",
 14921 => x"C0C0C0F99990A4F9",
 14922 => x"C0C0C0F99990A4A4",
 14923 => x"C0C0C0F99990A4B0",
 14924 => x"C0C0C0F99990A499",
 14925 => x"C0C0C0F99990A492",
 14926 => x"C0C0C0F99990A482",
 14927 => x"C0C0C0F99990A4F8",
 14928 => x"C0C0C0F99990A480",
 14929 => x"C0C0C0F99990A490",
 14930 => x"C0C0C0F99990B0C0",
 14931 => x"C0C0C0F99990B0F9",
 14932 => x"C0C0C0F99990B0A4",
 14933 => x"C0C0C0F99990B0B0",
 14934 => x"C0C0C0F99990B099",
 14935 => x"C0C0C0F99990B092",
 14936 => x"C0C0C0F99990B082",
 14937 => x"C0C0C0F99990B0F8",
 14938 => x"C0C0C0F99990B080",
 14939 => x"C0C0C0F99990B090",
 14940 => x"C0C0C0F9999099C0",
 14941 => x"C0C0C0F9999099F9",
 14942 => x"C0C0C0F9999099A4",
 14943 => x"C0C0C0F9999099B0",
 14944 => x"C0C0C0F999909999",
 14945 => x"C0C0C0F999909992",
 14946 => x"C0C0C0F999909982",
 14947 => x"C0C0C0F9999099F8",
 14948 => x"C0C0C0F999909980",
 14949 => x"C0C0C0F999909990",
 14950 => x"C0C0C0F9999092C0",
 14951 => x"C0C0C0F9999092F9",
 14952 => x"C0C0C0F9999092A4",
 14953 => x"C0C0C0F9999092B0",
 14954 => x"C0C0C0F999909299",
 14955 => x"C0C0C0F999909292",
 14956 => x"C0C0C0F999909282",
 14957 => x"C0C0C0F9999092F8",
 14958 => x"C0C0C0F999909280",
 14959 => x"C0C0C0F999909290",
 14960 => x"C0C0C0F9999082C0",
 14961 => x"C0C0C0F9999082F9",
 14962 => x"C0C0C0F9999082A4",
 14963 => x"C0C0C0F9999082B0",
 14964 => x"C0C0C0F999908299",
 14965 => x"C0C0C0F999908292",
 14966 => x"C0C0C0F999908282",
 14967 => x"C0C0C0F9999082F8",
 14968 => x"C0C0C0F999908280",
 14969 => x"C0C0C0F999908290",
 14970 => x"C0C0C0F99990F8C0",
 14971 => x"C0C0C0F99990F8F9",
 14972 => x"C0C0C0F99990F8A4",
 14973 => x"C0C0C0F99990F8B0",
 14974 => x"C0C0C0F99990F899",
 14975 => x"C0C0C0F99990F892",
 14976 => x"C0C0C0F99990F882",
 14977 => x"C0C0C0F99990F8F8",
 14978 => x"C0C0C0F99990F880",
 14979 => x"C0C0C0F99990F890",
 14980 => x"C0C0C0F9999080C0",
 14981 => x"C0C0C0F9999080F9",
 14982 => x"C0C0C0F9999080A4",
 14983 => x"C0C0C0F9999080B0",
 14984 => x"C0C0C0F999908099",
 14985 => x"C0C0C0F999908092",
 14986 => x"C0C0C0F999908082",
 14987 => x"C0C0C0F9999080F8",
 14988 => x"C0C0C0F999908080",
 14989 => x"C0C0C0F999908090",
 14990 => x"C0C0C0F9999090C0",
 14991 => x"C0C0C0F9999090F9",
 14992 => x"C0C0C0F9999090A4",
 14993 => x"C0C0C0F9999090B0",
 14994 => x"C0C0C0F999909099",
 14995 => x"C0C0C0F999909092",
 14996 => x"C0C0C0F999909082",
 14997 => x"C0C0C0F9999090F8",
 14998 => x"C0C0C0F999909080",
 14999 => x"C0C0C0F999909090",
 15000 => x"C0C0C0F992C0C0C0",
 15001 => x"C0C0C0F992C0C0F9",
 15002 => x"C0C0C0F992C0C0A4",
 15003 => x"C0C0C0F992C0C0B0",
 15004 => x"C0C0C0F992C0C099",
 15005 => x"C0C0C0F992C0C092",
 15006 => x"C0C0C0F992C0C082",
 15007 => x"C0C0C0F992C0C0F8",
 15008 => x"C0C0C0F992C0C080",
 15009 => x"C0C0C0F992C0C090",
 15010 => x"C0C0C0F992C0F9C0",
 15011 => x"C0C0C0F992C0F9F9",
 15012 => x"C0C0C0F992C0F9A4",
 15013 => x"C0C0C0F992C0F9B0",
 15014 => x"C0C0C0F992C0F999",
 15015 => x"C0C0C0F992C0F992",
 15016 => x"C0C0C0F992C0F982",
 15017 => x"C0C0C0F992C0F9F8",
 15018 => x"C0C0C0F992C0F980",
 15019 => x"C0C0C0F992C0F990",
 15020 => x"C0C0C0F992C0A4C0",
 15021 => x"C0C0C0F992C0A4F9",
 15022 => x"C0C0C0F992C0A4A4",
 15023 => x"C0C0C0F992C0A4B0",
 15024 => x"C0C0C0F992C0A499",
 15025 => x"C0C0C0F992C0A492",
 15026 => x"C0C0C0F992C0A482",
 15027 => x"C0C0C0F992C0A4F8",
 15028 => x"C0C0C0F992C0A480",
 15029 => x"C0C0C0F992C0A490",
 15030 => x"C0C0C0F992C0B0C0",
 15031 => x"C0C0C0F992C0B0F9",
 15032 => x"C0C0C0F992C0B0A4",
 15033 => x"C0C0C0F992C0B0B0",
 15034 => x"C0C0C0F992C0B099",
 15035 => x"C0C0C0F992C0B092",
 15036 => x"C0C0C0F992C0B082",
 15037 => x"C0C0C0F992C0B0F8",
 15038 => x"C0C0C0F992C0B080",
 15039 => x"C0C0C0F992C0B090",
 15040 => x"C0C0C0F992C099C0",
 15041 => x"C0C0C0F992C099F9",
 15042 => x"C0C0C0F992C099A4",
 15043 => x"C0C0C0F992C099B0",
 15044 => x"C0C0C0F992C09999",
 15045 => x"C0C0C0F992C09992",
 15046 => x"C0C0C0F992C09982",
 15047 => x"C0C0C0F992C099F8",
 15048 => x"C0C0C0F992C09980",
 15049 => x"C0C0C0F992C09990",
 15050 => x"C0C0C0F992C092C0",
 15051 => x"C0C0C0F992C092F9",
 15052 => x"C0C0C0F992C092A4",
 15053 => x"C0C0C0F992C092B0",
 15054 => x"C0C0C0F992C09299",
 15055 => x"C0C0C0F992C09292",
 15056 => x"C0C0C0F992C09282",
 15057 => x"C0C0C0F992C092F8",
 15058 => x"C0C0C0F992C09280",
 15059 => x"C0C0C0F992C09290",
 15060 => x"C0C0C0F992C082C0",
 15061 => x"C0C0C0F992C082F9",
 15062 => x"C0C0C0F992C082A4",
 15063 => x"C0C0C0F992C082B0",
 15064 => x"C0C0C0F992C08299",
 15065 => x"C0C0C0F992C08292",
 15066 => x"C0C0C0F992C08282",
 15067 => x"C0C0C0F992C082F8",
 15068 => x"C0C0C0F992C08280",
 15069 => x"C0C0C0F992C08290",
 15070 => x"C0C0C0F992C0F8C0",
 15071 => x"C0C0C0F992C0F8F9",
 15072 => x"C0C0C0F992C0F8A4",
 15073 => x"C0C0C0F992C0F8B0",
 15074 => x"C0C0C0F992C0F899",
 15075 => x"C0C0C0F992C0F892",
 15076 => x"C0C0C0F992C0F882",
 15077 => x"C0C0C0F992C0F8F8",
 15078 => x"C0C0C0F992C0F880",
 15079 => x"C0C0C0F992C0F890",
 15080 => x"C0C0C0F992C080C0",
 15081 => x"C0C0C0F992C080F9",
 15082 => x"C0C0C0F992C080A4",
 15083 => x"C0C0C0F992C080B0",
 15084 => x"C0C0C0F992C08099",
 15085 => x"C0C0C0F992C08092",
 15086 => x"C0C0C0F992C08082",
 15087 => x"C0C0C0F992C080F8",
 15088 => x"C0C0C0F992C08080",
 15089 => x"C0C0C0F992C08090",
 15090 => x"C0C0C0F992C090C0",
 15091 => x"C0C0C0F992C090F9",
 15092 => x"C0C0C0F992C090A4",
 15093 => x"C0C0C0F992C090B0",
 15094 => x"C0C0C0F992C09099",
 15095 => x"C0C0C0F992C09092",
 15096 => x"C0C0C0F992C09082",
 15097 => x"C0C0C0F992C090F8",
 15098 => x"C0C0C0F992C09080",
 15099 => x"C0C0C0F992C09090",
 15100 => x"C0C0C0F992F9C0C0",
 15101 => x"C0C0C0F992F9C0F9",
 15102 => x"C0C0C0F992F9C0A4",
 15103 => x"C0C0C0F992F9C0B0",
 15104 => x"C0C0C0F992F9C099",
 15105 => x"C0C0C0F992F9C092",
 15106 => x"C0C0C0F992F9C082",
 15107 => x"C0C0C0F992F9C0F8",
 15108 => x"C0C0C0F992F9C080",
 15109 => x"C0C0C0F992F9C090",
 15110 => x"C0C0C0F992F9F9C0",
 15111 => x"C0C0C0F992F9F9F9",
 15112 => x"C0C0C0F992F9F9A4",
 15113 => x"C0C0C0F992F9F9B0",
 15114 => x"C0C0C0F992F9F999",
 15115 => x"C0C0C0F992F9F992",
 15116 => x"C0C0C0F992F9F982",
 15117 => x"C0C0C0F992F9F9F8",
 15118 => x"C0C0C0F992F9F980",
 15119 => x"C0C0C0F992F9F990",
 15120 => x"C0C0C0F992F9A4C0",
 15121 => x"C0C0C0F992F9A4F9",
 15122 => x"C0C0C0F992F9A4A4",
 15123 => x"C0C0C0F992F9A4B0",
 15124 => x"C0C0C0F992F9A499",
 15125 => x"C0C0C0F992F9A492",
 15126 => x"C0C0C0F992F9A482",
 15127 => x"C0C0C0F992F9A4F8",
 15128 => x"C0C0C0F992F9A480",
 15129 => x"C0C0C0F992F9A490",
 15130 => x"C0C0C0F992F9B0C0",
 15131 => x"C0C0C0F992F9B0F9",
 15132 => x"C0C0C0F992F9B0A4",
 15133 => x"C0C0C0F992F9B0B0",
 15134 => x"C0C0C0F992F9B099",
 15135 => x"C0C0C0F992F9B092",
 15136 => x"C0C0C0F992F9B082",
 15137 => x"C0C0C0F992F9B0F8",
 15138 => x"C0C0C0F992F9B080",
 15139 => x"C0C0C0F992F9B090",
 15140 => x"C0C0C0F992F999C0",
 15141 => x"C0C0C0F992F999F9",
 15142 => x"C0C0C0F992F999A4",
 15143 => x"C0C0C0F992F999B0",
 15144 => x"C0C0C0F992F99999",
 15145 => x"C0C0C0F992F99992",
 15146 => x"C0C0C0F992F99982",
 15147 => x"C0C0C0F992F999F8",
 15148 => x"C0C0C0F992F99980",
 15149 => x"C0C0C0F992F99990",
 15150 => x"C0C0C0F992F992C0",
 15151 => x"C0C0C0F992F992F9",
 15152 => x"C0C0C0F992F992A4",
 15153 => x"C0C0C0F992F992B0",
 15154 => x"C0C0C0F992F99299",
 15155 => x"C0C0C0F992F99292",
 15156 => x"C0C0C0F992F99282",
 15157 => x"C0C0C0F992F992F8",
 15158 => x"C0C0C0F992F99280",
 15159 => x"C0C0C0F992F99290",
 15160 => x"C0C0C0F992F982C0",
 15161 => x"C0C0C0F992F982F9",
 15162 => x"C0C0C0F992F982A4",
 15163 => x"C0C0C0F992F982B0",
 15164 => x"C0C0C0F992F98299",
 15165 => x"C0C0C0F992F98292",
 15166 => x"C0C0C0F992F98282",
 15167 => x"C0C0C0F992F982F8",
 15168 => x"C0C0C0F992F98280",
 15169 => x"C0C0C0F992F98290",
 15170 => x"C0C0C0F992F9F8C0",
 15171 => x"C0C0C0F992F9F8F9",
 15172 => x"C0C0C0F992F9F8A4",
 15173 => x"C0C0C0F992F9F8B0",
 15174 => x"C0C0C0F992F9F899",
 15175 => x"C0C0C0F992F9F892",
 15176 => x"C0C0C0F992F9F882",
 15177 => x"C0C0C0F992F9F8F8",
 15178 => x"C0C0C0F992F9F880",
 15179 => x"C0C0C0F992F9F890",
 15180 => x"C0C0C0F992F980C0",
 15181 => x"C0C0C0F992F980F9",
 15182 => x"C0C0C0F992F980A4",
 15183 => x"C0C0C0F992F980B0",
 15184 => x"C0C0C0F992F98099",
 15185 => x"C0C0C0F992F98092",
 15186 => x"C0C0C0F992F98082",
 15187 => x"C0C0C0F992F980F8",
 15188 => x"C0C0C0F992F98080",
 15189 => x"C0C0C0F992F98090",
 15190 => x"C0C0C0F992F990C0",
 15191 => x"C0C0C0F992F990F9",
 15192 => x"C0C0C0F992F990A4",
 15193 => x"C0C0C0F992F990B0",
 15194 => x"C0C0C0F992F99099",
 15195 => x"C0C0C0F992F99092",
 15196 => x"C0C0C0F992F99082",
 15197 => x"C0C0C0F992F990F8",
 15198 => x"C0C0C0F992F99080",
 15199 => x"C0C0C0F992F99090",
 15200 => x"C0C0C0F992A4C0C0",
 15201 => x"C0C0C0F992A4C0F9",
 15202 => x"C0C0C0F992A4C0A4",
 15203 => x"C0C0C0F992A4C0B0",
 15204 => x"C0C0C0F992A4C099",
 15205 => x"C0C0C0F992A4C092",
 15206 => x"C0C0C0F992A4C082",
 15207 => x"C0C0C0F992A4C0F8",
 15208 => x"C0C0C0F992A4C080",
 15209 => x"C0C0C0F992A4C090",
 15210 => x"C0C0C0F992A4F9C0",
 15211 => x"C0C0C0F992A4F9F9",
 15212 => x"C0C0C0F992A4F9A4",
 15213 => x"C0C0C0F992A4F9B0",
 15214 => x"C0C0C0F992A4F999",
 15215 => x"C0C0C0F992A4F992",
 15216 => x"C0C0C0F992A4F982",
 15217 => x"C0C0C0F992A4F9F8",
 15218 => x"C0C0C0F992A4F980",
 15219 => x"C0C0C0F992A4F990",
 15220 => x"C0C0C0F992A4A4C0",
 15221 => x"C0C0C0F992A4A4F9",
 15222 => x"C0C0C0F992A4A4A4",
 15223 => x"C0C0C0F992A4A4B0",
 15224 => x"C0C0C0F992A4A499",
 15225 => x"C0C0C0F992A4A492",
 15226 => x"C0C0C0F992A4A482",
 15227 => x"C0C0C0F992A4A4F8",
 15228 => x"C0C0C0F992A4A480",
 15229 => x"C0C0C0F992A4A490",
 15230 => x"C0C0C0F992A4B0C0",
 15231 => x"C0C0C0F992A4B0F9",
 15232 => x"C0C0C0F992A4B0A4",
 15233 => x"C0C0C0F992A4B0B0",
 15234 => x"C0C0C0F992A4B099",
 15235 => x"C0C0C0F992A4B092",
 15236 => x"C0C0C0F992A4B082",
 15237 => x"C0C0C0F992A4B0F8",
 15238 => x"C0C0C0F992A4B080",
 15239 => x"C0C0C0F992A4B090",
 15240 => x"C0C0C0F992A499C0",
 15241 => x"C0C0C0F992A499F9",
 15242 => x"C0C0C0F992A499A4",
 15243 => x"C0C0C0F992A499B0",
 15244 => x"C0C0C0F992A49999",
 15245 => x"C0C0C0F992A49992",
 15246 => x"C0C0C0F992A49982",
 15247 => x"C0C0C0F992A499F8",
 15248 => x"C0C0C0F992A49980",
 15249 => x"C0C0C0F992A49990",
 15250 => x"C0C0C0F992A492C0",
 15251 => x"C0C0C0F992A492F9",
 15252 => x"C0C0C0F992A492A4",
 15253 => x"C0C0C0F992A492B0",
 15254 => x"C0C0C0F992A49299",
 15255 => x"C0C0C0F992A49292",
 15256 => x"C0C0C0F992A49282",
 15257 => x"C0C0C0F992A492F8",
 15258 => x"C0C0C0F992A49280",
 15259 => x"C0C0C0F992A49290",
 15260 => x"C0C0C0F992A482C0",
 15261 => x"C0C0C0F992A482F9",
 15262 => x"C0C0C0F992A482A4",
 15263 => x"C0C0C0F992A482B0",
 15264 => x"C0C0C0F992A48299",
 15265 => x"C0C0C0F992A48292",
 15266 => x"C0C0C0F992A48282",
 15267 => x"C0C0C0F992A482F8",
 15268 => x"C0C0C0F992A48280",
 15269 => x"C0C0C0F992A48290",
 15270 => x"C0C0C0F992A4F8C0",
 15271 => x"C0C0C0F992A4F8F9",
 15272 => x"C0C0C0F992A4F8A4",
 15273 => x"C0C0C0F992A4F8B0",
 15274 => x"C0C0C0F992A4F899",
 15275 => x"C0C0C0F992A4F892",
 15276 => x"C0C0C0F992A4F882",
 15277 => x"C0C0C0F992A4F8F8",
 15278 => x"C0C0C0F992A4F880",
 15279 => x"C0C0C0F992A4F890",
 15280 => x"C0C0C0F992A480C0",
 15281 => x"C0C0C0F992A480F9",
 15282 => x"C0C0C0F992A480A4",
 15283 => x"C0C0C0F992A480B0",
 15284 => x"C0C0C0F992A48099",
 15285 => x"C0C0C0F992A48092",
 15286 => x"C0C0C0F992A48082",
 15287 => x"C0C0C0F992A480F8",
 15288 => x"C0C0C0F992A48080",
 15289 => x"C0C0C0F992A48090",
 15290 => x"C0C0C0F992A490C0",
 15291 => x"C0C0C0F992A490F9",
 15292 => x"C0C0C0F992A490A4",
 15293 => x"C0C0C0F992A490B0",
 15294 => x"C0C0C0F992A49099",
 15295 => x"C0C0C0F992A49092",
 15296 => x"C0C0C0F992A49082",
 15297 => x"C0C0C0F992A490F8",
 15298 => x"C0C0C0F992A49080",
 15299 => x"C0C0C0F992A49090",
 15300 => x"C0C0C0F992B0C0C0",
 15301 => x"C0C0C0F992B0C0F9",
 15302 => x"C0C0C0F992B0C0A4",
 15303 => x"C0C0C0F992B0C0B0",
 15304 => x"C0C0C0F992B0C099",
 15305 => x"C0C0C0F992B0C092",
 15306 => x"C0C0C0F992B0C082",
 15307 => x"C0C0C0F992B0C0F8",
 15308 => x"C0C0C0F992B0C080",
 15309 => x"C0C0C0F992B0C090",
 15310 => x"C0C0C0F992B0F9C0",
 15311 => x"C0C0C0F992B0F9F9",
 15312 => x"C0C0C0F992B0F9A4",
 15313 => x"C0C0C0F992B0F9B0",
 15314 => x"C0C0C0F992B0F999",
 15315 => x"C0C0C0F992B0F992",
 15316 => x"C0C0C0F992B0F982",
 15317 => x"C0C0C0F992B0F9F8",
 15318 => x"C0C0C0F992B0F980",
 15319 => x"C0C0C0F992B0F990",
 15320 => x"C0C0C0F992B0A4C0",
 15321 => x"C0C0C0F992B0A4F9",
 15322 => x"C0C0C0F992B0A4A4",
 15323 => x"C0C0C0F992B0A4B0",
 15324 => x"C0C0C0F992B0A499",
 15325 => x"C0C0C0F992B0A492",
 15326 => x"C0C0C0F992B0A482",
 15327 => x"C0C0C0F992B0A4F8",
 15328 => x"C0C0C0F992B0A480",
 15329 => x"C0C0C0F992B0A490",
 15330 => x"C0C0C0F992B0B0C0",
 15331 => x"C0C0C0F992B0B0F9",
 15332 => x"C0C0C0F992B0B0A4",
 15333 => x"C0C0C0F992B0B0B0",
 15334 => x"C0C0C0F992B0B099",
 15335 => x"C0C0C0F992B0B092",
 15336 => x"C0C0C0F992B0B082",
 15337 => x"C0C0C0F992B0B0F8",
 15338 => x"C0C0C0F992B0B080",
 15339 => x"C0C0C0F992B0B090",
 15340 => x"C0C0C0F992B099C0",
 15341 => x"C0C0C0F992B099F9",
 15342 => x"C0C0C0F992B099A4",
 15343 => x"C0C0C0F992B099B0",
 15344 => x"C0C0C0F992B09999",
 15345 => x"C0C0C0F992B09992",
 15346 => x"C0C0C0F992B09982",
 15347 => x"C0C0C0F992B099F8",
 15348 => x"C0C0C0F992B09980",
 15349 => x"C0C0C0F992B09990",
 15350 => x"C0C0C0F992B092C0",
 15351 => x"C0C0C0F992B092F9",
 15352 => x"C0C0C0F992B092A4",
 15353 => x"C0C0C0F992B092B0",
 15354 => x"C0C0C0F992B09299",
 15355 => x"C0C0C0F992B09292",
 15356 => x"C0C0C0F992B09282",
 15357 => x"C0C0C0F992B092F8",
 15358 => x"C0C0C0F992B09280",
 15359 => x"C0C0C0F992B09290",
 15360 => x"C0C0C0F992B082C0",
 15361 => x"C0C0C0F992B082F9",
 15362 => x"C0C0C0F992B082A4",
 15363 => x"C0C0C0F992B082B0",
 15364 => x"C0C0C0F992B08299",
 15365 => x"C0C0C0F992B08292",
 15366 => x"C0C0C0F992B08282",
 15367 => x"C0C0C0F992B082F8",
 15368 => x"C0C0C0F992B08280",
 15369 => x"C0C0C0F992B08290",
 15370 => x"C0C0C0F992B0F8C0",
 15371 => x"C0C0C0F992B0F8F9",
 15372 => x"C0C0C0F992B0F8A4",
 15373 => x"C0C0C0F992B0F8B0",
 15374 => x"C0C0C0F992B0F899",
 15375 => x"C0C0C0F992B0F892",
 15376 => x"C0C0C0F992B0F882",
 15377 => x"C0C0C0F992B0F8F8",
 15378 => x"C0C0C0F992B0F880",
 15379 => x"C0C0C0F992B0F890",
 15380 => x"C0C0C0F992B080C0",
 15381 => x"C0C0C0F992B080F9",
 15382 => x"C0C0C0F992B080A4",
 15383 => x"C0C0C0F992B080B0",
 15384 => x"C0C0C0F992B08099",
 15385 => x"C0C0C0F992B08092",
 15386 => x"C0C0C0F992B08082",
 15387 => x"C0C0C0F992B080F8",
 15388 => x"C0C0C0F992B08080",
 15389 => x"C0C0C0F992B08090",
 15390 => x"C0C0C0F992B090C0",
 15391 => x"C0C0C0F992B090F9",
 15392 => x"C0C0C0F992B090A4",
 15393 => x"C0C0C0F992B090B0",
 15394 => x"C0C0C0F992B09099",
 15395 => x"C0C0C0F992B09092",
 15396 => x"C0C0C0F992B09082",
 15397 => x"C0C0C0F992B090F8",
 15398 => x"C0C0C0F992B09080",
 15399 => x"C0C0C0F992B09090",
 15400 => x"C0C0C0F99299C0C0",
 15401 => x"C0C0C0F99299C0F9",
 15402 => x"C0C0C0F99299C0A4",
 15403 => x"C0C0C0F99299C0B0",
 15404 => x"C0C0C0F99299C099",
 15405 => x"C0C0C0F99299C092",
 15406 => x"C0C0C0F99299C082",
 15407 => x"C0C0C0F99299C0F8",
 15408 => x"C0C0C0F99299C080",
 15409 => x"C0C0C0F99299C090",
 15410 => x"C0C0C0F99299F9C0",
 15411 => x"C0C0C0F99299F9F9",
 15412 => x"C0C0C0F99299F9A4",
 15413 => x"C0C0C0F99299F9B0",
 15414 => x"C0C0C0F99299F999",
 15415 => x"C0C0C0F99299F992",
 15416 => x"C0C0C0F99299F982",
 15417 => x"C0C0C0F99299F9F8",
 15418 => x"C0C0C0F99299F980",
 15419 => x"C0C0C0F99299F990",
 15420 => x"C0C0C0F99299A4C0",
 15421 => x"C0C0C0F99299A4F9",
 15422 => x"C0C0C0F99299A4A4",
 15423 => x"C0C0C0F99299A4B0",
 15424 => x"C0C0C0F99299A499",
 15425 => x"C0C0C0F99299A492",
 15426 => x"C0C0C0F99299A482",
 15427 => x"C0C0C0F99299A4F8",
 15428 => x"C0C0C0F99299A480",
 15429 => x"C0C0C0F99299A490",
 15430 => x"C0C0C0F99299B0C0",
 15431 => x"C0C0C0F99299B0F9",
 15432 => x"C0C0C0F99299B0A4",
 15433 => x"C0C0C0F99299B0B0",
 15434 => x"C0C0C0F99299B099",
 15435 => x"C0C0C0F99299B092",
 15436 => x"C0C0C0F99299B082",
 15437 => x"C0C0C0F99299B0F8",
 15438 => x"C0C0C0F99299B080",
 15439 => x"C0C0C0F99299B090",
 15440 => x"C0C0C0F9929999C0",
 15441 => x"C0C0C0F9929999F9",
 15442 => x"C0C0C0F9929999A4",
 15443 => x"C0C0C0F9929999B0",
 15444 => x"C0C0C0F992999999",
 15445 => x"C0C0C0F992999992",
 15446 => x"C0C0C0F992999982",
 15447 => x"C0C0C0F9929999F8",
 15448 => x"C0C0C0F992999980",
 15449 => x"C0C0C0F992999990",
 15450 => x"C0C0C0F9929992C0",
 15451 => x"C0C0C0F9929992F9",
 15452 => x"C0C0C0F9929992A4",
 15453 => x"C0C0C0F9929992B0",
 15454 => x"C0C0C0F992999299",
 15455 => x"C0C0C0F992999292",
 15456 => x"C0C0C0F992999282",
 15457 => x"C0C0C0F9929992F8",
 15458 => x"C0C0C0F992999280",
 15459 => x"C0C0C0F992999290",
 15460 => x"C0C0C0F9929982C0",
 15461 => x"C0C0C0F9929982F9",
 15462 => x"C0C0C0F9929982A4",
 15463 => x"C0C0C0F9929982B0",
 15464 => x"C0C0C0F992998299",
 15465 => x"C0C0C0F992998292",
 15466 => x"C0C0C0F992998282",
 15467 => x"C0C0C0F9929982F8",
 15468 => x"C0C0C0F992998280",
 15469 => x"C0C0C0F992998290",
 15470 => x"C0C0C0F99299F8C0",
 15471 => x"C0C0C0F99299F8F9",
 15472 => x"C0C0C0F99299F8A4",
 15473 => x"C0C0C0F99299F8B0",
 15474 => x"C0C0C0F99299F899",
 15475 => x"C0C0C0F99299F892",
 15476 => x"C0C0C0F99299F882",
 15477 => x"C0C0C0F99299F8F8",
 15478 => x"C0C0C0F99299F880",
 15479 => x"C0C0C0F99299F890",
 15480 => x"C0C0C0F9929980C0",
 15481 => x"C0C0C0F9929980F9",
 15482 => x"C0C0C0F9929980A4",
 15483 => x"C0C0C0F9929980B0",
 15484 => x"C0C0C0F992998099",
 15485 => x"C0C0C0F992998092",
 15486 => x"C0C0C0F992998082",
 15487 => x"C0C0C0F9929980F8",
 15488 => x"C0C0C0F992998080",
 15489 => x"C0C0C0F992998090",
 15490 => x"C0C0C0F9929990C0",
 15491 => x"C0C0C0F9929990F9",
 15492 => x"C0C0C0F9929990A4",
 15493 => x"C0C0C0F9929990B0",
 15494 => x"C0C0C0F992999099",
 15495 => x"C0C0C0F992999092",
 15496 => x"C0C0C0F992999082",
 15497 => x"C0C0C0F9929990F8",
 15498 => x"C0C0C0F992999080",
 15499 => x"C0C0C0F992999090",
 15500 => x"C0C0C0F99292C0C0",
 15501 => x"C0C0C0F99292C0F9",
 15502 => x"C0C0C0F99292C0A4",
 15503 => x"C0C0C0F99292C0B0",
 15504 => x"C0C0C0F99292C099",
 15505 => x"C0C0C0F99292C092",
 15506 => x"C0C0C0F99292C082",
 15507 => x"C0C0C0F99292C0F8",
 15508 => x"C0C0C0F99292C080",
 15509 => x"C0C0C0F99292C090",
 15510 => x"C0C0C0F99292F9C0",
 15511 => x"C0C0C0F99292F9F9",
 15512 => x"C0C0C0F99292F9A4",
 15513 => x"C0C0C0F99292F9B0",
 15514 => x"C0C0C0F99292F999",
 15515 => x"C0C0C0F99292F992",
 15516 => x"C0C0C0F99292F982",
 15517 => x"C0C0C0F99292F9F8",
 15518 => x"C0C0C0F99292F980",
 15519 => x"C0C0C0F99292F990",
 15520 => x"C0C0C0F99292A4C0",
 15521 => x"C0C0C0F99292A4F9",
 15522 => x"C0C0C0F99292A4A4",
 15523 => x"C0C0C0F99292A4B0",
 15524 => x"C0C0C0F99292A499",
 15525 => x"C0C0C0F99292A492",
 15526 => x"C0C0C0F99292A482",
 15527 => x"C0C0C0F99292A4F8",
 15528 => x"C0C0C0F99292A480",
 15529 => x"C0C0C0F99292A490",
 15530 => x"C0C0C0F99292B0C0",
 15531 => x"C0C0C0F99292B0F9",
 15532 => x"C0C0C0F99292B0A4",
 15533 => x"C0C0C0F99292B0B0",
 15534 => x"C0C0C0F99292B099",
 15535 => x"C0C0C0F99292B092",
 15536 => x"C0C0C0F99292B082",
 15537 => x"C0C0C0F99292B0F8",
 15538 => x"C0C0C0F99292B080",
 15539 => x"C0C0C0F99292B090",
 15540 => x"C0C0C0F9929299C0",
 15541 => x"C0C0C0F9929299F9",
 15542 => x"C0C0C0F9929299A4",
 15543 => x"C0C0C0F9929299B0",
 15544 => x"C0C0C0F992929999",
 15545 => x"C0C0C0F992929992",
 15546 => x"C0C0C0F992929982",
 15547 => x"C0C0C0F9929299F8",
 15548 => x"C0C0C0F992929980",
 15549 => x"C0C0C0F992929990",
 15550 => x"C0C0C0F9929292C0",
 15551 => x"C0C0C0F9929292F9",
 15552 => x"C0C0C0F9929292A4",
 15553 => x"C0C0C0F9929292B0",
 15554 => x"C0C0C0F992929299",
 15555 => x"C0C0C0F992929292",
 15556 => x"C0C0C0F992929282",
 15557 => x"C0C0C0F9929292F8",
 15558 => x"C0C0C0F992929280",
 15559 => x"C0C0C0F992929290",
 15560 => x"C0C0C0F9929282C0",
 15561 => x"C0C0C0F9929282F9",
 15562 => x"C0C0C0F9929282A4",
 15563 => x"C0C0C0F9929282B0",
 15564 => x"C0C0C0F992928299",
 15565 => x"C0C0C0F992928292",
 15566 => x"C0C0C0F992928282",
 15567 => x"C0C0C0F9929282F8",
 15568 => x"C0C0C0F992928280",
 15569 => x"C0C0C0F992928290",
 15570 => x"C0C0C0F99292F8C0",
 15571 => x"C0C0C0F99292F8F9",
 15572 => x"C0C0C0F99292F8A4",
 15573 => x"C0C0C0F99292F8B0",
 15574 => x"C0C0C0F99292F899",
 15575 => x"C0C0C0F99292F892",
 15576 => x"C0C0C0F99292F882",
 15577 => x"C0C0C0F99292F8F8",
 15578 => x"C0C0C0F99292F880",
 15579 => x"C0C0C0F99292F890",
 15580 => x"C0C0C0F9929280C0",
 15581 => x"C0C0C0F9929280F9",
 15582 => x"C0C0C0F9929280A4",
 15583 => x"C0C0C0F9929280B0",
 15584 => x"C0C0C0F992928099",
 15585 => x"C0C0C0F992928092",
 15586 => x"C0C0C0F992928082",
 15587 => x"C0C0C0F9929280F8",
 15588 => x"C0C0C0F992928080",
 15589 => x"C0C0C0F992928090",
 15590 => x"C0C0C0F9929290C0",
 15591 => x"C0C0C0F9929290F9",
 15592 => x"C0C0C0F9929290A4",
 15593 => x"C0C0C0F9929290B0",
 15594 => x"C0C0C0F992929099",
 15595 => x"C0C0C0F992929092",
 15596 => x"C0C0C0F992929082",
 15597 => x"C0C0C0F9929290F8",
 15598 => x"C0C0C0F992929080",
 15599 => x"C0C0C0F992929090",
 15600 => x"C0C0C0F99282C0C0",
 15601 => x"C0C0C0F99282C0F9",
 15602 => x"C0C0C0F99282C0A4",
 15603 => x"C0C0C0F99282C0B0",
 15604 => x"C0C0C0F99282C099",
 15605 => x"C0C0C0F99282C092",
 15606 => x"C0C0C0F99282C082",
 15607 => x"C0C0C0F99282C0F8",
 15608 => x"C0C0C0F99282C080",
 15609 => x"C0C0C0F99282C090",
 15610 => x"C0C0C0F99282F9C0",
 15611 => x"C0C0C0F99282F9F9",
 15612 => x"C0C0C0F99282F9A4",
 15613 => x"C0C0C0F99282F9B0",
 15614 => x"C0C0C0F99282F999",
 15615 => x"C0C0C0F99282F992",
 15616 => x"C0C0C0F99282F982",
 15617 => x"C0C0C0F99282F9F8",
 15618 => x"C0C0C0F99282F980",
 15619 => x"C0C0C0F99282F990",
 15620 => x"C0C0C0F99282A4C0",
 15621 => x"C0C0C0F99282A4F9",
 15622 => x"C0C0C0F99282A4A4",
 15623 => x"C0C0C0F99282A4B0",
 15624 => x"C0C0C0F99282A499",
 15625 => x"C0C0C0F99282A492",
 15626 => x"C0C0C0F99282A482",
 15627 => x"C0C0C0F99282A4F8",
 15628 => x"C0C0C0F99282A480",
 15629 => x"C0C0C0F99282A490",
 15630 => x"C0C0C0F99282B0C0",
 15631 => x"C0C0C0F99282B0F9",
 15632 => x"C0C0C0F99282B0A4",
 15633 => x"C0C0C0F99282B0B0",
 15634 => x"C0C0C0F99282B099",
 15635 => x"C0C0C0F99282B092",
 15636 => x"C0C0C0F99282B082",
 15637 => x"C0C0C0F99282B0F8",
 15638 => x"C0C0C0F99282B080",
 15639 => x"C0C0C0F99282B090",
 15640 => x"C0C0C0F9928299C0",
 15641 => x"C0C0C0F9928299F9",
 15642 => x"C0C0C0F9928299A4",
 15643 => x"C0C0C0F9928299B0",
 15644 => x"C0C0C0F992829999",
 15645 => x"C0C0C0F992829992",
 15646 => x"C0C0C0F992829982",
 15647 => x"C0C0C0F9928299F8",
 15648 => x"C0C0C0F992829980",
 15649 => x"C0C0C0F992829990",
 15650 => x"C0C0C0F9928292C0",
 15651 => x"C0C0C0F9928292F9",
 15652 => x"C0C0C0F9928292A4",
 15653 => x"C0C0C0F9928292B0",
 15654 => x"C0C0C0F992829299",
 15655 => x"C0C0C0F992829292",
 15656 => x"C0C0C0F992829282",
 15657 => x"C0C0C0F9928292F8",
 15658 => x"C0C0C0F992829280",
 15659 => x"C0C0C0F992829290",
 15660 => x"C0C0C0F9928282C0",
 15661 => x"C0C0C0F9928282F9",
 15662 => x"C0C0C0F9928282A4",
 15663 => x"C0C0C0F9928282B0",
 15664 => x"C0C0C0F992828299",
 15665 => x"C0C0C0F992828292",
 15666 => x"C0C0C0F992828282",
 15667 => x"C0C0C0F9928282F8",
 15668 => x"C0C0C0F992828280",
 15669 => x"C0C0C0F992828290",
 15670 => x"C0C0C0F99282F8C0",
 15671 => x"C0C0C0F99282F8F9",
 15672 => x"C0C0C0F99282F8A4",
 15673 => x"C0C0C0F99282F8B0",
 15674 => x"C0C0C0F99282F899",
 15675 => x"C0C0C0F99282F892",
 15676 => x"C0C0C0F99282F882",
 15677 => x"C0C0C0F99282F8F8",
 15678 => x"C0C0C0F99282F880",
 15679 => x"C0C0C0F99282F890",
 15680 => x"C0C0C0F9928280C0",
 15681 => x"C0C0C0F9928280F9",
 15682 => x"C0C0C0F9928280A4",
 15683 => x"C0C0C0F9928280B0",
 15684 => x"C0C0C0F992828099",
 15685 => x"C0C0C0F992828092",
 15686 => x"C0C0C0F992828082",
 15687 => x"C0C0C0F9928280F8",
 15688 => x"C0C0C0F992828080",
 15689 => x"C0C0C0F992828090",
 15690 => x"C0C0C0F9928290C0",
 15691 => x"C0C0C0F9928290F9",
 15692 => x"C0C0C0F9928290A4",
 15693 => x"C0C0C0F9928290B0",
 15694 => x"C0C0C0F992829099",
 15695 => x"C0C0C0F992829092",
 15696 => x"C0C0C0F992829082",
 15697 => x"C0C0C0F9928290F8",
 15698 => x"C0C0C0F992829080",
 15699 => x"C0C0C0F992829090",
 15700 => x"C0C0C0F992F8C0C0",
 15701 => x"C0C0C0F992F8C0F9",
 15702 => x"C0C0C0F992F8C0A4",
 15703 => x"C0C0C0F992F8C0B0",
 15704 => x"C0C0C0F992F8C099",
 15705 => x"C0C0C0F992F8C092",
 15706 => x"C0C0C0F992F8C082",
 15707 => x"C0C0C0F992F8C0F8",
 15708 => x"C0C0C0F992F8C080",
 15709 => x"C0C0C0F992F8C090",
 15710 => x"C0C0C0F992F8F9C0",
 15711 => x"C0C0C0F992F8F9F9",
 15712 => x"C0C0C0F992F8F9A4",
 15713 => x"C0C0C0F992F8F9B0",
 15714 => x"C0C0C0F992F8F999",
 15715 => x"C0C0C0F992F8F992",
 15716 => x"C0C0C0F992F8F982",
 15717 => x"C0C0C0F992F8F9F8",
 15718 => x"C0C0C0F992F8F980",
 15719 => x"C0C0C0F992F8F990",
 15720 => x"C0C0C0F992F8A4C0",
 15721 => x"C0C0C0F992F8A4F9",
 15722 => x"C0C0C0F992F8A4A4",
 15723 => x"C0C0C0F992F8A4B0",
 15724 => x"C0C0C0F992F8A499",
 15725 => x"C0C0C0F992F8A492",
 15726 => x"C0C0C0F992F8A482",
 15727 => x"C0C0C0F992F8A4F8",
 15728 => x"C0C0C0F992F8A480",
 15729 => x"C0C0C0F992F8A490",
 15730 => x"C0C0C0F992F8B0C0",
 15731 => x"C0C0C0F992F8B0F9",
 15732 => x"C0C0C0F992F8B0A4",
 15733 => x"C0C0C0F992F8B0B0",
 15734 => x"C0C0C0F992F8B099",
 15735 => x"C0C0C0F992F8B092",
 15736 => x"C0C0C0F992F8B082",
 15737 => x"C0C0C0F992F8B0F8",
 15738 => x"C0C0C0F992F8B080",
 15739 => x"C0C0C0F992F8B090",
 15740 => x"C0C0C0F992F899C0",
 15741 => x"C0C0C0F992F899F9",
 15742 => x"C0C0C0F992F899A4",
 15743 => x"C0C0C0F992F899B0",
 15744 => x"C0C0C0F992F89999",
 15745 => x"C0C0C0F992F89992",
 15746 => x"C0C0C0F992F89982",
 15747 => x"C0C0C0F992F899F8",
 15748 => x"C0C0C0F992F89980",
 15749 => x"C0C0C0F992F89990",
 15750 => x"C0C0C0F992F892C0",
 15751 => x"C0C0C0F992F892F9",
 15752 => x"C0C0C0F992F892A4",
 15753 => x"C0C0C0F992F892B0",
 15754 => x"C0C0C0F992F89299",
 15755 => x"C0C0C0F992F89292",
 15756 => x"C0C0C0F992F89282",
 15757 => x"C0C0C0F992F892F8",
 15758 => x"C0C0C0F992F89280",
 15759 => x"C0C0C0F992F89290",
 15760 => x"C0C0C0F992F882C0",
 15761 => x"C0C0C0F992F882F9",
 15762 => x"C0C0C0F992F882A4",
 15763 => x"C0C0C0F992F882B0",
 15764 => x"C0C0C0F992F88299",
 15765 => x"C0C0C0F992F88292",
 15766 => x"C0C0C0F992F88282",
 15767 => x"C0C0C0F992F882F8",
 15768 => x"C0C0C0F992F88280",
 15769 => x"C0C0C0F992F88290",
 15770 => x"C0C0C0F992F8F8C0",
 15771 => x"C0C0C0F992F8F8F9",
 15772 => x"C0C0C0F992F8F8A4",
 15773 => x"C0C0C0F992F8F8B0",
 15774 => x"C0C0C0F992F8F899",
 15775 => x"C0C0C0F992F8F892",
 15776 => x"C0C0C0F992F8F882",
 15777 => x"C0C0C0F992F8F8F8",
 15778 => x"C0C0C0F992F8F880",
 15779 => x"C0C0C0F992F8F890",
 15780 => x"C0C0C0F992F880C0",
 15781 => x"C0C0C0F992F880F9",
 15782 => x"C0C0C0F992F880A4",
 15783 => x"C0C0C0F992F880B0",
 15784 => x"C0C0C0F992F88099",
 15785 => x"C0C0C0F992F88092",
 15786 => x"C0C0C0F992F88082",
 15787 => x"C0C0C0F992F880F8",
 15788 => x"C0C0C0F992F88080",
 15789 => x"C0C0C0F992F88090",
 15790 => x"C0C0C0F992F890C0",
 15791 => x"C0C0C0F992F890F9",
 15792 => x"C0C0C0F992F890A4",
 15793 => x"C0C0C0F992F890B0",
 15794 => x"C0C0C0F992F89099",
 15795 => x"C0C0C0F992F89092",
 15796 => x"C0C0C0F992F89082",
 15797 => x"C0C0C0F992F890F8",
 15798 => x"C0C0C0F992F89080",
 15799 => x"C0C0C0F992F89090",
 15800 => x"C0C0C0F99280C0C0",
 15801 => x"C0C0C0F99280C0F9",
 15802 => x"C0C0C0F99280C0A4",
 15803 => x"C0C0C0F99280C0B0",
 15804 => x"C0C0C0F99280C099",
 15805 => x"C0C0C0F99280C092",
 15806 => x"C0C0C0F99280C082",
 15807 => x"C0C0C0F99280C0F8",
 15808 => x"C0C0C0F99280C080",
 15809 => x"C0C0C0F99280C090",
 15810 => x"C0C0C0F99280F9C0",
 15811 => x"C0C0C0F99280F9F9",
 15812 => x"C0C0C0F99280F9A4",
 15813 => x"C0C0C0F99280F9B0",
 15814 => x"C0C0C0F99280F999",
 15815 => x"C0C0C0F99280F992",
 15816 => x"C0C0C0F99280F982",
 15817 => x"C0C0C0F99280F9F8",
 15818 => x"C0C0C0F99280F980",
 15819 => x"C0C0C0F99280F990",
 15820 => x"C0C0C0F99280A4C0",
 15821 => x"C0C0C0F99280A4F9",
 15822 => x"C0C0C0F99280A4A4",
 15823 => x"C0C0C0F99280A4B0",
 15824 => x"C0C0C0F99280A499",
 15825 => x"C0C0C0F99280A492",
 15826 => x"C0C0C0F99280A482",
 15827 => x"C0C0C0F99280A4F8",
 15828 => x"C0C0C0F99280A480",
 15829 => x"C0C0C0F99280A490",
 15830 => x"C0C0C0F99280B0C0",
 15831 => x"C0C0C0F99280B0F9",
 15832 => x"C0C0C0F99280B0A4",
 15833 => x"C0C0C0F99280B0B0",
 15834 => x"C0C0C0F99280B099",
 15835 => x"C0C0C0F99280B092",
 15836 => x"C0C0C0F99280B082",
 15837 => x"C0C0C0F99280B0F8",
 15838 => x"C0C0C0F99280B080",
 15839 => x"C0C0C0F99280B090",
 15840 => x"C0C0C0F9928099C0",
 15841 => x"C0C0C0F9928099F9",
 15842 => x"C0C0C0F9928099A4",
 15843 => x"C0C0C0F9928099B0",
 15844 => x"C0C0C0F992809999",
 15845 => x"C0C0C0F992809992",
 15846 => x"C0C0C0F992809982",
 15847 => x"C0C0C0F9928099F8",
 15848 => x"C0C0C0F992809980",
 15849 => x"C0C0C0F992809990",
 15850 => x"C0C0C0F9928092C0",
 15851 => x"C0C0C0F9928092F9",
 15852 => x"C0C0C0F9928092A4",
 15853 => x"C0C0C0F9928092B0",
 15854 => x"C0C0C0F992809299",
 15855 => x"C0C0C0F992809292",
 15856 => x"C0C0C0F992809282",
 15857 => x"C0C0C0F9928092F8",
 15858 => x"C0C0C0F992809280",
 15859 => x"C0C0C0F992809290",
 15860 => x"C0C0C0F9928082C0",
 15861 => x"C0C0C0F9928082F9",
 15862 => x"C0C0C0F9928082A4",
 15863 => x"C0C0C0F9928082B0",
 15864 => x"C0C0C0F992808299",
 15865 => x"C0C0C0F992808292",
 15866 => x"C0C0C0F992808282",
 15867 => x"C0C0C0F9928082F8",
 15868 => x"C0C0C0F992808280",
 15869 => x"C0C0C0F992808290",
 15870 => x"C0C0C0F99280F8C0",
 15871 => x"C0C0C0F99280F8F9",
 15872 => x"C0C0C0F99280F8A4",
 15873 => x"C0C0C0F99280F8B0",
 15874 => x"C0C0C0F99280F899",
 15875 => x"C0C0C0F99280F892",
 15876 => x"C0C0C0F99280F882",
 15877 => x"C0C0C0F99280F8F8",
 15878 => x"C0C0C0F99280F880",
 15879 => x"C0C0C0F99280F890",
 15880 => x"C0C0C0F9928080C0",
 15881 => x"C0C0C0F9928080F9",
 15882 => x"C0C0C0F9928080A4",
 15883 => x"C0C0C0F9928080B0",
 15884 => x"C0C0C0F992808099",
 15885 => x"C0C0C0F992808092",
 15886 => x"C0C0C0F992808082",
 15887 => x"C0C0C0F9928080F8",
 15888 => x"C0C0C0F992808080",
 15889 => x"C0C0C0F992808090",
 15890 => x"C0C0C0F9928090C0",
 15891 => x"C0C0C0F9928090F9",
 15892 => x"C0C0C0F9928090A4",
 15893 => x"C0C0C0F9928090B0",
 15894 => x"C0C0C0F992809099",
 15895 => x"C0C0C0F992809092",
 15896 => x"C0C0C0F992809082",
 15897 => x"C0C0C0F9928090F8",
 15898 => x"C0C0C0F992809080",
 15899 => x"C0C0C0F992809090",
 15900 => x"C0C0C0F99290C0C0",
 15901 => x"C0C0C0F99290C0F9",
 15902 => x"C0C0C0F99290C0A4",
 15903 => x"C0C0C0F99290C0B0",
 15904 => x"C0C0C0F99290C099",
 15905 => x"C0C0C0F99290C092",
 15906 => x"C0C0C0F99290C082",
 15907 => x"C0C0C0F99290C0F8",
 15908 => x"C0C0C0F99290C080",
 15909 => x"C0C0C0F99290C090",
 15910 => x"C0C0C0F99290F9C0",
 15911 => x"C0C0C0F99290F9F9",
 15912 => x"C0C0C0F99290F9A4",
 15913 => x"C0C0C0F99290F9B0",
 15914 => x"C0C0C0F99290F999",
 15915 => x"C0C0C0F99290F992",
 15916 => x"C0C0C0F99290F982",
 15917 => x"C0C0C0F99290F9F8",
 15918 => x"C0C0C0F99290F980",
 15919 => x"C0C0C0F99290F990",
 15920 => x"C0C0C0F99290A4C0",
 15921 => x"C0C0C0F99290A4F9",
 15922 => x"C0C0C0F99290A4A4",
 15923 => x"C0C0C0F99290A4B0",
 15924 => x"C0C0C0F99290A499",
 15925 => x"C0C0C0F99290A492",
 15926 => x"C0C0C0F99290A482",
 15927 => x"C0C0C0F99290A4F8",
 15928 => x"C0C0C0F99290A480",
 15929 => x"C0C0C0F99290A490",
 15930 => x"C0C0C0F99290B0C0",
 15931 => x"C0C0C0F99290B0F9",
 15932 => x"C0C0C0F99290B0A4",
 15933 => x"C0C0C0F99290B0B0",
 15934 => x"C0C0C0F99290B099",
 15935 => x"C0C0C0F99290B092",
 15936 => x"C0C0C0F99290B082",
 15937 => x"C0C0C0F99290B0F8",
 15938 => x"C0C0C0F99290B080",
 15939 => x"C0C0C0F99290B090",
 15940 => x"C0C0C0F9929099C0",
 15941 => x"C0C0C0F9929099F9",
 15942 => x"C0C0C0F9929099A4",
 15943 => x"C0C0C0F9929099B0",
 15944 => x"C0C0C0F992909999",
 15945 => x"C0C0C0F992909992",
 15946 => x"C0C0C0F992909982",
 15947 => x"C0C0C0F9929099F8",
 15948 => x"C0C0C0F992909980",
 15949 => x"C0C0C0F992909990",
 15950 => x"C0C0C0F9929092C0",
 15951 => x"C0C0C0F9929092F9",
 15952 => x"C0C0C0F9929092A4",
 15953 => x"C0C0C0F9929092B0",
 15954 => x"C0C0C0F992909299",
 15955 => x"C0C0C0F992909292",
 15956 => x"C0C0C0F992909282",
 15957 => x"C0C0C0F9929092F8",
 15958 => x"C0C0C0F992909280",
 15959 => x"C0C0C0F992909290",
 15960 => x"C0C0C0F9929082C0",
 15961 => x"C0C0C0F9929082F9",
 15962 => x"C0C0C0F9929082A4",
 15963 => x"C0C0C0F9929082B0",
 15964 => x"C0C0C0F992908299",
 15965 => x"C0C0C0F992908292",
 15966 => x"C0C0C0F992908282",
 15967 => x"C0C0C0F9929082F8",
 15968 => x"C0C0C0F992908280",
 15969 => x"C0C0C0F992908290",
 15970 => x"C0C0C0F99290F8C0",
 15971 => x"C0C0C0F99290F8F9",
 15972 => x"C0C0C0F99290F8A4",
 15973 => x"C0C0C0F99290F8B0",
 15974 => x"C0C0C0F99290F899",
 15975 => x"C0C0C0F99290F892",
 15976 => x"C0C0C0F99290F882",
 15977 => x"C0C0C0F99290F8F8",
 15978 => x"C0C0C0F99290F880",
 15979 => x"C0C0C0F99290F890",
 15980 => x"C0C0C0F9929080C0",
 15981 => x"C0C0C0F9929080F9",
 15982 => x"C0C0C0F9929080A4",
 15983 => x"C0C0C0F9929080B0",
 15984 => x"C0C0C0F992908099",
 15985 => x"C0C0C0F992908092",
 15986 => x"C0C0C0F992908082",
 15987 => x"C0C0C0F9929080F8",
 15988 => x"C0C0C0F992908080",
 15989 => x"C0C0C0F992908090",
 15990 => x"C0C0C0F9929090C0",
 15991 => x"C0C0C0F9929090F9",
 15992 => x"C0C0C0F9929090A4",
 15993 => x"C0C0C0F9929090B0",
 15994 => x"C0C0C0F992909099",
 15995 => x"C0C0C0F992909092",
 15996 => x"C0C0C0F992909082",
 15997 => x"C0C0C0F9929090F8",
 15998 => x"C0C0C0F992909080",
 15999 => x"C0C0C0F992909090",
 16000 => x"C0C0C0F982C0C0C0",
 16001 => x"C0C0C0F982C0C0F9",
 16002 => x"C0C0C0F982C0C0A4",
 16003 => x"C0C0C0F982C0C0B0",
 16004 => x"C0C0C0F982C0C099",
 16005 => x"C0C0C0F982C0C092",
 16006 => x"C0C0C0F982C0C082",
 16007 => x"C0C0C0F982C0C0F8",
 16008 => x"C0C0C0F982C0C080",
 16009 => x"C0C0C0F982C0C090",
 16010 => x"C0C0C0F982C0F9C0",
 16011 => x"C0C0C0F982C0F9F9",
 16012 => x"C0C0C0F982C0F9A4",
 16013 => x"C0C0C0F982C0F9B0",
 16014 => x"C0C0C0F982C0F999",
 16015 => x"C0C0C0F982C0F992",
 16016 => x"C0C0C0F982C0F982",
 16017 => x"C0C0C0F982C0F9F8",
 16018 => x"C0C0C0F982C0F980",
 16019 => x"C0C0C0F982C0F990",
 16020 => x"C0C0C0F982C0A4C0",
 16021 => x"C0C0C0F982C0A4F9",
 16022 => x"C0C0C0F982C0A4A4",
 16023 => x"C0C0C0F982C0A4B0",
 16024 => x"C0C0C0F982C0A499",
 16025 => x"C0C0C0F982C0A492",
 16026 => x"C0C0C0F982C0A482",
 16027 => x"C0C0C0F982C0A4F8",
 16028 => x"C0C0C0F982C0A480",
 16029 => x"C0C0C0F982C0A490",
 16030 => x"C0C0C0F982C0B0C0",
 16031 => x"C0C0C0F982C0B0F9",
 16032 => x"C0C0C0F982C0B0A4",
 16033 => x"C0C0C0F982C0B0B0",
 16034 => x"C0C0C0F982C0B099",
 16035 => x"C0C0C0F982C0B092",
 16036 => x"C0C0C0F982C0B082",
 16037 => x"C0C0C0F982C0B0F8",
 16038 => x"C0C0C0F982C0B080",
 16039 => x"C0C0C0F982C0B090",
 16040 => x"C0C0C0F982C099C0",
 16041 => x"C0C0C0F982C099F9",
 16042 => x"C0C0C0F982C099A4",
 16043 => x"C0C0C0F982C099B0",
 16044 => x"C0C0C0F982C09999",
 16045 => x"C0C0C0F982C09992",
 16046 => x"C0C0C0F982C09982",
 16047 => x"C0C0C0F982C099F8",
 16048 => x"C0C0C0F982C09980",
 16049 => x"C0C0C0F982C09990",
 16050 => x"C0C0C0F982C092C0",
 16051 => x"C0C0C0F982C092F9",
 16052 => x"C0C0C0F982C092A4",
 16053 => x"C0C0C0F982C092B0",
 16054 => x"C0C0C0F982C09299",
 16055 => x"C0C0C0F982C09292",
 16056 => x"C0C0C0F982C09282",
 16057 => x"C0C0C0F982C092F8",
 16058 => x"C0C0C0F982C09280",
 16059 => x"C0C0C0F982C09290",
 16060 => x"C0C0C0F982C082C0",
 16061 => x"C0C0C0F982C082F9",
 16062 => x"C0C0C0F982C082A4",
 16063 => x"C0C0C0F982C082B0",
 16064 => x"C0C0C0F982C08299",
 16065 => x"C0C0C0F982C08292",
 16066 => x"C0C0C0F982C08282",
 16067 => x"C0C0C0F982C082F8",
 16068 => x"C0C0C0F982C08280",
 16069 => x"C0C0C0F982C08290",
 16070 => x"C0C0C0F982C0F8C0",
 16071 => x"C0C0C0F982C0F8F9",
 16072 => x"C0C0C0F982C0F8A4",
 16073 => x"C0C0C0F982C0F8B0",
 16074 => x"C0C0C0F982C0F899",
 16075 => x"C0C0C0F982C0F892",
 16076 => x"C0C0C0F982C0F882",
 16077 => x"C0C0C0F982C0F8F8",
 16078 => x"C0C0C0F982C0F880",
 16079 => x"C0C0C0F982C0F890",
 16080 => x"C0C0C0F982C080C0",
 16081 => x"C0C0C0F982C080F9",
 16082 => x"C0C0C0F982C080A4",
 16083 => x"C0C0C0F982C080B0",
 16084 => x"C0C0C0F982C08099",
 16085 => x"C0C0C0F982C08092",
 16086 => x"C0C0C0F982C08082",
 16087 => x"C0C0C0F982C080F8",
 16088 => x"C0C0C0F982C08080",
 16089 => x"C0C0C0F982C08090",
 16090 => x"C0C0C0F982C090C0",
 16091 => x"C0C0C0F982C090F9",
 16092 => x"C0C0C0F982C090A4",
 16093 => x"C0C0C0F982C090B0",
 16094 => x"C0C0C0F982C09099",
 16095 => x"C0C0C0F982C09092",
 16096 => x"C0C0C0F982C09082",
 16097 => x"C0C0C0F982C090F8",
 16098 => x"C0C0C0F982C09080",
 16099 => x"C0C0C0F982C09090",
 16100 => x"C0C0C0F982F9C0C0",
 16101 => x"C0C0C0F982F9C0F9",
 16102 => x"C0C0C0F982F9C0A4",
 16103 => x"C0C0C0F982F9C0B0",
 16104 => x"C0C0C0F982F9C099",
 16105 => x"C0C0C0F982F9C092",
 16106 => x"C0C0C0F982F9C082",
 16107 => x"C0C0C0F982F9C0F8",
 16108 => x"C0C0C0F982F9C080",
 16109 => x"C0C0C0F982F9C090",
 16110 => x"C0C0C0F982F9F9C0",
 16111 => x"C0C0C0F982F9F9F9",
 16112 => x"C0C0C0F982F9F9A4",
 16113 => x"C0C0C0F982F9F9B0",
 16114 => x"C0C0C0F982F9F999",
 16115 => x"C0C0C0F982F9F992",
 16116 => x"C0C0C0F982F9F982",
 16117 => x"C0C0C0F982F9F9F8",
 16118 => x"C0C0C0F982F9F980",
 16119 => x"C0C0C0F982F9F990",
 16120 => x"C0C0C0F982F9A4C0",
 16121 => x"C0C0C0F982F9A4F9",
 16122 => x"C0C0C0F982F9A4A4",
 16123 => x"C0C0C0F982F9A4B0",
 16124 => x"C0C0C0F982F9A499",
 16125 => x"C0C0C0F982F9A492",
 16126 => x"C0C0C0F982F9A482",
 16127 => x"C0C0C0F982F9A4F8",
 16128 => x"C0C0C0F982F9A480",
 16129 => x"C0C0C0F982F9A490",
 16130 => x"C0C0C0F982F9B0C0",
 16131 => x"C0C0C0F982F9B0F9",
 16132 => x"C0C0C0F982F9B0A4",
 16133 => x"C0C0C0F982F9B0B0",
 16134 => x"C0C0C0F982F9B099",
 16135 => x"C0C0C0F982F9B092",
 16136 => x"C0C0C0F982F9B082",
 16137 => x"C0C0C0F982F9B0F8",
 16138 => x"C0C0C0F982F9B080",
 16139 => x"C0C0C0F982F9B090",
 16140 => x"C0C0C0F982F999C0",
 16141 => x"C0C0C0F982F999F9",
 16142 => x"C0C0C0F982F999A4",
 16143 => x"C0C0C0F982F999B0",
 16144 => x"C0C0C0F982F99999",
 16145 => x"C0C0C0F982F99992",
 16146 => x"C0C0C0F982F99982",
 16147 => x"C0C0C0F982F999F8",
 16148 => x"C0C0C0F982F99980",
 16149 => x"C0C0C0F982F99990",
 16150 => x"C0C0C0F982F992C0",
 16151 => x"C0C0C0F982F992F9",
 16152 => x"C0C0C0F982F992A4",
 16153 => x"C0C0C0F982F992B0",
 16154 => x"C0C0C0F982F99299",
 16155 => x"C0C0C0F982F99292",
 16156 => x"C0C0C0F982F99282",
 16157 => x"C0C0C0F982F992F8",
 16158 => x"C0C0C0F982F99280",
 16159 => x"C0C0C0F982F99290",
 16160 => x"C0C0C0F982F982C0",
 16161 => x"C0C0C0F982F982F9",
 16162 => x"C0C0C0F982F982A4",
 16163 => x"C0C0C0F982F982B0",
 16164 => x"C0C0C0F982F98299",
 16165 => x"C0C0C0F982F98292",
 16166 => x"C0C0C0F982F98282",
 16167 => x"C0C0C0F982F982F8",
 16168 => x"C0C0C0F982F98280",
 16169 => x"C0C0C0F982F98290",
 16170 => x"C0C0C0F982F9F8C0",
 16171 => x"C0C0C0F982F9F8F9",
 16172 => x"C0C0C0F982F9F8A4",
 16173 => x"C0C0C0F982F9F8B0",
 16174 => x"C0C0C0F982F9F899",
 16175 => x"C0C0C0F982F9F892",
 16176 => x"C0C0C0F982F9F882",
 16177 => x"C0C0C0F982F9F8F8",
 16178 => x"C0C0C0F982F9F880",
 16179 => x"C0C0C0F982F9F890",
 16180 => x"C0C0C0F982F980C0",
 16181 => x"C0C0C0F982F980F9",
 16182 => x"C0C0C0F982F980A4",
 16183 => x"C0C0C0F982F980B0",
 16184 => x"C0C0C0F982F98099",
 16185 => x"C0C0C0F982F98092",
 16186 => x"C0C0C0F982F98082",
 16187 => x"C0C0C0F982F980F8",
 16188 => x"C0C0C0F982F98080",
 16189 => x"C0C0C0F982F98090",
 16190 => x"C0C0C0F982F990C0",
 16191 => x"C0C0C0F982F990F9",
 16192 => x"C0C0C0F982F990A4",
 16193 => x"C0C0C0F982F990B0",
 16194 => x"C0C0C0F982F99099",
 16195 => x"C0C0C0F982F99092",
 16196 => x"C0C0C0F982F99082",
 16197 => x"C0C0C0F982F990F8",
 16198 => x"C0C0C0F982F99080",
 16199 => x"C0C0C0F982F99090",
 16200 => x"C0C0C0F982A4C0C0",
 16201 => x"C0C0C0F982A4C0F9",
 16202 => x"C0C0C0F982A4C0A4",
 16203 => x"C0C0C0F982A4C0B0",
 16204 => x"C0C0C0F982A4C099",
 16205 => x"C0C0C0F982A4C092",
 16206 => x"C0C0C0F982A4C082",
 16207 => x"C0C0C0F982A4C0F8",
 16208 => x"C0C0C0F982A4C080",
 16209 => x"C0C0C0F982A4C090",
 16210 => x"C0C0C0F982A4F9C0",
 16211 => x"C0C0C0F982A4F9F9",
 16212 => x"C0C0C0F982A4F9A4",
 16213 => x"C0C0C0F982A4F9B0",
 16214 => x"C0C0C0F982A4F999",
 16215 => x"C0C0C0F982A4F992",
 16216 => x"C0C0C0F982A4F982",
 16217 => x"C0C0C0F982A4F9F8",
 16218 => x"C0C0C0F982A4F980",
 16219 => x"C0C0C0F982A4F990",
 16220 => x"C0C0C0F982A4A4C0",
 16221 => x"C0C0C0F982A4A4F9",
 16222 => x"C0C0C0F982A4A4A4",
 16223 => x"C0C0C0F982A4A4B0",
 16224 => x"C0C0C0F982A4A499",
 16225 => x"C0C0C0F982A4A492",
 16226 => x"C0C0C0F982A4A482",
 16227 => x"C0C0C0F982A4A4F8",
 16228 => x"C0C0C0F982A4A480",
 16229 => x"C0C0C0F982A4A490",
 16230 => x"C0C0C0F982A4B0C0",
 16231 => x"C0C0C0F982A4B0F9",
 16232 => x"C0C0C0F982A4B0A4",
 16233 => x"C0C0C0F982A4B0B0",
 16234 => x"C0C0C0F982A4B099",
 16235 => x"C0C0C0F982A4B092",
 16236 => x"C0C0C0F982A4B082",
 16237 => x"C0C0C0F982A4B0F8",
 16238 => x"C0C0C0F982A4B080",
 16239 => x"C0C0C0F982A4B090",
 16240 => x"C0C0C0F982A499C0",
 16241 => x"C0C0C0F982A499F9",
 16242 => x"C0C0C0F982A499A4",
 16243 => x"C0C0C0F982A499B0",
 16244 => x"C0C0C0F982A49999",
 16245 => x"C0C0C0F982A49992",
 16246 => x"C0C0C0F982A49982",
 16247 => x"C0C0C0F982A499F8",
 16248 => x"C0C0C0F982A49980",
 16249 => x"C0C0C0F982A49990",
 16250 => x"C0C0C0F982A492C0",
 16251 => x"C0C0C0F982A492F9",
 16252 => x"C0C0C0F982A492A4",
 16253 => x"C0C0C0F982A492B0",
 16254 => x"C0C0C0F982A49299",
 16255 => x"C0C0C0F982A49292",
 16256 => x"C0C0C0F982A49282",
 16257 => x"C0C0C0F982A492F8",
 16258 => x"C0C0C0F982A49280",
 16259 => x"C0C0C0F982A49290",
 16260 => x"C0C0C0F982A482C0",
 16261 => x"C0C0C0F982A482F9",
 16262 => x"C0C0C0F982A482A4",
 16263 => x"C0C0C0F982A482B0",
 16264 => x"C0C0C0F982A48299",
 16265 => x"C0C0C0F982A48292",
 16266 => x"C0C0C0F982A48282",
 16267 => x"C0C0C0F982A482F8",
 16268 => x"C0C0C0F982A48280",
 16269 => x"C0C0C0F982A48290",
 16270 => x"C0C0C0F982A4F8C0",
 16271 => x"C0C0C0F982A4F8F9",
 16272 => x"C0C0C0F982A4F8A4",
 16273 => x"C0C0C0F982A4F8B0",
 16274 => x"C0C0C0F982A4F899",
 16275 => x"C0C0C0F982A4F892",
 16276 => x"C0C0C0F982A4F882",
 16277 => x"C0C0C0F982A4F8F8",
 16278 => x"C0C0C0F982A4F880",
 16279 => x"C0C0C0F982A4F890",
 16280 => x"C0C0C0F982A480C0",
 16281 => x"C0C0C0F982A480F9",
 16282 => x"C0C0C0F982A480A4",
 16283 => x"C0C0C0F982A480B0",
 16284 => x"C0C0C0F982A48099",
 16285 => x"C0C0C0F982A48092",
 16286 => x"C0C0C0F982A48082",
 16287 => x"C0C0C0F982A480F8",
 16288 => x"C0C0C0F982A48080",
 16289 => x"C0C0C0F982A48090",
 16290 => x"C0C0C0F982A490C0",
 16291 => x"C0C0C0F982A490F9",
 16292 => x"C0C0C0F982A490A4",
 16293 => x"C0C0C0F982A490B0",
 16294 => x"C0C0C0F982A49099",
 16295 => x"C0C0C0F982A49092",
 16296 => x"C0C0C0F982A49082",
 16297 => x"C0C0C0F982A490F8",
 16298 => x"C0C0C0F982A49080",
 16299 => x"C0C0C0F982A49090",
 16300 => x"C0C0C0F982B0C0C0",
 16301 => x"C0C0C0F982B0C0F9",
 16302 => x"C0C0C0F982B0C0A4",
 16303 => x"C0C0C0F982B0C0B0",
 16304 => x"C0C0C0F982B0C099",
 16305 => x"C0C0C0F982B0C092",
 16306 => x"C0C0C0F982B0C082",
 16307 => x"C0C0C0F982B0C0F8",
 16308 => x"C0C0C0F982B0C080",
 16309 => x"C0C0C0F982B0C090",
 16310 => x"C0C0C0F982B0F9C0",
 16311 => x"C0C0C0F982B0F9F9",
 16312 => x"C0C0C0F982B0F9A4",
 16313 => x"C0C0C0F982B0F9B0",
 16314 => x"C0C0C0F982B0F999",
 16315 => x"C0C0C0F982B0F992",
 16316 => x"C0C0C0F982B0F982",
 16317 => x"C0C0C0F982B0F9F8",
 16318 => x"C0C0C0F982B0F980",
 16319 => x"C0C0C0F982B0F990",
 16320 => x"C0C0C0F982B0A4C0",
 16321 => x"C0C0C0F982B0A4F9",
 16322 => x"C0C0C0F982B0A4A4",
 16323 => x"C0C0C0F982B0A4B0",
 16324 => x"C0C0C0F982B0A499",
 16325 => x"C0C0C0F982B0A492",
 16326 => x"C0C0C0F982B0A482",
 16327 => x"C0C0C0F982B0A4F8",
 16328 => x"C0C0C0F982B0A480",
 16329 => x"C0C0C0F982B0A490",
 16330 => x"C0C0C0F982B0B0C0",
 16331 => x"C0C0C0F982B0B0F9",
 16332 => x"C0C0C0F982B0B0A4",
 16333 => x"C0C0C0F982B0B0B0",
 16334 => x"C0C0C0F982B0B099",
 16335 => x"C0C0C0F982B0B092",
 16336 => x"C0C0C0F982B0B082",
 16337 => x"C0C0C0F982B0B0F8",
 16338 => x"C0C0C0F982B0B080",
 16339 => x"C0C0C0F982B0B090",
 16340 => x"C0C0C0F982B099C0",
 16341 => x"C0C0C0F982B099F9",
 16342 => x"C0C0C0F982B099A4",
 16343 => x"C0C0C0F982B099B0",
 16344 => x"C0C0C0F982B09999",
 16345 => x"C0C0C0F982B09992",
 16346 => x"C0C0C0F982B09982",
 16347 => x"C0C0C0F982B099F8",
 16348 => x"C0C0C0F982B09980",
 16349 => x"C0C0C0F982B09990",
 16350 => x"C0C0C0F982B092C0",
 16351 => x"C0C0C0F982B092F9",
 16352 => x"C0C0C0F982B092A4",
 16353 => x"C0C0C0F982B092B0",
 16354 => x"C0C0C0F982B09299",
 16355 => x"C0C0C0F982B09292",
 16356 => x"C0C0C0F982B09282",
 16357 => x"C0C0C0F982B092F8",
 16358 => x"C0C0C0F982B09280",
 16359 => x"C0C0C0F982B09290",
 16360 => x"C0C0C0F982B082C0",
 16361 => x"C0C0C0F982B082F9",
 16362 => x"C0C0C0F982B082A4",
 16363 => x"C0C0C0F982B082B0",
 16364 => x"C0C0C0F982B08299",
 16365 => x"C0C0C0F982B08292",
 16366 => x"C0C0C0F982B08282",
 16367 => x"C0C0C0F982B082F8",
 16368 => x"C0C0C0F982B08280",
 16369 => x"C0C0C0F982B08290",
 16370 => x"C0C0C0F982B0F8C0",
 16371 => x"C0C0C0F982B0F8F9",
 16372 => x"C0C0C0F982B0F8A4",
 16373 => x"C0C0C0F982B0F8B0",
 16374 => x"C0C0C0F982B0F899",
 16375 => x"C0C0C0F982B0F892",
 16376 => x"C0C0C0F982B0F882",
 16377 => x"C0C0C0F982B0F8F8",
 16378 => x"C0C0C0F982B0F880",
 16379 => x"C0C0C0F982B0F890",
 16380 => x"C0C0C0F982B080C0",
 16381 => x"C0C0C0F982B080F9",
 16382 => x"C0C0C0F982B080A4",
 16383 => x"C0C0C0F982B080B0",
 16384 => x"C0C0C0F982B08099",
 16385 => x"C0C0C0F982B08092",
 16386 => x"C0C0C0F982B08082",
 16387 => x"C0C0C0F982B080F8",
 16388 => x"C0C0C0F982B08080",
 16389 => x"C0C0C0F982B08090",
 16390 => x"C0C0C0F982B090C0",
 16391 => x"C0C0C0F982B090F9",
 16392 => x"C0C0C0F982B090A4",
 16393 => x"C0C0C0F982B090B0",
 16394 => x"C0C0C0F982B09099",
 16395 => x"C0C0C0F982B09092",
 16396 => x"C0C0C0F982B09082",
 16397 => x"C0C0C0F982B090F8",
 16398 => x"C0C0C0F982B09080",
 16399 => x"C0C0C0F982B09090",
 16400 => x"C0C0C0F98299C0C0",
 16401 => x"C0C0C0F98299C0F9",
 16402 => x"C0C0C0F98299C0A4",
 16403 => x"C0C0C0F98299C0B0",
 16404 => x"C0C0C0F98299C099",
 16405 => x"C0C0C0F98299C092",
 16406 => x"C0C0C0F98299C082",
 16407 => x"C0C0C0F98299C0F8",
 16408 => x"C0C0C0F98299C080",
 16409 => x"C0C0C0F98299C090",
 16410 => x"C0C0C0F98299F9C0",
 16411 => x"C0C0C0F98299F9F9",
 16412 => x"C0C0C0F98299F9A4",
 16413 => x"C0C0C0F98299F9B0",
 16414 => x"C0C0C0F98299F999",
 16415 => x"C0C0C0F98299F992",
 16416 => x"C0C0C0F98299F982",
 16417 => x"C0C0C0F98299F9F8",
 16418 => x"C0C0C0F98299F980",
 16419 => x"C0C0C0F98299F990",
 16420 => x"C0C0C0F98299A4C0",
 16421 => x"C0C0C0F98299A4F9",
 16422 => x"C0C0C0F98299A4A4",
 16423 => x"C0C0C0F98299A4B0",
 16424 => x"C0C0C0F98299A499",
 16425 => x"C0C0C0F98299A492",
 16426 => x"C0C0C0F98299A482",
 16427 => x"C0C0C0F98299A4F8",
 16428 => x"C0C0C0F98299A480",
 16429 => x"C0C0C0F98299A490",
 16430 => x"C0C0C0F98299B0C0",
 16431 => x"C0C0C0F98299B0F9",
 16432 => x"C0C0C0F98299B0A4",
 16433 => x"C0C0C0F98299B0B0",
 16434 => x"C0C0C0F98299B099",
 16435 => x"C0C0C0F98299B092",
 16436 => x"C0C0C0F98299B082",
 16437 => x"C0C0C0F98299B0F8",
 16438 => x"C0C0C0F98299B080",
 16439 => x"C0C0C0F98299B090",
 16440 => x"C0C0C0F9829999C0",
 16441 => x"C0C0C0F9829999F9",
 16442 => x"C0C0C0F9829999A4",
 16443 => x"C0C0C0F9829999B0",
 16444 => x"C0C0C0F982999999",
 16445 => x"C0C0C0F982999992",
 16446 => x"C0C0C0F982999982",
 16447 => x"C0C0C0F9829999F8",
 16448 => x"C0C0C0F982999980",
 16449 => x"C0C0C0F982999990",
 16450 => x"C0C0C0F9829992C0",
 16451 => x"C0C0C0F9829992F9",
 16452 => x"C0C0C0F9829992A4",
 16453 => x"C0C0C0F9829992B0",
 16454 => x"C0C0C0F982999299",
 16455 => x"C0C0C0F982999292",
 16456 => x"C0C0C0F982999282",
 16457 => x"C0C0C0F9829992F8",
 16458 => x"C0C0C0F982999280",
 16459 => x"C0C0C0F982999290",
 16460 => x"C0C0C0F9829982C0",
 16461 => x"C0C0C0F9829982F9",
 16462 => x"C0C0C0F9829982A4",
 16463 => x"C0C0C0F9829982B0",
 16464 => x"C0C0C0F982998299",
 16465 => x"C0C0C0F982998292",
 16466 => x"C0C0C0F982998282",
 16467 => x"C0C0C0F9829982F8",
 16468 => x"C0C0C0F982998280",
 16469 => x"C0C0C0F982998290",
 16470 => x"C0C0C0F98299F8C0",
 16471 => x"C0C0C0F98299F8F9",
 16472 => x"C0C0C0F98299F8A4",
 16473 => x"C0C0C0F98299F8B0",
 16474 => x"C0C0C0F98299F899",
 16475 => x"C0C0C0F98299F892",
 16476 => x"C0C0C0F98299F882",
 16477 => x"C0C0C0F98299F8F8",
 16478 => x"C0C0C0F98299F880",
 16479 => x"C0C0C0F98299F890",
 16480 => x"C0C0C0F9829980C0",
 16481 => x"C0C0C0F9829980F9",
 16482 => x"C0C0C0F9829980A4",
 16483 => x"C0C0C0F9829980B0",
 16484 => x"C0C0C0F982998099",
 16485 => x"C0C0C0F982998092",
 16486 => x"C0C0C0F982998082",
 16487 => x"C0C0C0F9829980F8",
 16488 => x"C0C0C0F982998080",
 16489 => x"C0C0C0F982998090",
 16490 => x"C0C0C0F9829990C0",
 16491 => x"C0C0C0F9829990F9",
 16492 => x"C0C0C0F9829990A4",
 16493 => x"C0C0C0F9829990B0",
 16494 => x"C0C0C0F982999099",
 16495 => x"C0C0C0F982999092",
 16496 => x"C0C0C0F982999082",
 16497 => x"C0C0C0F9829990F8",
 16498 => x"C0C0C0F982999080",
 16499 => x"C0C0C0F982999090",
 16500 => x"C0C0C0F98292C0C0",
 16501 => x"C0C0C0F98292C0F9",
 16502 => x"C0C0C0F98292C0A4",
 16503 => x"C0C0C0F98292C0B0",
 16504 => x"C0C0C0F98292C099",
 16505 => x"C0C0C0F98292C092",
 16506 => x"C0C0C0F98292C082",
 16507 => x"C0C0C0F98292C0F8",
 16508 => x"C0C0C0F98292C080",
 16509 => x"C0C0C0F98292C090",
 16510 => x"C0C0C0F98292F9C0",
 16511 => x"C0C0C0F98292F9F9",
 16512 => x"C0C0C0F98292F9A4",
 16513 => x"C0C0C0F98292F9B0",
 16514 => x"C0C0C0F98292F999",
 16515 => x"C0C0C0F98292F992",
 16516 => x"C0C0C0F98292F982",
 16517 => x"C0C0C0F98292F9F8",
 16518 => x"C0C0C0F98292F980",
 16519 => x"C0C0C0F98292F990",
 16520 => x"C0C0C0F98292A4C0",
 16521 => x"C0C0C0F98292A4F9",
 16522 => x"C0C0C0F98292A4A4",
 16523 => x"C0C0C0F98292A4B0",
 16524 => x"C0C0C0F98292A499",
 16525 => x"C0C0C0F98292A492",
 16526 => x"C0C0C0F98292A482",
 16527 => x"C0C0C0F98292A4F8",
 16528 => x"C0C0C0F98292A480",
 16529 => x"C0C0C0F98292A490",
 16530 => x"C0C0C0F98292B0C0",
 16531 => x"C0C0C0F98292B0F9",
 16532 => x"C0C0C0F98292B0A4",
 16533 => x"C0C0C0F98292B0B0",
 16534 => x"C0C0C0F98292B099",
 16535 => x"C0C0C0F98292B092",
 16536 => x"C0C0C0F98292B082",
 16537 => x"C0C0C0F98292B0F8",
 16538 => x"C0C0C0F98292B080",
 16539 => x"C0C0C0F98292B090",
 16540 => x"C0C0C0F9829299C0",
 16541 => x"C0C0C0F9829299F9",
 16542 => x"C0C0C0F9829299A4",
 16543 => x"C0C0C0F9829299B0",
 16544 => x"C0C0C0F982929999",
 16545 => x"C0C0C0F982929992",
 16546 => x"C0C0C0F982929982",
 16547 => x"C0C0C0F9829299F8",
 16548 => x"C0C0C0F982929980",
 16549 => x"C0C0C0F982929990",
 16550 => x"C0C0C0F9829292C0",
 16551 => x"C0C0C0F9829292F9",
 16552 => x"C0C0C0F9829292A4",
 16553 => x"C0C0C0F9829292B0",
 16554 => x"C0C0C0F982929299",
 16555 => x"C0C0C0F982929292",
 16556 => x"C0C0C0F982929282",
 16557 => x"C0C0C0F9829292F8",
 16558 => x"C0C0C0F982929280",
 16559 => x"C0C0C0F982929290",
 16560 => x"C0C0C0F9829282C0",
 16561 => x"C0C0C0F9829282F9",
 16562 => x"C0C0C0F9829282A4",
 16563 => x"C0C0C0F9829282B0",
 16564 => x"C0C0C0F982928299",
 16565 => x"C0C0C0F982928292",
 16566 => x"C0C0C0F982928282",
 16567 => x"C0C0C0F9829282F8",
 16568 => x"C0C0C0F982928280",
 16569 => x"C0C0C0F982928290",
 16570 => x"C0C0C0F98292F8C0",
 16571 => x"C0C0C0F98292F8F9",
 16572 => x"C0C0C0F98292F8A4",
 16573 => x"C0C0C0F98292F8B0",
 16574 => x"C0C0C0F98292F899",
 16575 => x"C0C0C0F98292F892",
 16576 => x"C0C0C0F98292F882",
 16577 => x"C0C0C0F98292F8F8",
 16578 => x"C0C0C0F98292F880",
 16579 => x"C0C0C0F98292F890",
 16580 => x"C0C0C0F9829280C0",
 16581 => x"C0C0C0F9829280F9",
 16582 => x"C0C0C0F9829280A4",
 16583 => x"C0C0C0F9829280B0",
 16584 => x"C0C0C0F982928099",
 16585 => x"C0C0C0F982928092",
 16586 => x"C0C0C0F982928082",
 16587 => x"C0C0C0F9829280F8",
 16588 => x"C0C0C0F982928080",
 16589 => x"C0C0C0F982928090",
 16590 => x"C0C0C0F9829290C0",
 16591 => x"C0C0C0F9829290F9",
 16592 => x"C0C0C0F9829290A4",
 16593 => x"C0C0C0F9829290B0",
 16594 => x"C0C0C0F982929099",
 16595 => x"C0C0C0F982929092",
 16596 => x"C0C0C0F982929082",
 16597 => x"C0C0C0F9829290F8",
 16598 => x"C0C0C0F982929080",
 16599 => x"C0C0C0F982929090",
 16600 => x"C0C0C0F98282C0C0",
 16601 => x"C0C0C0F98282C0F9",
 16602 => x"C0C0C0F98282C0A4",
 16603 => x"C0C0C0F98282C0B0",
 16604 => x"C0C0C0F98282C099",
 16605 => x"C0C0C0F98282C092",
 16606 => x"C0C0C0F98282C082",
 16607 => x"C0C0C0F98282C0F8",
 16608 => x"C0C0C0F98282C080",
 16609 => x"C0C0C0F98282C090",
 16610 => x"C0C0C0F98282F9C0",
 16611 => x"C0C0C0F98282F9F9",
 16612 => x"C0C0C0F98282F9A4",
 16613 => x"C0C0C0F98282F9B0",
 16614 => x"C0C0C0F98282F999",
 16615 => x"C0C0C0F98282F992",
 16616 => x"C0C0C0F98282F982",
 16617 => x"C0C0C0F98282F9F8",
 16618 => x"C0C0C0F98282F980",
 16619 => x"C0C0C0F98282F990",
 16620 => x"C0C0C0F98282A4C0",
 16621 => x"C0C0C0F98282A4F9",
 16622 => x"C0C0C0F98282A4A4",
 16623 => x"C0C0C0F98282A4B0",
 16624 => x"C0C0C0F98282A499",
 16625 => x"C0C0C0F98282A492",
 16626 => x"C0C0C0F98282A482",
 16627 => x"C0C0C0F98282A4F8",
 16628 => x"C0C0C0F98282A480",
 16629 => x"C0C0C0F98282A490",
 16630 => x"C0C0C0F98282B0C0",
 16631 => x"C0C0C0F98282B0F9",
 16632 => x"C0C0C0F98282B0A4",
 16633 => x"C0C0C0F98282B0B0",
 16634 => x"C0C0C0F98282B099",
 16635 => x"C0C0C0F98282B092",
 16636 => x"C0C0C0F98282B082",
 16637 => x"C0C0C0F98282B0F8",
 16638 => x"C0C0C0F98282B080",
 16639 => x"C0C0C0F98282B090",
 16640 => x"C0C0C0F9828299C0",
 16641 => x"C0C0C0F9828299F9",
 16642 => x"C0C0C0F9828299A4",
 16643 => x"C0C0C0F9828299B0",
 16644 => x"C0C0C0F982829999",
 16645 => x"C0C0C0F982829992",
 16646 => x"C0C0C0F982829982",
 16647 => x"C0C0C0F9828299F8",
 16648 => x"C0C0C0F982829980",
 16649 => x"C0C0C0F982829990",
 16650 => x"C0C0C0F9828292C0",
 16651 => x"C0C0C0F9828292F9",
 16652 => x"C0C0C0F9828292A4",
 16653 => x"C0C0C0F9828292B0",
 16654 => x"C0C0C0F982829299",
 16655 => x"C0C0C0F982829292",
 16656 => x"C0C0C0F982829282",
 16657 => x"C0C0C0F9828292F8",
 16658 => x"C0C0C0F982829280",
 16659 => x"C0C0C0F982829290",
 16660 => x"C0C0C0F9828282C0",
 16661 => x"C0C0C0F9828282F9",
 16662 => x"C0C0C0F9828282A4",
 16663 => x"C0C0C0F9828282B0",
 16664 => x"C0C0C0F982828299",
 16665 => x"C0C0C0F982828292",
 16666 => x"C0C0C0F982828282",
 16667 => x"C0C0C0F9828282F8",
 16668 => x"C0C0C0F982828280",
 16669 => x"C0C0C0F982828290",
 16670 => x"C0C0C0F98282F8C0",
 16671 => x"C0C0C0F98282F8F9",
 16672 => x"C0C0C0F98282F8A4",
 16673 => x"C0C0C0F98282F8B0",
 16674 => x"C0C0C0F98282F899",
 16675 => x"C0C0C0F98282F892",
 16676 => x"C0C0C0F98282F882",
 16677 => x"C0C0C0F98282F8F8",
 16678 => x"C0C0C0F98282F880",
 16679 => x"C0C0C0F98282F890",
 16680 => x"C0C0C0F9828280C0",
 16681 => x"C0C0C0F9828280F9",
 16682 => x"C0C0C0F9828280A4",
 16683 => x"C0C0C0F9828280B0",
 16684 => x"C0C0C0F982828099",
 16685 => x"C0C0C0F982828092",
 16686 => x"C0C0C0F982828082",
 16687 => x"C0C0C0F9828280F8",
 16688 => x"C0C0C0F982828080",
 16689 => x"C0C0C0F982828090",
 16690 => x"C0C0C0F9828290C0",
 16691 => x"C0C0C0F9828290F9",
 16692 => x"C0C0C0F9828290A4",
 16693 => x"C0C0C0F9828290B0",
 16694 => x"C0C0C0F982829099",
 16695 => x"C0C0C0F982829092",
 16696 => x"C0C0C0F982829082",
 16697 => x"C0C0C0F9828290F8",
 16698 => x"C0C0C0F982829080",
 16699 => x"C0C0C0F982829090",
 16700 => x"C0C0C0F982F8C0C0",
 16701 => x"C0C0C0F982F8C0F9",
 16702 => x"C0C0C0F982F8C0A4",
 16703 => x"C0C0C0F982F8C0B0",
 16704 => x"C0C0C0F982F8C099",
 16705 => x"C0C0C0F982F8C092",
 16706 => x"C0C0C0F982F8C082",
 16707 => x"C0C0C0F982F8C0F8",
 16708 => x"C0C0C0F982F8C080",
 16709 => x"C0C0C0F982F8C090",
 16710 => x"C0C0C0F982F8F9C0",
 16711 => x"C0C0C0F982F8F9F9",
 16712 => x"C0C0C0F982F8F9A4",
 16713 => x"C0C0C0F982F8F9B0",
 16714 => x"C0C0C0F982F8F999",
 16715 => x"C0C0C0F982F8F992",
 16716 => x"C0C0C0F982F8F982",
 16717 => x"C0C0C0F982F8F9F8",
 16718 => x"C0C0C0F982F8F980",
 16719 => x"C0C0C0F982F8F990",
 16720 => x"C0C0C0F982F8A4C0",
 16721 => x"C0C0C0F982F8A4F9",
 16722 => x"C0C0C0F982F8A4A4",
 16723 => x"C0C0C0F982F8A4B0",
 16724 => x"C0C0C0F982F8A499",
 16725 => x"C0C0C0F982F8A492",
 16726 => x"C0C0C0F982F8A482",
 16727 => x"C0C0C0F982F8A4F8",
 16728 => x"C0C0C0F982F8A480",
 16729 => x"C0C0C0F982F8A490",
 16730 => x"C0C0C0F982F8B0C0",
 16731 => x"C0C0C0F982F8B0F9",
 16732 => x"C0C0C0F982F8B0A4",
 16733 => x"C0C0C0F982F8B0B0",
 16734 => x"C0C0C0F982F8B099",
 16735 => x"C0C0C0F982F8B092",
 16736 => x"C0C0C0F982F8B082",
 16737 => x"C0C0C0F982F8B0F8",
 16738 => x"C0C0C0F982F8B080",
 16739 => x"C0C0C0F982F8B090",
 16740 => x"C0C0C0F982F899C0",
 16741 => x"C0C0C0F982F899F9",
 16742 => x"C0C0C0F982F899A4",
 16743 => x"C0C0C0F982F899B0",
 16744 => x"C0C0C0F982F89999",
 16745 => x"C0C0C0F982F89992",
 16746 => x"C0C0C0F982F89982",
 16747 => x"C0C0C0F982F899F8",
 16748 => x"C0C0C0F982F89980",
 16749 => x"C0C0C0F982F89990",
 16750 => x"C0C0C0F982F892C0",
 16751 => x"C0C0C0F982F892F9",
 16752 => x"C0C0C0F982F892A4",
 16753 => x"C0C0C0F982F892B0",
 16754 => x"C0C0C0F982F89299",
 16755 => x"C0C0C0F982F89292",
 16756 => x"C0C0C0F982F89282",
 16757 => x"C0C0C0F982F892F8",
 16758 => x"C0C0C0F982F89280",
 16759 => x"C0C0C0F982F89290",
 16760 => x"C0C0C0F982F882C0",
 16761 => x"C0C0C0F982F882F9",
 16762 => x"C0C0C0F982F882A4",
 16763 => x"C0C0C0F982F882B0",
 16764 => x"C0C0C0F982F88299",
 16765 => x"C0C0C0F982F88292",
 16766 => x"C0C0C0F982F88282",
 16767 => x"C0C0C0F982F882F8",
 16768 => x"C0C0C0F982F88280",
 16769 => x"C0C0C0F982F88290",
 16770 => x"C0C0C0F982F8F8C0",
 16771 => x"C0C0C0F982F8F8F9",
 16772 => x"C0C0C0F982F8F8A4",
 16773 => x"C0C0C0F982F8F8B0",
 16774 => x"C0C0C0F982F8F899",
 16775 => x"C0C0C0F982F8F892",
 16776 => x"C0C0C0F982F8F882",
 16777 => x"C0C0C0F982F8F8F8",
 16778 => x"C0C0C0F982F8F880",
 16779 => x"C0C0C0F982F8F890",
 16780 => x"C0C0C0F982F880C0",
 16781 => x"C0C0C0F982F880F9",
 16782 => x"C0C0C0F982F880A4",
 16783 => x"C0C0C0F982F880B0",
 16784 => x"C0C0C0F982F88099",
 16785 => x"C0C0C0F982F88092",
 16786 => x"C0C0C0F982F88082",
 16787 => x"C0C0C0F982F880F8",
 16788 => x"C0C0C0F982F88080",
 16789 => x"C0C0C0F982F88090",
 16790 => x"C0C0C0F982F890C0",
 16791 => x"C0C0C0F982F890F9",
 16792 => x"C0C0C0F982F890A4",
 16793 => x"C0C0C0F982F890B0",
 16794 => x"C0C0C0F982F89099",
 16795 => x"C0C0C0F982F89092",
 16796 => x"C0C0C0F982F89082",
 16797 => x"C0C0C0F982F890F8",
 16798 => x"C0C0C0F982F89080",
 16799 => x"C0C0C0F982F89090",
 16800 => x"C0C0C0F98280C0C0",
 16801 => x"C0C0C0F98280C0F9",
 16802 => x"C0C0C0F98280C0A4",
 16803 => x"C0C0C0F98280C0B0",
 16804 => x"C0C0C0F98280C099",
 16805 => x"C0C0C0F98280C092",
 16806 => x"C0C0C0F98280C082",
 16807 => x"C0C0C0F98280C0F8",
 16808 => x"C0C0C0F98280C080",
 16809 => x"C0C0C0F98280C090",
 16810 => x"C0C0C0F98280F9C0",
 16811 => x"C0C0C0F98280F9F9",
 16812 => x"C0C0C0F98280F9A4",
 16813 => x"C0C0C0F98280F9B0",
 16814 => x"C0C0C0F98280F999",
 16815 => x"C0C0C0F98280F992",
 16816 => x"C0C0C0F98280F982",
 16817 => x"C0C0C0F98280F9F8",
 16818 => x"C0C0C0F98280F980",
 16819 => x"C0C0C0F98280F990",
 16820 => x"C0C0C0F98280A4C0",
 16821 => x"C0C0C0F98280A4F9",
 16822 => x"C0C0C0F98280A4A4",
 16823 => x"C0C0C0F98280A4B0",
 16824 => x"C0C0C0F98280A499",
 16825 => x"C0C0C0F98280A492",
 16826 => x"C0C0C0F98280A482",
 16827 => x"C0C0C0F98280A4F8",
 16828 => x"C0C0C0F98280A480",
 16829 => x"C0C0C0F98280A490",
 16830 => x"C0C0C0F98280B0C0",
 16831 => x"C0C0C0F98280B0F9",
 16832 => x"C0C0C0F98280B0A4",
 16833 => x"C0C0C0F98280B0B0",
 16834 => x"C0C0C0F98280B099",
 16835 => x"C0C0C0F98280B092",
 16836 => x"C0C0C0F98280B082",
 16837 => x"C0C0C0F98280B0F8",
 16838 => x"C0C0C0F98280B080",
 16839 => x"C0C0C0F98280B090",
 16840 => x"C0C0C0F9828099C0",
 16841 => x"C0C0C0F9828099F9",
 16842 => x"C0C0C0F9828099A4",
 16843 => x"C0C0C0F9828099B0",
 16844 => x"C0C0C0F982809999",
 16845 => x"C0C0C0F982809992",
 16846 => x"C0C0C0F982809982",
 16847 => x"C0C0C0F9828099F8",
 16848 => x"C0C0C0F982809980",
 16849 => x"C0C0C0F982809990",
 16850 => x"C0C0C0F9828092C0",
 16851 => x"C0C0C0F9828092F9",
 16852 => x"C0C0C0F9828092A4",
 16853 => x"C0C0C0F9828092B0",
 16854 => x"C0C0C0F982809299",
 16855 => x"C0C0C0F982809292",
 16856 => x"C0C0C0F982809282",
 16857 => x"C0C0C0F9828092F8",
 16858 => x"C0C0C0F982809280",
 16859 => x"C0C0C0F982809290",
 16860 => x"C0C0C0F9828082C0",
 16861 => x"C0C0C0F9828082F9",
 16862 => x"C0C0C0F9828082A4",
 16863 => x"C0C0C0F9828082B0",
 16864 => x"C0C0C0F982808299",
 16865 => x"C0C0C0F982808292",
 16866 => x"C0C0C0F982808282",
 16867 => x"C0C0C0F9828082F8",
 16868 => x"C0C0C0F982808280",
 16869 => x"C0C0C0F982808290",
 16870 => x"C0C0C0F98280F8C0",
 16871 => x"C0C0C0F98280F8F9",
 16872 => x"C0C0C0F98280F8A4",
 16873 => x"C0C0C0F98280F8B0",
 16874 => x"C0C0C0F98280F899",
 16875 => x"C0C0C0F98280F892",
 16876 => x"C0C0C0F98280F882",
 16877 => x"C0C0C0F98280F8F8",
 16878 => x"C0C0C0F98280F880",
 16879 => x"C0C0C0F98280F890",
 16880 => x"C0C0C0F9828080C0",
 16881 => x"C0C0C0F9828080F9",
 16882 => x"C0C0C0F9828080A4",
 16883 => x"C0C0C0F9828080B0",
 16884 => x"C0C0C0F982808099",
 16885 => x"C0C0C0F982808092",
 16886 => x"C0C0C0F982808082",
 16887 => x"C0C0C0F9828080F8",
 16888 => x"C0C0C0F982808080",
 16889 => x"C0C0C0F982808090",
 16890 => x"C0C0C0F9828090C0",
 16891 => x"C0C0C0F9828090F9",
 16892 => x"C0C0C0F9828090A4",
 16893 => x"C0C0C0F9828090B0",
 16894 => x"C0C0C0F982809099",
 16895 => x"C0C0C0F982809092",
 16896 => x"C0C0C0F982809082",
 16897 => x"C0C0C0F9828090F8",
 16898 => x"C0C0C0F982809080",
 16899 => x"C0C0C0F982809090",
 16900 => x"C0C0C0F98290C0C0",
 16901 => x"C0C0C0F98290C0F9",
 16902 => x"C0C0C0F98290C0A4",
 16903 => x"C0C0C0F98290C0B0",
 16904 => x"C0C0C0F98290C099",
 16905 => x"C0C0C0F98290C092",
 16906 => x"C0C0C0F98290C082",
 16907 => x"C0C0C0F98290C0F8",
 16908 => x"C0C0C0F98290C080",
 16909 => x"C0C0C0F98290C090",
 16910 => x"C0C0C0F98290F9C0",
 16911 => x"C0C0C0F98290F9F9",
 16912 => x"C0C0C0F98290F9A4",
 16913 => x"C0C0C0F98290F9B0",
 16914 => x"C0C0C0F98290F999",
 16915 => x"C0C0C0F98290F992",
 16916 => x"C0C0C0F98290F982",
 16917 => x"C0C0C0F98290F9F8",
 16918 => x"C0C0C0F98290F980",
 16919 => x"C0C0C0F98290F990",
 16920 => x"C0C0C0F98290A4C0",
 16921 => x"C0C0C0F98290A4F9",
 16922 => x"C0C0C0F98290A4A4",
 16923 => x"C0C0C0F98290A4B0",
 16924 => x"C0C0C0F98290A499",
 16925 => x"C0C0C0F98290A492",
 16926 => x"C0C0C0F98290A482",
 16927 => x"C0C0C0F98290A4F8",
 16928 => x"C0C0C0F98290A480",
 16929 => x"C0C0C0F98290A490",
 16930 => x"C0C0C0F98290B0C0",
 16931 => x"C0C0C0F98290B0F9",
 16932 => x"C0C0C0F98290B0A4",
 16933 => x"C0C0C0F98290B0B0",
 16934 => x"C0C0C0F98290B099",
 16935 => x"C0C0C0F98290B092",
 16936 => x"C0C0C0F98290B082",
 16937 => x"C0C0C0F98290B0F8",
 16938 => x"C0C0C0F98290B080",
 16939 => x"C0C0C0F98290B090",
 16940 => x"C0C0C0F9829099C0",
 16941 => x"C0C0C0F9829099F9",
 16942 => x"C0C0C0F9829099A4",
 16943 => x"C0C0C0F9829099B0",
 16944 => x"C0C0C0F982909999",
 16945 => x"C0C0C0F982909992",
 16946 => x"C0C0C0F982909982",
 16947 => x"C0C0C0F9829099F8",
 16948 => x"C0C0C0F982909980",
 16949 => x"C0C0C0F982909990",
 16950 => x"C0C0C0F9829092C0",
 16951 => x"C0C0C0F9829092F9",
 16952 => x"C0C0C0F9829092A4",
 16953 => x"C0C0C0F9829092B0",
 16954 => x"C0C0C0F982909299",
 16955 => x"C0C0C0F982909292",
 16956 => x"C0C0C0F982909282",
 16957 => x"C0C0C0F9829092F8",
 16958 => x"C0C0C0F982909280",
 16959 => x"C0C0C0F982909290",
 16960 => x"C0C0C0F9829082C0",
 16961 => x"C0C0C0F9829082F9",
 16962 => x"C0C0C0F9829082A4",
 16963 => x"C0C0C0F9829082B0",
 16964 => x"C0C0C0F982908299",
 16965 => x"C0C0C0F982908292",
 16966 => x"C0C0C0F982908282",
 16967 => x"C0C0C0F9829082F8",
 16968 => x"C0C0C0F982908280",
 16969 => x"C0C0C0F982908290",
 16970 => x"C0C0C0F98290F8C0",
 16971 => x"C0C0C0F98290F8F9",
 16972 => x"C0C0C0F98290F8A4",
 16973 => x"C0C0C0F98290F8B0",
 16974 => x"C0C0C0F98290F899",
 16975 => x"C0C0C0F98290F892",
 16976 => x"C0C0C0F98290F882",
 16977 => x"C0C0C0F98290F8F8",
 16978 => x"C0C0C0F98290F880",
 16979 => x"C0C0C0F98290F890",
 16980 => x"C0C0C0F9829080C0",
 16981 => x"C0C0C0F9829080F9",
 16982 => x"C0C0C0F9829080A4",
 16983 => x"C0C0C0F9829080B0",
 16984 => x"C0C0C0F982908099",
 16985 => x"C0C0C0F982908092",
 16986 => x"C0C0C0F982908082",
 16987 => x"C0C0C0F9829080F8",
 16988 => x"C0C0C0F982908080",
 16989 => x"C0C0C0F982908090",
 16990 => x"C0C0C0F9829090C0",
 16991 => x"C0C0C0F9829090F9",
 16992 => x"C0C0C0F9829090A4",
 16993 => x"C0C0C0F9829090B0",
 16994 => x"C0C0C0F982909099",
 16995 => x"C0C0C0F982909092",
 16996 => x"C0C0C0F982909082",
 16997 => x"C0C0C0F9829090F8",
 16998 => x"C0C0C0F982909080",
 16999 => x"C0C0C0F982909090",
 17000 => x"C0C0C0F9F8C0C0C0",
 17001 => x"C0C0C0F9F8C0C0F9",
 17002 => x"C0C0C0F9F8C0C0A4",
 17003 => x"C0C0C0F9F8C0C0B0",
 17004 => x"C0C0C0F9F8C0C099",
 17005 => x"C0C0C0F9F8C0C092",
 17006 => x"C0C0C0F9F8C0C082",
 17007 => x"C0C0C0F9F8C0C0F8",
 17008 => x"C0C0C0F9F8C0C080",
 17009 => x"C0C0C0F9F8C0C090",
 17010 => x"C0C0C0F9F8C0F9C0",
 17011 => x"C0C0C0F9F8C0F9F9",
 17012 => x"C0C0C0F9F8C0F9A4",
 17013 => x"C0C0C0F9F8C0F9B0",
 17014 => x"C0C0C0F9F8C0F999",
 17015 => x"C0C0C0F9F8C0F992",
 17016 => x"C0C0C0F9F8C0F982",
 17017 => x"C0C0C0F9F8C0F9F8",
 17018 => x"C0C0C0F9F8C0F980",
 17019 => x"C0C0C0F9F8C0F990",
 17020 => x"C0C0C0F9F8C0A4C0",
 17021 => x"C0C0C0F9F8C0A4F9",
 17022 => x"C0C0C0F9F8C0A4A4",
 17023 => x"C0C0C0F9F8C0A4B0",
 17024 => x"C0C0C0F9F8C0A499",
 17025 => x"C0C0C0F9F8C0A492",
 17026 => x"C0C0C0F9F8C0A482",
 17027 => x"C0C0C0F9F8C0A4F8",
 17028 => x"C0C0C0F9F8C0A480",
 17029 => x"C0C0C0F9F8C0A490",
 17030 => x"C0C0C0F9F8C0B0C0",
 17031 => x"C0C0C0F9F8C0B0F9",
 17032 => x"C0C0C0F9F8C0B0A4",
 17033 => x"C0C0C0F9F8C0B0B0",
 17034 => x"C0C0C0F9F8C0B099",
 17035 => x"C0C0C0F9F8C0B092",
 17036 => x"C0C0C0F9F8C0B082",
 17037 => x"C0C0C0F9F8C0B0F8",
 17038 => x"C0C0C0F9F8C0B080",
 17039 => x"C0C0C0F9F8C0B090",
 17040 => x"C0C0C0F9F8C099C0",
 17041 => x"C0C0C0F9F8C099F9",
 17042 => x"C0C0C0F9F8C099A4",
 17043 => x"C0C0C0F9F8C099B0",
 17044 => x"C0C0C0F9F8C09999",
 17045 => x"C0C0C0F9F8C09992",
 17046 => x"C0C0C0F9F8C09982",
 17047 => x"C0C0C0F9F8C099F8",
 17048 => x"C0C0C0F9F8C09980",
 17049 => x"C0C0C0F9F8C09990",
 17050 => x"C0C0C0F9F8C092C0",
 17051 => x"C0C0C0F9F8C092F9",
 17052 => x"C0C0C0F9F8C092A4",
 17053 => x"C0C0C0F9F8C092B0",
 17054 => x"C0C0C0F9F8C09299",
 17055 => x"C0C0C0F9F8C09292",
 17056 => x"C0C0C0F9F8C09282",
 17057 => x"C0C0C0F9F8C092F8",
 17058 => x"C0C0C0F9F8C09280",
 17059 => x"C0C0C0F9F8C09290",
 17060 => x"C0C0C0F9F8C082C0",
 17061 => x"C0C0C0F9F8C082F9",
 17062 => x"C0C0C0F9F8C082A4",
 17063 => x"C0C0C0F9F8C082B0",
 17064 => x"C0C0C0F9F8C08299",
 17065 => x"C0C0C0F9F8C08292",
 17066 => x"C0C0C0F9F8C08282",
 17067 => x"C0C0C0F9F8C082F8",
 17068 => x"C0C0C0F9F8C08280",
 17069 => x"C0C0C0F9F8C08290",
 17070 => x"C0C0C0F9F8C0F8C0",
 17071 => x"C0C0C0F9F8C0F8F9",
 17072 => x"C0C0C0F9F8C0F8A4",
 17073 => x"C0C0C0F9F8C0F8B0",
 17074 => x"C0C0C0F9F8C0F899",
 17075 => x"C0C0C0F9F8C0F892",
 17076 => x"C0C0C0F9F8C0F882",
 17077 => x"C0C0C0F9F8C0F8F8",
 17078 => x"C0C0C0F9F8C0F880",
 17079 => x"C0C0C0F9F8C0F890",
 17080 => x"C0C0C0F9F8C080C0",
 17081 => x"C0C0C0F9F8C080F9",
 17082 => x"C0C0C0F9F8C080A4",
 17083 => x"C0C0C0F9F8C080B0",
 17084 => x"C0C0C0F9F8C08099",
 17085 => x"C0C0C0F9F8C08092",
 17086 => x"C0C0C0F9F8C08082",
 17087 => x"C0C0C0F9F8C080F8",
 17088 => x"C0C0C0F9F8C08080",
 17089 => x"C0C0C0F9F8C08090",
 17090 => x"C0C0C0F9F8C090C0",
 17091 => x"C0C0C0F9F8C090F9",
 17092 => x"C0C0C0F9F8C090A4",
 17093 => x"C0C0C0F9F8C090B0",
 17094 => x"C0C0C0F9F8C09099",
 17095 => x"C0C0C0F9F8C09092",
 17096 => x"C0C0C0F9F8C09082",
 17097 => x"C0C0C0F9F8C090F8",
 17098 => x"C0C0C0F9F8C09080",
 17099 => x"C0C0C0F9F8C09090",
 17100 => x"C0C0C0F9F8F9C0C0",
 17101 => x"C0C0C0F9F8F9C0F9",
 17102 => x"C0C0C0F9F8F9C0A4",
 17103 => x"C0C0C0F9F8F9C0B0",
 17104 => x"C0C0C0F9F8F9C099",
 17105 => x"C0C0C0F9F8F9C092",
 17106 => x"C0C0C0F9F8F9C082",
 17107 => x"C0C0C0F9F8F9C0F8",
 17108 => x"C0C0C0F9F8F9C080",
 17109 => x"C0C0C0F9F8F9C090",
 17110 => x"C0C0C0F9F8F9F9C0",
 17111 => x"C0C0C0F9F8F9F9F9",
 17112 => x"C0C0C0F9F8F9F9A4",
 17113 => x"C0C0C0F9F8F9F9B0",
 17114 => x"C0C0C0F9F8F9F999",
 17115 => x"C0C0C0F9F8F9F992",
 17116 => x"C0C0C0F9F8F9F982",
 17117 => x"C0C0C0F9F8F9F9F8",
 17118 => x"C0C0C0F9F8F9F980",
 17119 => x"C0C0C0F9F8F9F990",
 17120 => x"C0C0C0F9F8F9A4C0",
 17121 => x"C0C0C0F9F8F9A4F9",
 17122 => x"C0C0C0F9F8F9A4A4",
 17123 => x"C0C0C0F9F8F9A4B0",
 17124 => x"C0C0C0F9F8F9A499",
 17125 => x"C0C0C0F9F8F9A492",
 17126 => x"C0C0C0F9F8F9A482",
 17127 => x"C0C0C0F9F8F9A4F8",
 17128 => x"C0C0C0F9F8F9A480",
 17129 => x"C0C0C0F9F8F9A490",
 17130 => x"C0C0C0F9F8F9B0C0",
 17131 => x"C0C0C0F9F8F9B0F9",
 17132 => x"C0C0C0F9F8F9B0A4",
 17133 => x"C0C0C0F9F8F9B0B0",
 17134 => x"C0C0C0F9F8F9B099",
 17135 => x"C0C0C0F9F8F9B092",
 17136 => x"C0C0C0F9F8F9B082",
 17137 => x"C0C0C0F9F8F9B0F8",
 17138 => x"C0C0C0F9F8F9B080",
 17139 => x"C0C0C0F9F8F9B090",
 17140 => x"C0C0C0F9F8F999C0",
 17141 => x"C0C0C0F9F8F999F9",
 17142 => x"C0C0C0F9F8F999A4",
 17143 => x"C0C0C0F9F8F999B0",
 17144 => x"C0C0C0F9F8F99999",
 17145 => x"C0C0C0F9F8F99992",
 17146 => x"C0C0C0F9F8F99982",
 17147 => x"C0C0C0F9F8F999F8",
 17148 => x"C0C0C0F9F8F99980",
 17149 => x"C0C0C0F9F8F99990",
 17150 => x"C0C0C0F9F8F992C0",
 17151 => x"C0C0C0F9F8F992F9",
 17152 => x"C0C0C0F9F8F992A4",
 17153 => x"C0C0C0F9F8F992B0",
 17154 => x"C0C0C0F9F8F99299",
 17155 => x"C0C0C0F9F8F99292",
 17156 => x"C0C0C0F9F8F99282",
 17157 => x"C0C0C0F9F8F992F8",
 17158 => x"C0C0C0F9F8F99280",
 17159 => x"C0C0C0F9F8F99290",
 17160 => x"C0C0C0F9F8F982C0",
 17161 => x"C0C0C0F9F8F982F9",
 17162 => x"C0C0C0F9F8F982A4",
 17163 => x"C0C0C0F9F8F982B0",
 17164 => x"C0C0C0F9F8F98299",
 17165 => x"C0C0C0F9F8F98292",
 17166 => x"C0C0C0F9F8F98282",
 17167 => x"C0C0C0F9F8F982F8",
 17168 => x"C0C0C0F9F8F98280",
 17169 => x"C0C0C0F9F8F98290",
 17170 => x"C0C0C0F9F8F9F8C0",
 17171 => x"C0C0C0F9F8F9F8F9",
 17172 => x"C0C0C0F9F8F9F8A4",
 17173 => x"C0C0C0F9F8F9F8B0",
 17174 => x"C0C0C0F9F8F9F899",
 17175 => x"C0C0C0F9F8F9F892",
 17176 => x"C0C0C0F9F8F9F882",
 17177 => x"C0C0C0F9F8F9F8F8",
 17178 => x"C0C0C0F9F8F9F880",
 17179 => x"C0C0C0F9F8F9F890",
 17180 => x"C0C0C0F9F8F980C0",
 17181 => x"C0C0C0F9F8F980F9",
 17182 => x"C0C0C0F9F8F980A4",
 17183 => x"C0C0C0F9F8F980B0",
 17184 => x"C0C0C0F9F8F98099",
 17185 => x"C0C0C0F9F8F98092",
 17186 => x"C0C0C0F9F8F98082",
 17187 => x"C0C0C0F9F8F980F8",
 17188 => x"C0C0C0F9F8F98080",
 17189 => x"C0C0C0F9F8F98090",
 17190 => x"C0C0C0F9F8F990C0",
 17191 => x"C0C0C0F9F8F990F9",
 17192 => x"C0C0C0F9F8F990A4",
 17193 => x"C0C0C0F9F8F990B0",
 17194 => x"C0C0C0F9F8F99099",
 17195 => x"C0C0C0F9F8F99092",
 17196 => x"C0C0C0F9F8F99082",
 17197 => x"C0C0C0F9F8F990F8",
 17198 => x"C0C0C0F9F8F99080",
 17199 => x"C0C0C0F9F8F99090",
 17200 => x"C0C0C0F9F8A4C0C0",
 17201 => x"C0C0C0F9F8A4C0F9",
 17202 => x"C0C0C0F9F8A4C0A4",
 17203 => x"C0C0C0F9F8A4C0B0",
 17204 => x"C0C0C0F9F8A4C099",
 17205 => x"C0C0C0F9F8A4C092",
 17206 => x"C0C0C0F9F8A4C082",
 17207 => x"C0C0C0F9F8A4C0F8",
 17208 => x"C0C0C0F9F8A4C080",
 17209 => x"C0C0C0F9F8A4C090",
 17210 => x"C0C0C0F9F8A4F9C0",
 17211 => x"C0C0C0F9F8A4F9F9",
 17212 => x"C0C0C0F9F8A4F9A4",
 17213 => x"C0C0C0F9F8A4F9B0",
 17214 => x"C0C0C0F9F8A4F999",
 17215 => x"C0C0C0F9F8A4F992",
 17216 => x"C0C0C0F9F8A4F982",
 17217 => x"C0C0C0F9F8A4F9F8",
 17218 => x"C0C0C0F9F8A4F980",
 17219 => x"C0C0C0F9F8A4F990",
 17220 => x"C0C0C0F9F8A4A4C0",
 17221 => x"C0C0C0F9F8A4A4F9",
 17222 => x"C0C0C0F9F8A4A4A4",
 17223 => x"C0C0C0F9F8A4A4B0",
 17224 => x"C0C0C0F9F8A4A499",
 17225 => x"C0C0C0F9F8A4A492",
 17226 => x"C0C0C0F9F8A4A482",
 17227 => x"C0C0C0F9F8A4A4F8",
 17228 => x"C0C0C0F9F8A4A480",
 17229 => x"C0C0C0F9F8A4A490",
 17230 => x"C0C0C0F9F8A4B0C0",
 17231 => x"C0C0C0F9F8A4B0F9",
 17232 => x"C0C0C0F9F8A4B0A4",
 17233 => x"C0C0C0F9F8A4B0B0",
 17234 => x"C0C0C0F9F8A4B099",
 17235 => x"C0C0C0F9F8A4B092",
 17236 => x"C0C0C0F9F8A4B082",
 17237 => x"C0C0C0F9F8A4B0F8",
 17238 => x"C0C0C0F9F8A4B080",
 17239 => x"C0C0C0F9F8A4B090",
 17240 => x"C0C0C0F9F8A499C0",
 17241 => x"C0C0C0F9F8A499F9",
 17242 => x"C0C0C0F9F8A499A4",
 17243 => x"C0C0C0F9F8A499B0",
 17244 => x"C0C0C0F9F8A49999",
 17245 => x"C0C0C0F9F8A49992",
 17246 => x"C0C0C0F9F8A49982",
 17247 => x"C0C0C0F9F8A499F8",
 17248 => x"C0C0C0F9F8A49980",
 17249 => x"C0C0C0F9F8A49990",
 17250 => x"C0C0C0F9F8A492C0",
 17251 => x"C0C0C0F9F8A492F9",
 17252 => x"C0C0C0F9F8A492A4",
 17253 => x"C0C0C0F9F8A492B0",
 17254 => x"C0C0C0F9F8A49299",
 17255 => x"C0C0C0F9F8A49292",
 17256 => x"C0C0C0F9F8A49282",
 17257 => x"C0C0C0F9F8A492F8",
 17258 => x"C0C0C0F9F8A49280",
 17259 => x"C0C0C0F9F8A49290",
 17260 => x"C0C0C0F9F8A482C0",
 17261 => x"C0C0C0F9F8A482F9",
 17262 => x"C0C0C0F9F8A482A4",
 17263 => x"C0C0C0F9F8A482B0",
 17264 => x"C0C0C0F9F8A48299",
 17265 => x"C0C0C0F9F8A48292",
 17266 => x"C0C0C0F9F8A48282",
 17267 => x"C0C0C0F9F8A482F8",
 17268 => x"C0C0C0F9F8A48280",
 17269 => x"C0C0C0F9F8A48290",
 17270 => x"C0C0C0F9F8A4F8C0",
 17271 => x"C0C0C0F9F8A4F8F9",
 17272 => x"C0C0C0F9F8A4F8A4",
 17273 => x"C0C0C0F9F8A4F8B0",
 17274 => x"C0C0C0F9F8A4F899",
 17275 => x"C0C0C0F9F8A4F892",
 17276 => x"C0C0C0F9F8A4F882",
 17277 => x"C0C0C0F9F8A4F8F8",
 17278 => x"C0C0C0F9F8A4F880",
 17279 => x"C0C0C0F9F8A4F890",
 17280 => x"C0C0C0F9F8A480C0",
 17281 => x"C0C0C0F9F8A480F9",
 17282 => x"C0C0C0F9F8A480A4",
 17283 => x"C0C0C0F9F8A480B0",
 17284 => x"C0C0C0F9F8A48099",
 17285 => x"C0C0C0F9F8A48092",
 17286 => x"C0C0C0F9F8A48082",
 17287 => x"C0C0C0F9F8A480F8",
 17288 => x"C0C0C0F9F8A48080",
 17289 => x"C0C0C0F9F8A48090",
 17290 => x"C0C0C0F9F8A490C0",
 17291 => x"C0C0C0F9F8A490F9",
 17292 => x"C0C0C0F9F8A490A4",
 17293 => x"C0C0C0F9F8A490B0",
 17294 => x"C0C0C0F9F8A49099",
 17295 => x"C0C0C0F9F8A49092",
 17296 => x"C0C0C0F9F8A49082",
 17297 => x"C0C0C0F9F8A490F8",
 17298 => x"C0C0C0F9F8A49080",
 17299 => x"C0C0C0F9F8A49090",
 17300 => x"C0C0C0F9F8B0C0C0",
 17301 => x"C0C0C0F9F8B0C0F9",
 17302 => x"C0C0C0F9F8B0C0A4",
 17303 => x"C0C0C0F9F8B0C0B0",
 17304 => x"C0C0C0F9F8B0C099",
 17305 => x"C0C0C0F9F8B0C092",
 17306 => x"C0C0C0F9F8B0C082",
 17307 => x"C0C0C0F9F8B0C0F8",
 17308 => x"C0C0C0F9F8B0C080",
 17309 => x"C0C0C0F9F8B0C090",
 17310 => x"C0C0C0F9F8B0F9C0",
 17311 => x"C0C0C0F9F8B0F9F9",
 17312 => x"C0C0C0F9F8B0F9A4",
 17313 => x"C0C0C0F9F8B0F9B0",
 17314 => x"C0C0C0F9F8B0F999",
 17315 => x"C0C0C0F9F8B0F992",
 17316 => x"C0C0C0F9F8B0F982",
 17317 => x"C0C0C0F9F8B0F9F8",
 17318 => x"C0C0C0F9F8B0F980",
 17319 => x"C0C0C0F9F8B0F990",
 17320 => x"C0C0C0F9F8B0A4C0",
 17321 => x"C0C0C0F9F8B0A4F9",
 17322 => x"C0C0C0F9F8B0A4A4",
 17323 => x"C0C0C0F9F8B0A4B0",
 17324 => x"C0C0C0F9F8B0A499",
 17325 => x"C0C0C0F9F8B0A492",
 17326 => x"C0C0C0F9F8B0A482",
 17327 => x"C0C0C0F9F8B0A4F8",
 17328 => x"C0C0C0F9F8B0A480",
 17329 => x"C0C0C0F9F8B0A490",
 17330 => x"C0C0C0F9F8B0B0C0",
 17331 => x"C0C0C0F9F8B0B0F9",
 17332 => x"C0C0C0F9F8B0B0A4",
 17333 => x"C0C0C0F9F8B0B0B0",
 17334 => x"C0C0C0F9F8B0B099",
 17335 => x"C0C0C0F9F8B0B092",
 17336 => x"C0C0C0F9F8B0B082",
 17337 => x"C0C0C0F9F8B0B0F8",
 17338 => x"C0C0C0F9F8B0B080",
 17339 => x"C0C0C0F9F8B0B090",
 17340 => x"C0C0C0F9F8B099C0",
 17341 => x"C0C0C0F9F8B099F9",
 17342 => x"C0C0C0F9F8B099A4",
 17343 => x"C0C0C0F9F8B099B0",
 17344 => x"C0C0C0F9F8B09999",
 17345 => x"C0C0C0F9F8B09992",
 17346 => x"C0C0C0F9F8B09982",
 17347 => x"C0C0C0F9F8B099F8",
 17348 => x"C0C0C0F9F8B09980",
 17349 => x"C0C0C0F9F8B09990",
 17350 => x"C0C0C0F9F8B092C0",
 17351 => x"C0C0C0F9F8B092F9",
 17352 => x"C0C0C0F9F8B092A4",
 17353 => x"C0C0C0F9F8B092B0",
 17354 => x"C0C0C0F9F8B09299",
 17355 => x"C0C0C0F9F8B09292",
 17356 => x"C0C0C0F9F8B09282",
 17357 => x"C0C0C0F9F8B092F8",
 17358 => x"C0C0C0F9F8B09280",
 17359 => x"C0C0C0F9F8B09290",
 17360 => x"C0C0C0F9F8B082C0",
 17361 => x"C0C0C0F9F8B082F9",
 17362 => x"C0C0C0F9F8B082A4",
 17363 => x"C0C0C0F9F8B082B0",
 17364 => x"C0C0C0F9F8B08299",
 17365 => x"C0C0C0F9F8B08292",
 17366 => x"C0C0C0F9F8B08282",
 17367 => x"C0C0C0F9F8B082F8",
 17368 => x"C0C0C0F9F8B08280",
 17369 => x"C0C0C0F9F8B08290",
 17370 => x"C0C0C0F9F8B0F8C0",
 17371 => x"C0C0C0F9F8B0F8F9",
 17372 => x"C0C0C0F9F8B0F8A4",
 17373 => x"C0C0C0F9F8B0F8B0",
 17374 => x"C0C0C0F9F8B0F899",
 17375 => x"C0C0C0F9F8B0F892",
 17376 => x"C0C0C0F9F8B0F882",
 17377 => x"C0C0C0F9F8B0F8F8",
 17378 => x"C0C0C0F9F8B0F880",
 17379 => x"C0C0C0F9F8B0F890",
 17380 => x"C0C0C0F9F8B080C0",
 17381 => x"C0C0C0F9F8B080F9",
 17382 => x"C0C0C0F9F8B080A4",
 17383 => x"C0C0C0F9F8B080B0",
 17384 => x"C0C0C0F9F8B08099",
 17385 => x"C0C0C0F9F8B08092",
 17386 => x"C0C0C0F9F8B08082",
 17387 => x"C0C0C0F9F8B080F8",
 17388 => x"C0C0C0F9F8B08080",
 17389 => x"C0C0C0F9F8B08090",
 17390 => x"C0C0C0F9F8B090C0",
 17391 => x"C0C0C0F9F8B090F9",
 17392 => x"C0C0C0F9F8B090A4",
 17393 => x"C0C0C0F9F8B090B0",
 17394 => x"C0C0C0F9F8B09099",
 17395 => x"C0C0C0F9F8B09092",
 17396 => x"C0C0C0F9F8B09082",
 17397 => x"C0C0C0F9F8B090F8",
 17398 => x"C0C0C0F9F8B09080",
 17399 => x"C0C0C0F9F8B09090",
 17400 => x"C0C0C0F9F899C0C0",
 17401 => x"C0C0C0F9F899C0F9",
 17402 => x"C0C0C0F9F899C0A4",
 17403 => x"C0C0C0F9F899C0B0",
 17404 => x"C0C0C0F9F899C099",
 17405 => x"C0C0C0F9F899C092",
 17406 => x"C0C0C0F9F899C082",
 17407 => x"C0C0C0F9F899C0F8",
 17408 => x"C0C0C0F9F899C080",
 17409 => x"C0C0C0F9F899C090",
 17410 => x"C0C0C0F9F899F9C0",
 17411 => x"C0C0C0F9F899F9F9",
 17412 => x"C0C0C0F9F899F9A4",
 17413 => x"C0C0C0F9F899F9B0",
 17414 => x"C0C0C0F9F899F999",
 17415 => x"C0C0C0F9F899F992",
 17416 => x"C0C0C0F9F899F982",
 17417 => x"C0C0C0F9F899F9F8",
 17418 => x"C0C0C0F9F899F980",
 17419 => x"C0C0C0F9F899F990",
 17420 => x"C0C0C0F9F899A4C0",
 17421 => x"C0C0C0F9F899A4F9",
 17422 => x"C0C0C0F9F899A4A4",
 17423 => x"C0C0C0F9F899A4B0",
 17424 => x"C0C0C0F9F899A499",
 17425 => x"C0C0C0F9F899A492",
 17426 => x"C0C0C0F9F899A482",
 17427 => x"C0C0C0F9F899A4F8",
 17428 => x"C0C0C0F9F899A480",
 17429 => x"C0C0C0F9F899A490",
 17430 => x"C0C0C0F9F899B0C0",
 17431 => x"C0C0C0F9F899B0F9",
 17432 => x"C0C0C0F9F899B0A4",
 17433 => x"C0C0C0F9F899B0B0",
 17434 => x"C0C0C0F9F899B099",
 17435 => x"C0C0C0F9F899B092",
 17436 => x"C0C0C0F9F899B082",
 17437 => x"C0C0C0F9F899B0F8",
 17438 => x"C0C0C0F9F899B080",
 17439 => x"C0C0C0F9F899B090",
 17440 => x"C0C0C0F9F89999C0",
 17441 => x"C0C0C0F9F89999F9",
 17442 => x"C0C0C0F9F89999A4",
 17443 => x"C0C0C0F9F89999B0",
 17444 => x"C0C0C0F9F8999999",
 17445 => x"C0C0C0F9F8999992",
 17446 => x"C0C0C0F9F8999982",
 17447 => x"C0C0C0F9F89999F8",
 17448 => x"C0C0C0F9F8999980",
 17449 => x"C0C0C0F9F8999990",
 17450 => x"C0C0C0F9F89992C0",
 17451 => x"C0C0C0F9F89992F9",
 17452 => x"C0C0C0F9F89992A4",
 17453 => x"C0C0C0F9F89992B0",
 17454 => x"C0C0C0F9F8999299",
 17455 => x"C0C0C0F9F8999292",
 17456 => x"C0C0C0F9F8999282",
 17457 => x"C0C0C0F9F89992F8",
 17458 => x"C0C0C0F9F8999280",
 17459 => x"C0C0C0F9F8999290",
 17460 => x"C0C0C0F9F89982C0",
 17461 => x"C0C0C0F9F89982F9",
 17462 => x"C0C0C0F9F89982A4",
 17463 => x"C0C0C0F9F89982B0",
 17464 => x"C0C0C0F9F8998299",
 17465 => x"C0C0C0F9F8998292",
 17466 => x"C0C0C0F9F8998282",
 17467 => x"C0C0C0F9F89982F8",
 17468 => x"C0C0C0F9F8998280",
 17469 => x"C0C0C0F9F8998290",
 17470 => x"C0C0C0F9F899F8C0",
 17471 => x"C0C0C0F9F899F8F9",
 17472 => x"C0C0C0F9F899F8A4",
 17473 => x"C0C0C0F9F899F8B0",
 17474 => x"C0C0C0F9F899F899",
 17475 => x"C0C0C0F9F899F892",
 17476 => x"C0C0C0F9F899F882",
 17477 => x"C0C0C0F9F899F8F8",
 17478 => x"C0C0C0F9F899F880",
 17479 => x"C0C0C0F9F899F890",
 17480 => x"C0C0C0F9F89980C0",
 17481 => x"C0C0C0F9F89980F9",
 17482 => x"C0C0C0F9F89980A4",
 17483 => x"C0C0C0F9F89980B0",
 17484 => x"C0C0C0F9F8998099",
 17485 => x"C0C0C0F9F8998092",
 17486 => x"C0C0C0F9F8998082",
 17487 => x"C0C0C0F9F89980F8",
 17488 => x"C0C0C0F9F8998080",
 17489 => x"C0C0C0F9F8998090",
 17490 => x"C0C0C0F9F89990C0",
 17491 => x"C0C0C0F9F89990F9",
 17492 => x"C0C0C0F9F89990A4",
 17493 => x"C0C0C0F9F89990B0",
 17494 => x"C0C0C0F9F8999099",
 17495 => x"C0C0C0F9F8999092",
 17496 => x"C0C0C0F9F8999082",
 17497 => x"C0C0C0F9F89990F8",
 17498 => x"C0C0C0F9F8999080",
 17499 => x"C0C0C0F9F8999090",
 17500 => x"C0C0C0F9F892C0C0",
 17501 => x"C0C0C0F9F892C0F9",
 17502 => x"C0C0C0F9F892C0A4",
 17503 => x"C0C0C0F9F892C0B0",
 17504 => x"C0C0C0F9F892C099",
 17505 => x"C0C0C0F9F892C092",
 17506 => x"C0C0C0F9F892C082",
 17507 => x"C0C0C0F9F892C0F8",
 17508 => x"C0C0C0F9F892C080",
 17509 => x"C0C0C0F9F892C090",
 17510 => x"C0C0C0F9F892F9C0",
 17511 => x"C0C0C0F9F892F9F9",
 17512 => x"C0C0C0F9F892F9A4",
 17513 => x"C0C0C0F9F892F9B0",
 17514 => x"C0C0C0F9F892F999",
 17515 => x"C0C0C0F9F892F992",
 17516 => x"C0C0C0F9F892F982",
 17517 => x"C0C0C0F9F892F9F8",
 17518 => x"C0C0C0F9F892F980",
 17519 => x"C0C0C0F9F892F990",
 17520 => x"C0C0C0F9F892A4C0",
 17521 => x"C0C0C0F9F892A4F9",
 17522 => x"C0C0C0F9F892A4A4",
 17523 => x"C0C0C0F9F892A4B0",
 17524 => x"C0C0C0F9F892A499",
 17525 => x"C0C0C0F9F892A492",
 17526 => x"C0C0C0F9F892A482",
 17527 => x"C0C0C0F9F892A4F8",
 17528 => x"C0C0C0F9F892A480",
 17529 => x"C0C0C0F9F892A490",
 17530 => x"C0C0C0F9F892B0C0",
 17531 => x"C0C0C0F9F892B0F9",
 17532 => x"C0C0C0F9F892B0A4",
 17533 => x"C0C0C0F9F892B0B0",
 17534 => x"C0C0C0F9F892B099",
 17535 => x"C0C0C0F9F892B092",
 17536 => x"C0C0C0F9F892B082",
 17537 => x"C0C0C0F9F892B0F8",
 17538 => x"C0C0C0F9F892B080",
 17539 => x"C0C0C0F9F892B090",
 17540 => x"C0C0C0F9F89299C0",
 17541 => x"C0C0C0F9F89299F9",
 17542 => x"C0C0C0F9F89299A4",
 17543 => x"C0C0C0F9F89299B0",
 17544 => x"C0C0C0F9F8929999",
 17545 => x"C0C0C0F9F8929992",
 17546 => x"C0C0C0F9F8929982",
 17547 => x"C0C0C0F9F89299F8",
 17548 => x"C0C0C0F9F8929980",
 17549 => x"C0C0C0F9F8929990",
 17550 => x"C0C0C0F9F89292C0",
 17551 => x"C0C0C0F9F89292F9",
 17552 => x"C0C0C0F9F89292A4",
 17553 => x"C0C0C0F9F89292B0",
 17554 => x"C0C0C0F9F8929299",
 17555 => x"C0C0C0F9F8929292",
 17556 => x"C0C0C0F9F8929282",
 17557 => x"C0C0C0F9F89292F8",
 17558 => x"C0C0C0F9F8929280",
 17559 => x"C0C0C0F9F8929290",
 17560 => x"C0C0C0F9F89282C0",
 17561 => x"C0C0C0F9F89282F9",
 17562 => x"C0C0C0F9F89282A4",
 17563 => x"C0C0C0F9F89282B0",
 17564 => x"C0C0C0F9F8928299",
 17565 => x"C0C0C0F9F8928292",
 17566 => x"C0C0C0F9F8928282",
 17567 => x"C0C0C0F9F89282F8",
 17568 => x"C0C0C0F9F8928280",
 17569 => x"C0C0C0F9F8928290",
 17570 => x"C0C0C0F9F892F8C0",
 17571 => x"C0C0C0F9F892F8F9",
 17572 => x"C0C0C0F9F892F8A4",
 17573 => x"C0C0C0F9F892F8B0",
 17574 => x"C0C0C0F9F892F899",
 17575 => x"C0C0C0F9F892F892",
 17576 => x"C0C0C0F9F892F882",
 17577 => x"C0C0C0F9F892F8F8",
 17578 => x"C0C0C0F9F892F880",
 17579 => x"C0C0C0F9F892F890",
 17580 => x"C0C0C0F9F89280C0",
 17581 => x"C0C0C0F9F89280F9",
 17582 => x"C0C0C0F9F89280A4",
 17583 => x"C0C0C0F9F89280B0",
 17584 => x"C0C0C0F9F8928099",
 17585 => x"C0C0C0F9F8928092",
 17586 => x"C0C0C0F9F8928082",
 17587 => x"C0C0C0F9F89280F8",
 17588 => x"C0C0C0F9F8928080",
 17589 => x"C0C0C0F9F8928090",
 17590 => x"C0C0C0F9F89290C0",
 17591 => x"C0C0C0F9F89290F9",
 17592 => x"C0C0C0F9F89290A4",
 17593 => x"C0C0C0F9F89290B0",
 17594 => x"C0C0C0F9F8929099",
 17595 => x"C0C0C0F9F8929092",
 17596 => x"C0C0C0F9F8929082",
 17597 => x"C0C0C0F9F89290F8",
 17598 => x"C0C0C0F9F8929080",
 17599 => x"C0C0C0F9F8929090",
 17600 => x"C0C0C0F9F882C0C0",
 17601 => x"C0C0C0F9F882C0F9",
 17602 => x"C0C0C0F9F882C0A4",
 17603 => x"C0C0C0F9F882C0B0",
 17604 => x"C0C0C0F9F882C099",
 17605 => x"C0C0C0F9F882C092",
 17606 => x"C0C0C0F9F882C082",
 17607 => x"C0C0C0F9F882C0F8",
 17608 => x"C0C0C0F9F882C080",
 17609 => x"C0C0C0F9F882C090",
 17610 => x"C0C0C0F9F882F9C0",
 17611 => x"C0C0C0F9F882F9F9",
 17612 => x"C0C0C0F9F882F9A4",
 17613 => x"C0C0C0F9F882F9B0",
 17614 => x"C0C0C0F9F882F999",
 17615 => x"C0C0C0F9F882F992",
 17616 => x"C0C0C0F9F882F982",
 17617 => x"C0C0C0F9F882F9F8",
 17618 => x"C0C0C0F9F882F980",
 17619 => x"C0C0C0F9F882F990",
 17620 => x"C0C0C0F9F882A4C0",
 17621 => x"C0C0C0F9F882A4F9",
 17622 => x"C0C0C0F9F882A4A4",
 17623 => x"C0C0C0F9F882A4B0",
 17624 => x"C0C0C0F9F882A499",
 17625 => x"C0C0C0F9F882A492",
 17626 => x"C0C0C0F9F882A482",
 17627 => x"C0C0C0F9F882A4F8",
 17628 => x"C0C0C0F9F882A480",
 17629 => x"C0C0C0F9F882A490",
 17630 => x"C0C0C0F9F882B0C0",
 17631 => x"C0C0C0F9F882B0F9",
 17632 => x"C0C0C0F9F882B0A4",
 17633 => x"C0C0C0F9F882B0B0",
 17634 => x"C0C0C0F9F882B099",
 17635 => x"C0C0C0F9F882B092",
 17636 => x"C0C0C0F9F882B082",
 17637 => x"C0C0C0F9F882B0F8",
 17638 => x"C0C0C0F9F882B080",
 17639 => x"C0C0C0F9F882B090",
 17640 => x"C0C0C0F9F88299C0",
 17641 => x"C0C0C0F9F88299F9",
 17642 => x"C0C0C0F9F88299A4",
 17643 => x"C0C0C0F9F88299B0",
 17644 => x"C0C0C0F9F8829999",
 17645 => x"C0C0C0F9F8829992",
 17646 => x"C0C0C0F9F8829982",
 17647 => x"C0C0C0F9F88299F8",
 17648 => x"C0C0C0F9F8829980",
 17649 => x"C0C0C0F9F8829990",
 17650 => x"C0C0C0F9F88292C0",
 17651 => x"C0C0C0F9F88292F9",
 17652 => x"C0C0C0F9F88292A4",
 17653 => x"C0C0C0F9F88292B0",
 17654 => x"C0C0C0F9F8829299",
 17655 => x"C0C0C0F9F8829292",
 17656 => x"C0C0C0F9F8829282",
 17657 => x"C0C0C0F9F88292F8",
 17658 => x"C0C0C0F9F8829280",
 17659 => x"C0C0C0F9F8829290",
 17660 => x"C0C0C0F9F88282C0",
 17661 => x"C0C0C0F9F88282F9",
 17662 => x"C0C0C0F9F88282A4",
 17663 => x"C0C0C0F9F88282B0",
 17664 => x"C0C0C0F9F8828299",
 17665 => x"C0C0C0F9F8828292",
 17666 => x"C0C0C0F9F8828282",
 17667 => x"C0C0C0F9F88282F8",
 17668 => x"C0C0C0F9F8828280",
 17669 => x"C0C0C0F9F8828290",
 17670 => x"C0C0C0F9F882F8C0",
 17671 => x"C0C0C0F9F882F8F9",
 17672 => x"C0C0C0F9F882F8A4",
 17673 => x"C0C0C0F9F882F8B0",
 17674 => x"C0C0C0F9F882F899",
 17675 => x"C0C0C0F9F882F892",
 17676 => x"C0C0C0F9F882F882",
 17677 => x"C0C0C0F9F882F8F8",
 17678 => x"C0C0C0F9F882F880",
 17679 => x"C0C0C0F9F882F890",
 17680 => x"C0C0C0F9F88280C0",
 17681 => x"C0C0C0F9F88280F9",
 17682 => x"C0C0C0F9F88280A4",
 17683 => x"C0C0C0F9F88280B0",
 17684 => x"C0C0C0F9F8828099",
 17685 => x"C0C0C0F9F8828092",
 17686 => x"C0C0C0F9F8828082",
 17687 => x"C0C0C0F9F88280F8",
 17688 => x"C0C0C0F9F8828080",
 17689 => x"C0C0C0F9F8828090",
 17690 => x"C0C0C0F9F88290C0",
 17691 => x"C0C0C0F9F88290F9",
 17692 => x"C0C0C0F9F88290A4",
 17693 => x"C0C0C0F9F88290B0",
 17694 => x"C0C0C0F9F8829099",
 17695 => x"C0C0C0F9F8829092",
 17696 => x"C0C0C0F9F8829082",
 17697 => x"C0C0C0F9F88290F8",
 17698 => x"C0C0C0F9F8829080",
 17699 => x"C0C0C0F9F8829090",
 17700 => x"C0C0C0F9F8F8C0C0",
 17701 => x"C0C0C0F9F8F8C0F9",
 17702 => x"C0C0C0F9F8F8C0A4",
 17703 => x"C0C0C0F9F8F8C0B0",
 17704 => x"C0C0C0F9F8F8C099",
 17705 => x"C0C0C0F9F8F8C092",
 17706 => x"C0C0C0F9F8F8C082",
 17707 => x"C0C0C0F9F8F8C0F8",
 17708 => x"C0C0C0F9F8F8C080",
 17709 => x"C0C0C0F9F8F8C090",
 17710 => x"C0C0C0F9F8F8F9C0",
 17711 => x"C0C0C0F9F8F8F9F9",
 17712 => x"C0C0C0F9F8F8F9A4",
 17713 => x"C0C0C0F9F8F8F9B0",
 17714 => x"C0C0C0F9F8F8F999",
 17715 => x"C0C0C0F9F8F8F992",
 17716 => x"C0C0C0F9F8F8F982",
 17717 => x"C0C0C0F9F8F8F9F8",
 17718 => x"C0C0C0F9F8F8F980",
 17719 => x"C0C0C0F9F8F8F990",
 17720 => x"C0C0C0F9F8F8A4C0",
 17721 => x"C0C0C0F9F8F8A4F9",
 17722 => x"C0C0C0F9F8F8A4A4",
 17723 => x"C0C0C0F9F8F8A4B0",
 17724 => x"C0C0C0F9F8F8A499",
 17725 => x"C0C0C0F9F8F8A492",
 17726 => x"C0C0C0F9F8F8A482",
 17727 => x"C0C0C0F9F8F8A4F8",
 17728 => x"C0C0C0F9F8F8A480",
 17729 => x"C0C0C0F9F8F8A490",
 17730 => x"C0C0C0F9F8F8B0C0",
 17731 => x"C0C0C0F9F8F8B0F9",
 17732 => x"C0C0C0F9F8F8B0A4",
 17733 => x"C0C0C0F9F8F8B0B0",
 17734 => x"C0C0C0F9F8F8B099",
 17735 => x"C0C0C0F9F8F8B092",
 17736 => x"C0C0C0F9F8F8B082",
 17737 => x"C0C0C0F9F8F8B0F8",
 17738 => x"C0C0C0F9F8F8B080",
 17739 => x"C0C0C0F9F8F8B090",
 17740 => x"C0C0C0F9F8F899C0",
 17741 => x"C0C0C0F9F8F899F9",
 17742 => x"C0C0C0F9F8F899A4",
 17743 => x"C0C0C0F9F8F899B0",
 17744 => x"C0C0C0F9F8F89999",
 17745 => x"C0C0C0F9F8F89992",
 17746 => x"C0C0C0F9F8F89982",
 17747 => x"C0C0C0F9F8F899F8",
 17748 => x"C0C0C0F9F8F89980",
 17749 => x"C0C0C0F9F8F89990",
 17750 => x"C0C0C0F9F8F892C0",
 17751 => x"C0C0C0F9F8F892F9",
 17752 => x"C0C0C0F9F8F892A4",
 17753 => x"C0C0C0F9F8F892B0",
 17754 => x"C0C0C0F9F8F89299",
 17755 => x"C0C0C0F9F8F89292",
 17756 => x"C0C0C0F9F8F89282",
 17757 => x"C0C0C0F9F8F892F8",
 17758 => x"C0C0C0F9F8F89280",
 17759 => x"C0C0C0F9F8F89290",
 17760 => x"C0C0C0F9F8F882C0",
 17761 => x"C0C0C0F9F8F882F9",
 17762 => x"C0C0C0F9F8F882A4",
 17763 => x"C0C0C0F9F8F882B0",
 17764 => x"C0C0C0F9F8F88299",
 17765 => x"C0C0C0F9F8F88292",
 17766 => x"C0C0C0F9F8F88282",
 17767 => x"C0C0C0F9F8F882F8",
 17768 => x"C0C0C0F9F8F88280",
 17769 => x"C0C0C0F9F8F88290",
 17770 => x"C0C0C0F9F8F8F8C0",
 17771 => x"C0C0C0F9F8F8F8F9",
 17772 => x"C0C0C0F9F8F8F8A4",
 17773 => x"C0C0C0F9F8F8F8B0",
 17774 => x"C0C0C0F9F8F8F899",
 17775 => x"C0C0C0F9F8F8F892",
 17776 => x"C0C0C0F9F8F8F882",
 17777 => x"C0C0C0F9F8F8F8F8",
 17778 => x"C0C0C0F9F8F8F880",
 17779 => x"C0C0C0F9F8F8F890",
 17780 => x"C0C0C0F9F8F880C0",
 17781 => x"C0C0C0F9F8F880F9",
 17782 => x"C0C0C0F9F8F880A4",
 17783 => x"C0C0C0F9F8F880B0",
 17784 => x"C0C0C0F9F8F88099",
 17785 => x"C0C0C0F9F8F88092",
 17786 => x"C0C0C0F9F8F88082",
 17787 => x"C0C0C0F9F8F880F8",
 17788 => x"C0C0C0F9F8F88080",
 17789 => x"C0C0C0F9F8F88090",
 17790 => x"C0C0C0F9F8F890C0",
 17791 => x"C0C0C0F9F8F890F9",
 17792 => x"C0C0C0F9F8F890A4",
 17793 => x"C0C0C0F9F8F890B0",
 17794 => x"C0C0C0F9F8F89099",
 17795 => x"C0C0C0F9F8F89092",
 17796 => x"C0C0C0F9F8F89082",
 17797 => x"C0C0C0F9F8F890F8",
 17798 => x"C0C0C0F9F8F89080",
 17799 => x"C0C0C0F9F8F89090",
 17800 => x"C0C0C0F9F880C0C0",
 17801 => x"C0C0C0F9F880C0F9",
 17802 => x"C0C0C0F9F880C0A4",
 17803 => x"C0C0C0F9F880C0B0",
 17804 => x"C0C0C0F9F880C099",
 17805 => x"C0C0C0F9F880C092",
 17806 => x"C0C0C0F9F880C082",
 17807 => x"C0C0C0F9F880C0F8",
 17808 => x"C0C0C0F9F880C080",
 17809 => x"C0C0C0F9F880C090",
 17810 => x"C0C0C0F9F880F9C0",
 17811 => x"C0C0C0F9F880F9F9",
 17812 => x"C0C0C0F9F880F9A4",
 17813 => x"C0C0C0F9F880F9B0",
 17814 => x"C0C0C0F9F880F999",
 17815 => x"C0C0C0F9F880F992",
 17816 => x"C0C0C0F9F880F982",
 17817 => x"C0C0C0F9F880F9F8",
 17818 => x"C0C0C0F9F880F980",
 17819 => x"C0C0C0F9F880F990",
 17820 => x"C0C0C0F9F880A4C0",
 17821 => x"C0C0C0F9F880A4F9",
 17822 => x"C0C0C0F9F880A4A4",
 17823 => x"C0C0C0F9F880A4B0",
 17824 => x"C0C0C0F9F880A499",
 17825 => x"C0C0C0F9F880A492",
 17826 => x"C0C0C0F9F880A482",
 17827 => x"C0C0C0F9F880A4F8",
 17828 => x"C0C0C0F9F880A480",
 17829 => x"C0C0C0F9F880A490",
 17830 => x"C0C0C0F9F880B0C0",
 17831 => x"C0C0C0F9F880B0F9",
 17832 => x"C0C0C0F9F880B0A4",
 17833 => x"C0C0C0F9F880B0B0",
 17834 => x"C0C0C0F9F880B099",
 17835 => x"C0C0C0F9F880B092",
 17836 => x"C0C0C0F9F880B082",
 17837 => x"C0C0C0F9F880B0F8",
 17838 => x"C0C0C0F9F880B080",
 17839 => x"C0C0C0F9F880B090",
 17840 => x"C0C0C0F9F88099C0",
 17841 => x"C0C0C0F9F88099F9",
 17842 => x"C0C0C0F9F88099A4",
 17843 => x"C0C0C0F9F88099B0",
 17844 => x"C0C0C0F9F8809999",
 17845 => x"C0C0C0F9F8809992",
 17846 => x"C0C0C0F9F8809982",
 17847 => x"C0C0C0F9F88099F8",
 17848 => x"C0C0C0F9F8809980",
 17849 => x"C0C0C0F9F8809990",
 17850 => x"C0C0C0F9F88092C0",
 17851 => x"C0C0C0F9F88092F9",
 17852 => x"C0C0C0F9F88092A4",
 17853 => x"C0C0C0F9F88092B0",
 17854 => x"C0C0C0F9F8809299",
 17855 => x"C0C0C0F9F8809292",
 17856 => x"C0C0C0F9F8809282",
 17857 => x"C0C0C0F9F88092F8",
 17858 => x"C0C0C0F9F8809280",
 17859 => x"C0C0C0F9F8809290",
 17860 => x"C0C0C0F9F88082C0",
 17861 => x"C0C0C0F9F88082F9",
 17862 => x"C0C0C0F9F88082A4",
 17863 => x"C0C0C0F9F88082B0",
 17864 => x"C0C0C0F9F8808299",
 17865 => x"C0C0C0F9F8808292",
 17866 => x"C0C0C0F9F8808282",
 17867 => x"C0C0C0F9F88082F8",
 17868 => x"C0C0C0F9F8808280",
 17869 => x"C0C0C0F9F8808290",
 17870 => x"C0C0C0F9F880F8C0",
 17871 => x"C0C0C0F9F880F8F9",
 17872 => x"C0C0C0F9F880F8A4",
 17873 => x"C0C0C0F9F880F8B0",
 17874 => x"C0C0C0F9F880F899",
 17875 => x"C0C0C0F9F880F892",
 17876 => x"C0C0C0F9F880F882",
 17877 => x"C0C0C0F9F880F8F8",
 17878 => x"C0C0C0F9F880F880",
 17879 => x"C0C0C0F9F880F890",
 17880 => x"C0C0C0F9F88080C0",
 17881 => x"C0C0C0F9F88080F9",
 17882 => x"C0C0C0F9F88080A4",
 17883 => x"C0C0C0F9F88080B0",
 17884 => x"C0C0C0F9F8808099",
 17885 => x"C0C0C0F9F8808092",
 17886 => x"C0C0C0F9F8808082",
 17887 => x"C0C0C0F9F88080F8",
 17888 => x"C0C0C0F9F8808080",
 17889 => x"C0C0C0F9F8808090",
 17890 => x"C0C0C0F9F88090C0",
 17891 => x"C0C0C0F9F88090F9",
 17892 => x"C0C0C0F9F88090A4",
 17893 => x"C0C0C0F9F88090B0",
 17894 => x"C0C0C0F9F8809099",
 17895 => x"C0C0C0F9F8809092",
 17896 => x"C0C0C0F9F8809082",
 17897 => x"C0C0C0F9F88090F8",
 17898 => x"C0C0C0F9F8809080",
 17899 => x"C0C0C0F9F8809090",
 17900 => x"C0C0C0F9F890C0C0",
 17901 => x"C0C0C0F9F890C0F9",
 17902 => x"C0C0C0F9F890C0A4",
 17903 => x"C0C0C0F9F890C0B0",
 17904 => x"C0C0C0F9F890C099",
 17905 => x"C0C0C0F9F890C092",
 17906 => x"C0C0C0F9F890C082",
 17907 => x"C0C0C0F9F890C0F8",
 17908 => x"C0C0C0F9F890C080",
 17909 => x"C0C0C0F9F890C090",
 17910 => x"C0C0C0F9F890F9C0",
 17911 => x"C0C0C0F9F890F9F9",
 17912 => x"C0C0C0F9F890F9A4",
 17913 => x"C0C0C0F9F890F9B0",
 17914 => x"C0C0C0F9F890F999",
 17915 => x"C0C0C0F9F890F992",
 17916 => x"C0C0C0F9F890F982",
 17917 => x"C0C0C0F9F890F9F8",
 17918 => x"C0C0C0F9F890F980",
 17919 => x"C0C0C0F9F890F990",
 17920 => x"C0C0C0F9F890A4C0",
 17921 => x"C0C0C0F9F890A4F9",
 17922 => x"C0C0C0F9F890A4A4",
 17923 => x"C0C0C0F9F890A4B0",
 17924 => x"C0C0C0F9F890A499",
 17925 => x"C0C0C0F9F890A492",
 17926 => x"C0C0C0F9F890A482",
 17927 => x"C0C0C0F9F890A4F8",
 17928 => x"C0C0C0F9F890A480",
 17929 => x"C0C0C0F9F890A490",
 17930 => x"C0C0C0F9F890B0C0",
 17931 => x"C0C0C0F9F890B0F9",
 17932 => x"C0C0C0F9F890B0A4",
 17933 => x"C0C0C0F9F890B0B0",
 17934 => x"C0C0C0F9F890B099",
 17935 => x"C0C0C0F9F890B092",
 17936 => x"C0C0C0F9F890B082",
 17937 => x"C0C0C0F9F890B0F8",
 17938 => x"C0C0C0F9F890B080",
 17939 => x"C0C0C0F9F890B090",
 17940 => x"C0C0C0F9F89099C0",
 17941 => x"C0C0C0F9F89099F9",
 17942 => x"C0C0C0F9F89099A4",
 17943 => x"C0C0C0F9F89099B0",
 17944 => x"C0C0C0F9F8909999",
 17945 => x"C0C0C0F9F8909992",
 17946 => x"C0C0C0F9F8909982",
 17947 => x"C0C0C0F9F89099F8",
 17948 => x"C0C0C0F9F8909980",
 17949 => x"C0C0C0F9F8909990",
 17950 => x"C0C0C0F9F89092C0",
 17951 => x"C0C0C0F9F89092F9",
 17952 => x"C0C0C0F9F89092A4",
 17953 => x"C0C0C0F9F89092B0",
 17954 => x"C0C0C0F9F8909299",
 17955 => x"C0C0C0F9F8909292",
 17956 => x"C0C0C0F9F8909282",
 17957 => x"C0C0C0F9F89092F8",
 17958 => x"C0C0C0F9F8909280",
 17959 => x"C0C0C0F9F8909290",
 17960 => x"C0C0C0F9F89082C0",
 17961 => x"C0C0C0F9F89082F9",
 17962 => x"C0C0C0F9F89082A4",
 17963 => x"C0C0C0F9F89082B0",
 17964 => x"C0C0C0F9F8908299",
 17965 => x"C0C0C0F9F8908292",
 17966 => x"C0C0C0F9F8908282",
 17967 => x"C0C0C0F9F89082F8",
 17968 => x"C0C0C0F9F8908280",
 17969 => x"C0C0C0F9F8908290",
 17970 => x"C0C0C0F9F890F8C0",
 17971 => x"C0C0C0F9F890F8F9",
 17972 => x"C0C0C0F9F890F8A4",
 17973 => x"C0C0C0F9F890F8B0",
 17974 => x"C0C0C0F9F890F899",
 17975 => x"C0C0C0F9F890F892",
 17976 => x"C0C0C0F9F890F882",
 17977 => x"C0C0C0F9F890F8F8",
 17978 => x"C0C0C0F9F890F880",
 17979 => x"C0C0C0F9F890F890",
 17980 => x"C0C0C0F9F89080C0",
 17981 => x"C0C0C0F9F89080F9",
 17982 => x"C0C0C0F9F89080A4",
 17983 => x"C0C0C0F9F89080B0",
 17984 => x"C0C0C0F9F8908099",
 17985 => x"C0C0C0F9F8908092",
 17986 => x"C0C0C0F9F8908082",
 17987 => x"C0C0C0F9F89080F8",
 17988 => x"C0C0C0F9F8908080",
 17989 => x"C0C0C0F9F8908090",
 17990 => x"C0C0C0F9F89090C0",
 17991 => x"C0C0C0F9F89090F9",
 17992 => x"C0C0C0F9F89090A4",
 17993 => x"C0C0C0F9F89090B0",
 17994 => x"C0C0C0F9F8909099",
 17995 => x"C0C0C0F9F8909092",
 17996 => x"C0C0C0F9F8909082",
 17997 => x"C0C0C0F9F89090F8",
 17998 => x"C0C0C0F9F8909080",
 17999 => x"C0C0C0F9F8909090",
 18000 => x"C0C0C0F980C0C0C0",
 18001 => x"C0C0C0F980C0C0F9",
 18002 => x"C0C0C0F980C0C0A4",
 18003 => x"C0C0C0F980C0C0B0",
 18004 => x"C0C0C0F980C0C099",
 18005 => x"C0C0C0F980C0C092",
 18006 => x"C0C0C0F980C0C082",
 18007 => x"C0C0C0F980C0C0F8",
 18008 => x"C0C0C0F980C0C080",
 18009 => x"C0C0C0F980C0C090",
 18010 => x"C0C0C0F980C0F9C0",
 18011 => x"C0C0C0F980C0F9F9",
 18012 => x"C0C0C0F980C0F9A4",
 18013 => x"C0C0C0F980C0F9B0",
 18014 => x"C0C0C0F980C0F999",
 18015 => x"C0C0C0F980C0F992",
 18016 => x"C0C0C0F980C0F982",
 18017 => x"C0C0C0F980C0F9F8",
 18018 => x"C0C0C0F980C0F980",
 18019 => x"C0C0C0F980C0F990",
 18020 => x"C0C0C0F980C0A4C0",
 18021 => x"C0C0C0F980C0A4F9",
 18022 => x"C0C0C0F980C0A4A4",
 18023 => x"C0C0C0F980C0A4B0",
 18024 => x"C0C0C0F980C0A499",
 18025 => x"C0C0C0F980C0A492",
 18026 => x"C0C0C0F980C0A482",
 18027 => x"C0C0C0F980C0A4F8",
 18028 => x"C0C0C0F980C0A480",
 18029 => x"C0C0C0F980C0A490",
 18030 => x"C0C0C0F980C0B0C0",
 18031 => x"C0C0C0F980C0B0F9",
 18032 => x"C0C0C0F980C0B0A4",
 18033 => x"C0C0C0F980C0B0B0",
 18034 => x"C0C0C0F980C0B099",
 18035 => x"C0C0C0F980C0B092",
 18036 => x"C0C0C0F980C0B082",
 18037 => x"C0C0C0F980C0B0F8",
 18038 => x"C0C0C0F980C0B080",
 18039 => x"C0C0C0F980C0B090",
 18040 => x"C0C0C0F980C099C0",
 18041 => x"C0C0C0F980C099F9",
 18042 => x"C0C0C0F980C099A4",
 18043 => x"C0C0C0F980C099B0",
 18044 => x"C0C0C0F980C09999",
 18045 => x"C0C0C0F980C09992",
 18046 => x"C0C0C0F980C09982",
 18047 => x"C0C0C0F980C099F8",
 18048 => x"C0C0C0F980C09980",
 18049 => x"C0C0C0F980C09990",
 18050 => x"C0C0C0F980C092C0",
 18051 => x"C0C0C0F980C092F9",
 18052 => x"C0C0C0F980C092A4",
 18053 => x"C0C0C0F980C092B0",
 18054 => x"C0C0C0F980C09299",
 18055 => x"C0C0C0F980C09292",
 18056 => x"C0C0C0F980C09282",
 18057 => x"C0C0C0F980C092F8",
 18058 => x"C0C0C0F980C09280",
 18059 => x"C0C0C0F980C09290",
 18060 => x"C0C0C0F980C082C0",
 18061 => x"C0C0C0F980C082F9",
 18062 => x"C0C0C0F980C082A4",
 18063 => x"C0C0C0F980C082B0",
 18064 => x"C0C0C0F980C08299",
 18065 => x"C0C0C0F980C08292",
 18066 => x"C0C0C0F980C08282",
 18067 => x"C0C0C0F980C082F8",
 18068 => x"C0C0C0F980C08280",
 18069 => x"C0C0C0F980C08290",
 18070 => x"C0C0C0F980C0F8C0",
 18071 => x"C0C0C0F980C0F8F9",
 18072 => x"C0C0C0F980C0F8A4",
 18073 => x"C0C0C0F980C0F8B0",
 18074 => x"C0C0C0F980C0F899",
 18075 => x"C0C0C0F980C0F892",
 18076 => x"C0C0C0F980C0F882",
 18077 => x"C0C0C0F980C0F8F8",
 18078 => x"C0C0C0F980C0F880",
 18079 => x"C0C0C0F980C0F890",
 18080 => x"C0C0C0F980C080C0",
 18081 => x"C0C0C0F980C080F9",
 18082 => x"C0C0C0F980C080A4",
 18083 => x"C0C0C0F980C080B0",
 18084 => x"C0C0C0F980C08099",
 18085 => x"C0C0C0F980C08092",
 18086 => x"C0C0C0F980C08082",
 18087 => x"C0C0C0F980C080F8",
 18088 => x"C0C0C0F980C08080",
 18089 => x"C0C0C0F980C08090",
 18090 => x"C0C0C0F980C090C0",
 18091 => x"C0C0C0F980C090F9",
 18092 => x"C0C0C0F980C090A4",
 18093 => x"C0C0C0F980C090B0",
 18094 => x"C0C0C0F980C09099",
 18095 => x"C0C0C0F980C09092",
 18096 => x"C0C0C0F980C09082",
 18097 => x"C0C0C0F980C090F8",
 18098 => x"C0C0C0F980C09080",
 18099 => x"C0C0C0F980C09090",
 18100 => x"C0C0C0F980F9C0C0",
 18101 => x"C0C0C0F980F9C0F9",
 18102 => x"C0C0C0F980F9C0A4",
 18103 => x"C0C0C0F980F9C0B0",
 18104 => x"C0C0C0F980F9C099",
 18105 => x"C0C0C0F980F9C092",
 18106 => x"C0C0C0F980F9C082",
 18107 => x"C0C0C0F980F9C0F8",
 18108 => x"C0C0C0F980F9C080",
 18109 => x"C0C0C0F980F9C090",
 18110 => x"C0C0C0F980F9F9C0",
 18111 => x"C0C0C0F980F9F9F9",
 18112 => x"C0C0C0F980F9F9A4",
 18113 => x"C0C0C0F980F9F9B0",
 18114 => x"C0C0C0F980F9F999",
 18115 => x"C0C0C0F980F9F992",
 18116 => x"C0C0C0F980F9F982",
 18117 => x"C0C0C0F980F9F9F8",
 18118 => x"C0C0C0F980F9F980",
 18119 => x"C0C0C0F980F9F990",
 18120 => x"C0C0C0F980F9A4C0",
 18121 => x"C0C0C0F980F9A4F9",
 18122 => x"C0C0C0F980F9A4A4",
 18123 => x"C0C0C0F980F9A4B0",
 18124 => x"C0C0C0F980F9A499",
 18125 => x"C0C0C0F980F9A492",
 18126 => x"C0C0C0F980F9A482",
 18127 => x"C0C0C0F980F9A4F8",
 18128 => x"C0C0C0F980F9A480",
 18129 => x"C0C0C0F980F9A490",
 18130 => x"C0C0C0F980F9B0C0",
 18131 => x"C0C0C0F980F9B0F9",
 18132 => x"C0C0C0F980F9B0A4",
 18133 => x"C0C0C0F980F9B0B0",
 18134 => x"C0C0C0F980F9B099",
 18135 => x"C0C0C0F980F9B092",
 18136 => x"C0C0C0F980F9B082",
 18137 => x"C0C0C0F980F9B0F8",
 18138 => x"C0C0C0F980F9B080",
 18139 => x"C0C0C0F980F9B090",
 18140 => x"C0C0C0F980F999C0",
 18141 => x"C0C0C0F980F999F9",
 18142 => x"C0C0C0F980F999A4",
 18143 => x"C0C0C0F980F999B0",
 18144 => x"C0C0C0F980F99999",
 18145 => x"C0C0C0F980F99992",
 18146 => x"C0C0C0F980F99982",
 18147 => x"C0C0C0F980F999F8",
 18148 => x"C0C0C0F980F99980",
 18149 => x"C0C0C0F980F99990",
 18150 => x"C0C0C0F980F992C0",
 18151 => x"C0C0C0F980F992F9",
 18152 => x"C0C0C0F980F992A4",
 18153 => x"C0C0C0F980F992B0",
 18154 => x"C0C0C0F980F99299",
 18155 => x"C0C0C0F980F99292",
 18156 => x"C0C0C0F980F99282",
 18157 => x"C0C0C0F980F992F8",
 18158 => x"C0C0C0F980F99280",
 18159 => x"C0C0C0F980F99290",
 18160 => x"C0C0C0F980F982C0",
 18161 => x"C0C0C0F980F982F9",
 18162 => x"C0C0C0F980F982A4",
 18163 => x"C0C0C0F980F982B0",
 18164 => x"C0C0C0F980F98299",
 18165 => x"C0C0C0F980F98292",
 18166 => x"C0C0C0F980F98282",
 18167 => x"C0C0C0F980F982F8",
 18168 => x"C0C0C0F980F98280",
 18169 => x"C0C0C0F980F98290",
 18170 => x"C0C0C0F980F9F8C0",
 18171 => x"C0C0C0F980F9F8F9",
 18172 => x"C0C0C0F980F9F8A4",
 18173 => x"C0C0C0F980F9F8B0",
 18174 => x"C0C0C0F980F9F899",
 18175 => x"C0C0C0F980F9F892",
 18176 => x"C0C0C0F980F9F882",
 18177 => x"C0C0C0F980F9F8F8",
 18178 => x"C0C0C0F980F9F880",
 18179 => x"C0C0C0F980F9F890",
 18180 => x"C0C0C0F980F980C0",
 18181 => x"C0C0C0F980F980F9",
 18182 => x"C0C0C0F980F980A4",
 18183 => x"C0C0C0F980F980B0",
 18184 => x"C0C0C0F980F98099",
 18185 => x"C0C0C0F980F98092",
 18186 => x"C0C0C0F980F98082",
 18187 => x"C0C0C0F980F980F8",
 18188 => x"C0C0C0F980F98080",
 18189 => x"C0C0C0F980F98090",
 18190 => x"C0C0C0F980F990C0",
 18191 => x"C0C0C0F980F990F9",
 18192 => x"C0C0C0F980F990A4",
 18193 => x"C0C0C0F980F990B0",
 18194 => x"C0C0C0F980F99099",
 18195 => x"C0C0C0F980F99092",
 18196 => x"C0C0C0F980F99082",
 18197 => x"C0C0C0F980F990F8",
 18198 => x"C0C0C0F980F99080",
 18199 => x"C0C0C0F980F99090",
 18200 => x"C0C0C0F980A4C0C0",
 18201 => x"C0C0C0F980A4C0F9",
 18202 => x"C0C0C0F980A4C0A4",
 18203 => x"C0C0C0F980A4C0B0",
 18204 => x"C0C0C0F980A4C099",
 18205 => x"C0C0C0F980A4C092",
 18206 => x"C0C0C0F980A4C082",
 18207 => x"C0C0C0F980A4C0F8",
 18208 => x"C0C0C0F980A4C080",
 18209 => x"C0C0C0F980A4C090",
 18210 => x"C0C0C0F980A4F9C0",
 18211 => x"C0C0C0F980A4F9F9",
 18212 => x"C0C0C0F980A4F9A4",
 18213 => x"C0C0C0F980A4F9B0",
 18214 => x"C0C0C0F980A4F999",
 18215 => x"C0C0C0F980A4F992",
 18216 => x"C0C0C0F980A4F982",
 18217 => x"C0C0C0F980A4F9F8",
 18218 => x"C0C0C0F980A4F980",
 18219 => x"C0C0C0F980A4F990",
 18220 => x"C0C0C0F980A4A4C0",
 18221 => x"C0C0C0F980A4A4F9",
 18222 => x"C0C0C0F980A4A4A4",
 18223 => x"C0C0C0F980A4A4B0",
 18224 => x"C0C0C0F980A4A499",
 18225 => x"C0C0C0F980A4A492",
 18226 => x"C0C0C0F980A4A482",
 18227 => x"C0C0C0F980A4A4F8",
 18228 => x"C0C0C0F980A4A480",
 18229 => x"C0C0C0F980A4A490",
 18230 => x"C0C0C0F980A4B0C0",
 18231 => x"C0C0C0F980A4B0F9",
 18232 => x"C0C0C0F980A4B0A4",
 18233 => x"C0C0C0F980A4B0B0",
 18234 => x"C0C0C0F980A4B099",
 18235 => x"C0C0C0F980A4B092",
 18236 => x"C0C0C0F980A4B082",
 18237 => x"C0C0C0F980A4B0F8",
 18238 => x"C0C0C0F980A4B080",
 18239 => x"C0C0C0F980A4B090",
 18240 => x"C0C0C0F980A499C0",
 18241 => x"C0C0C0F980A499F9",
 18242 => x"C0C0C0F980A499A4",
 18243 => x"C0C0C0F980A499B0",
 18244 => x"C0C0C0F980A49999",
 18245 => x"C0C0C0F980A49992",
 18246 => x"C0C0C0F980A49982",
 18247 => x"C0C0C0F980A499F8",
 18248 => x"C0C0C0F980A49980",
 18249 => x"C0C0C0F980A49990",
 18250 => x"C0C0C0F980A492C0",
 18251 => x"C0C0C0F980A492F9",
 18252 => x"C0C0C0F980A492A4",
 18253 => x"C0C0C0F980A492B0",
 18254 => x"C0C0C0F980A49299",
 18255 => x"C0C0C0F980A49292",
 18256 => x"C0C0C0F980A49282",
 18257 => x"C0C0C0F980A492F8",
 18258 => x"C0C0C0F980A49280",
 18259 => x"C0C0C0F980A49290",
 18260 => x"C0C0C0F980A482C0",
 18261 => x"C0C0C0F980A482F9",
 18262 => x"C0C0C0F980A482A4",
 18263 => x"C0C0C0F980A482B0",
 18264 => x"C0C0C0F980A48299",
 18265 => x"C0C0C0F980A48292",
 18266 => x"C0C0C0F980A48282",
 18267 => x"C0C0C0F980A482F8",
 18268 => x"C0C0C0F980A48280",
 18269 => x"C0C0C0F980A48290",
 18270 => x"C0C0C0F980A4F8C0",
 18271 => x"C0C0C0F980A4F8F9",
 18272 => x"C0C0C0F980A4F8A4",
 18273 => x"C0C0C0F980A4F8B0",
 18274 => x"C0C0C0F980A4F899",
 18275 => x"C0C0C0F980A4F892",
 18276 => x"C0C0C0F980A4F882",
 18277 => x"C0C0C0F980A4F8F8",
 18278 => x"C0C0C0F980A4F880",
 18279 => x"C0C0C0F980A4F890",
 18280 => x"C0C0C0F980A480C0",
 18281 => x"C0C0C0F980A480F9",
 18282 => x"C0C0C0F980A480A4",
 18283 => x"C0C0C0F980A480B0",
 18284 => x"C0C0C0F980A48099",
 18285 => x"C0C0C0F980A48092",
 18286 => x"C0C0C0F980A48082",
 18287 => x"C0C0C0F980A480F8",
 18288 => x"C0C0C0F980A48080",
 18289 => x"C0C0C0F980A48090",
 18290 => x"C0C0C0F980A490C0",
 18291 => x"C0C0C0F980A490F9",
 18292 => x"C0C0C0F980A490A4",
 18293 => x"C0C0C0F980A490B0",
 18294 => x"C0C0C0F980A49099",
 18295 => x"C0C0C0F980A49092",
 18296 => x"C0C0C0F980A49082",
 18297 => x"C0C0C0F980A490F8",
 18298 => x"C0C0C0F980A49080",
 18299 => x"C0C0C0F980A49090",
 18300 => x"C0C0C0F980B0C0C0",
 18301 => x"C0C0C0F980B0C0F9",
 18302 => x"C0C0C0F980B0C0A4",
 18303 => x"C0C0C0F980B0C0B0",
 18304 => x"C0C0C0F980B0C099",
 18305 => x"C0C0C0F980B0C092",
 18306 => x"C0C0C0F980B0C082",
 18307 => x"C0C0C0F980B0C0F8",
 18308 => x"C0C0C0F980B0C080",
 18309 => x"C0C0C0F980B0C090",
 18310 => x"C0C0C0F980B0F9C0",
 18311 => x"C0C0C0F980B0F9F9",
 18312 => x"C0C0C0F980B0F9A4",
 18313 => x"C0C0C0F980B0F9B0",
 18314 => x"C0C0C0F980B0F999",
 18315 => x"C0C0C0F980B0F992",
 18316 => x"C0C0C0F980B0F982",
 18317 => x"C0C0C0F980B0F9F8",
 18318 => x"C0C0C0F980B0F980",
 18319 => x"C0C0C0F980B0F990",
 18320 => x"C0C0C0F980B0A4C0",
 18321 => x"C0C0C0F980B0A4F9",
 18322 => x"C0C0C0F980B0A4A4",
 18323 => x"C0C0C0F980B0A4B0",
 18324 => x"C0C0C0F980B0A499",
 18325 => x"C0C0C0F980B0A492",
 18326 => x"C0C0C0F980B0A482",
 18327 => x"C0C0C0F980B0A4F8",
 18328 => x"C0C0C0F980B0A480",
 18329 => x"C0C0C0F980B0A490",
 18330 => x"C0C0C0F980B0B0C0",
 18331 => x"C0C0C0F980B0B0F9",
 18332 => x"C0C0C0F980B0B0A4",
 18333 => x"C0C0C0F980B0B0B0",
 18334 => x"C0C0C0F980B0B099",
 18335 => x"C0C0C0F980B0B092",
 18336 => x"C0C0C0F980B0B082",
 18337 => x"C0C0C0F980B0B0F8",
 18338 => x"C0C0C0F980B0B080",
 18339 => x"C0C0C0F980B0B090",
 18340 => x"C0C0C0F980B099C0",
 18341 => x"C0C0C0F980B099F9",
 18342 => x"C0C0C0F980B099A4",
 18343 => x"C0C0C0F980B099B0",
 18344 => x"C0C0C0F980B09999",
 18345 => x"C0C0C0F980B09992",
 18346 => x"C0C0C0F980B09982",
 18347 => x"C0C0C0F980B099F8",
 18348 => x"C0C0C0F980B09980",
 18349 => x"C0C0C0F980B09990",
 18350 => x"C0C0C0F980B092C0",
 18351 => x"C0C0C0F980B092F9",
 18352 => x"C0C0C0F980B092A4",
 18353 => x"C0C0C0F980B092B0",
 18354 => x"C0C0C0F980B09299",
 18355 => x"C0C0C0F980B09292",
 18356 => x"C0C0C0F980B09282",
 18357 => x"C0C0C0F980B092F8",
 18358 => x"C0C0C0F980B09280",
 18359 => x"C0C0C0F980B09290",
 18360 => x"C0C0C0F980B082C0",
 18361 => x"C0C0C0F980B082F9",
 18362 => x"C0C0C0F980B082A4",
 18363 => x"C0C0C0F980B082B0",
 18364 => x"C0C0C0F980B08299",
 18365 => x"C0C0C0F980B08292",
 18366 => x"C0C0C0F980B08282",
 18367 => x"C0C0C0F980B082F8",
 18368 => x"C0C0C0F980B08280",
 18369 => x"C0C0C0F980B08290",
 18370 => x"C0C0C0F980B0F8C0",
 18371 => x"C0C0C0F980B0F8F9",
 18372 => x"C0C0C0F980B0F8A4",
 18373 => x"C0C0C0F980B0F8B0",
 18374 => x"C0C0C0F980B0F899",
 18375 => x"C0C0C0F980B0F892",
 18376 => x"C0C0C0F980B0F882",
 18377 => x"C0C0C0F980B0F8F8",
 18378 => x"C0C0C0F980B0F880",
 18379 => x"C0C0C0F980B0F890",
 18380 => x"C0C0C0F980B080C0",
 18381 => x"C0C0C0F980B080F9",
 18382 => x"C0C0C0F980B080A4",
 18383 => x"C0C0C0F980B080B0",
 18384 => x"C0C0C0F980B08099",
 18385 => x"C0C0C0F980B08092",
 18386 => x"C0C0C0F980B08082",
 18387 => x"C0C0C0F980B080F8",
 18388 => x"C0C0C0F980B08080",
 18389 => x"C0C0C0F980B08090",
 18390 => x"C0C0C0F980B090C0",
 18391 => x"C0C0C0F980B090F9",
 18392 => x"C0C0C0F980B090A4",
 18393 => x"C0C0C0F980B090B0",
 18394 => x"C0C0C0F980B09099",
 18395 => x"C0C0C0F980B09092",
 18396 => x"C0C0C0F980B09082",
 18397 => x"C0C0C0F980B090F8",
 18398 => x"C0C0C0F980B09080",
 18399 => x"C0C0C0F980B09090",
 18400 => x"C0C0C0F98099C0C0",
 18401 => x"C0C0C0F98099C0F9",
 18402 => x"C0C0C0F98099C0A4",
 18403 => x"C0C0C0F98099C0B0",
 18404 => x"C0C0C0F98099C099",
 18405 => x"C0C0C0F98099C092",
 18406 => x"C0C0C0F98099C082",
 18407 => x"C0C0C0F98099C0F8",
 18408 => x"C0C0C0F98099C080",
 18409 => x"C0C0C0F98099C090",
 18410 => x"C0C0C0F98099F9C0",
 18411 => x"C0C0C0F98099F9F9",
 18412 => x"C0C0C0F98099F9A4",
 18413 => x"C0C0C0F98099F9B0",
 18414 => x"C0C0C0F98099F999",
 18415 => x"C0C0C0F98099F992",
 18416 => x"C0C0C0F98099F982",
 18417 => x"C0C0C0F98099F9F8",
 18418 => x"C0C0C0F98099F980",
 18419 => x"C0C0C0F98099F990",
 18420 => x"C0C0C0F98099A4C0",
 18421 => x"C0C0C0F98099A4F9",
 18422 => x"C0C0C0F98099A4A4",
 18423 => x"C0C0C0F98099A4B0",
 18424 => x"C0C0C0F98099A499",
 18425 => x"C0C0C0F98099A492",
 18426 => x"C0C0C0F98099A482",
 18427 => x"C0C0C0F98099A4F8",
 18428 => x"C0C0C0F98099A480",
 18429 => x"C0C0C0F98099A490",
 18430 => x"C0C0C0F98099B0C0",
 18431 => x"C0C0C0F98099B0F9",
 18432 => x"C0C0C0F98099B0A4",
 18433 => x"C0C0C0F98099B0B0",
 18434 => x"C0C0C0F98099B099",
 18435 => x"C0C0C0F98099B092",
 18436 => x"C0C0C0F98099B082",
 18437 => x"C0C0C0F98099B0F8",
 18438 => x"C0C0C0F98099B080",
 18439 => x"C0C0C0F98099B090",
 18440 => x"C0C0C0F9809999C0",
 18441 => x"C0C0C0F9809999F9",
 18442 => x"C0C0C0F9809999A4",
 18443 => x"C0C0C0F9809999B0",
 18444 => x"C0C0C0F980999999",
 18445 => x"C0C0C0F980999992",
 18446 => x"C0C0C0F980999982",
 18447 => x"C0C0C0F9809999F8",
 18448 => x"C0C0C0F980999980",
 18449 => x"C0C0C0F980999990",
 18450 => x"C0C0C0F9809992C0",
 18451 => x"C0C0C0F9809992F9",
 18452 => x"C0C0C0F9809992A4",
 18453 => x"C0C0C0F9809992B0",
 18454 => x"C0C0C0F980999299",
 18455 => x"C0C0C0F980999292",
 18456 => x"C0C0C0F980999282",
 18457 => x"C0C0C0F9809992F8",
 18458 => x"C0C0C0F980999280",
 18459 => x"C0C0C0F980999290",
 18460 => x"C0C0C0F9809982C0",
 18461 => x"C0C0C0F9809982F9",
 18462 => x"C0C0C0F9809982A4",
 18463 => x"C0C0C0F9809982B0",
 18464 => x"C0C0C0F980998299",
 18465 => x"C0C0C0F980998292",
 18466 => x"C0C0C0F980998282",
 18467 => x"C0C0C0F9809982F8",
 18468 => x"C0C0C0F980998280",
 18469 => x"C0C0C0F980998290",
 18470 => x"C0C0C0F98099F8C0",
 18471 => x"C0C0C0F98099F8F9",
 18472 => x"C0C0C0F98099F8A4",
 18473 => x"C0C0C0F98099F8B0",
 18474 => x"C0C0C0F98099F899",
 18475 => x"C0C0C0F98099F892",
 18476 => x"C0C0C0F98099F882",
 18477 => x"C0C0C0F98099F8F8",
 18478 => x"C0C0C0F98099F880",
 18479 => x"C0C0C0F98099F890",
 18480 => x"C0C0C0F9809980C0",
 18481 => x"C0C0C0F9809980F9",
 18482 => x"C0C0C0F9809980A4",
 18483 => x"C0C0C0F9809980B0",
 18484 => x"C0C0C0F980998099",
 18485 => x"C0C0C0F980998092",
 18486 => x"C0C0C0F980998082",
 18487 => x"C0C0C0F9809980F8",
 18488 => x"C0C0C0F980998080",
 18489 => x"C0C0C0F980998090",
 18490 => x"C0C0C0F9809990C0",
 18491 => x"C0C0C0F9809990F9",
 18492 => x"C0C0C0F9809990A4",
 18493 => x"C0C0C0F9809990B0",
 18494 => x"C0C0C0F980999099",
 18495 => x"C0C0C0F980999092",
 18496 => x"C0C0C0F980999082",
 18497 => x"C0C0C0F9809990F8",
 18498 => x"C0C0C0F980999080",
 18499 => x"C0C0C0F980999090",
 18500 => x"C0C0C0F98092C0C0",
 18501 => x"C0C0C0F98092C0F9",
 18502 => x"C0C0C0F98092C0A4",
 18503 => x"C0C0C0F98092C0B0",
 18504 => x"C0C0C0F98092C099",
 18505 => x"C0C0C0F98092C092",
 18506 => x"C0C0C0F98092C082",
 18507 => x"C0C0C0F98092C0F8",
 18508 => x"C0C0C0F98092C080",
 18509 => x"C0C0C0F98092C090",
 18510 => x"C0C0C0F98092F9C0",
 18511 => x"C0C0C0F98092F9F9",
 18512 => x"C0C0C0F98092F9A4",
 18513 => x"C0C0C0F98092F9B0",
 18514 => x"C0C0C0F98092F999",
 18515 => x"C0C0C0F98092F992",
 18516 => x"C0C0C0F98092F982",
 18517 => x"C0C0C0F98092F9F8",
 18518 => x"C0C0C0F98092F980",
 18519 => x"C0C0C0F98092F990",
 18520 => x"C0C0C0F98092A4C0",
 18521 => x"C0C0C0F98092A4F9",
 18522 => x"C0C0C0F98092A4A4",
 18523 => x"C0C0C0F98092A4B0",
 18524 => x"C0C0C0F98092A499",
 18525 => x"C0C0C0F98092A492",
 18526 => x"C0C0C0F98092A482",
 18527 => x"C0C0C0F98092A4F8",
 18528 => x"C0C0C0F98092A480",
 18529 => x"C0C0C0F98092A490",
 18530 => x"C0C0C0F98092B0C0",
 18531 => x"C0C0C0F98092B0F9",
 18532 => x"C0C0C0F98092B0A4",
 18533 => x"C0C0C0F98092B0B0",
 18534 => x"C0C0C0F98092B099",
 18535 => x"C0C0C0F98092B092",
 18536 => x"C0C0C0F98092B082",
 18537 => x"C0C0C0F98092B0F8",
 18538 => x"C0C0C0F98092B080",
 18539 => x"C0C0C0F98092B090",
 18540 => x"C0C0C0F9809299C0",
 18541 => x"C0C0C0F9809299F9",
 18542 => x"C0C0C0F9809299A4",
 18543 => x"C0C0C0F9809299B0",
 18544 => x"C0C0C0F980929999",
 18545 => x"C0C0C0F980929992",
 18546 => x"C0C0C0F980929982",
 18547 => x"C0C0C0F9809299F8",
 18548 => x"C0C0C0F980929980",
 18549 => x"C0C0C0F980929990",
 18550 => x"C0C0C0F9809292C0",
 18551 => x"C0C0C0F9809292F9",
 18552 => x"C0C0C0F9809292A4",
 18553 => x"C0C0C0F9809292B0",
 18554 => x"C0C0C0F980929299",
 18555 => x"C0C0C0F980929292",
 18556 => x"C0C0C0F980929282",
 18557 => x"C0C0C0F9809292F8",
 18558 => x"C0C0C0F980929280",
 18559 => x"C0C0C0F980929290",
 18560 => x"C0C0C0F9809282C0",
 18561 => x"C0C0C0F9809282F9",
 18562 => x"C0C0C0F9809282A4",
 18563 => x"C0C0C0F9809282B0",
 18564 => x"C0C0C0F980928299",
 18565 => x"C0C0C0F980928292",
 18566 => x"C0C0C0F980928282",
 18567 => x"C0C0C0F9809282F8",
 18568 => x"C0C0C0F980928280",
 18569 => x"C0C0C0F980928290",
 18570 => x"C0C0C0F98092F8C0",
 18571 => x"C0C0C0F98092F8F9",
 18572 => x"C0C0C0F98092F8A4",
 18573 => x"C0C0C0F98092F8B0",
 18574 => x"C0C0C0F98092F899",
 18575 => x"C0C0C0F98092F892",
 18576 => x"C0C0C0F98092F882",
 18577 => x"C0C0C0F98092F8F8",
 18578 => x"C0C0C0F98092F880",
 18579 => x"C0C0C0F98092F890",
 18580 => x"C0C0C0F9809280C0",
 18581 => x"C0C0C0F9809280F9",
 18582 => x"C0C0C0F9809280A4",
 18583 => x"C0C0C0F9809280B0",
 18584 => x"C0C0C0F980928099",
 18585 => x"C0C0C0F980928092",
 18586 => x"C0C0C0F980928082",
 18587 => x"C0C0C0F9809280F8",
 18588 => x"C0C0C0F980928080",
 18589 => x"C0C0C0F980928090",
 18590 => x"C0C0C0F9809290C0",
 18591 => x"C0C0C0F9809290F9",
 18592 => x"C0C0C0F9809290A4",
 18593 => x"C0C0C0F9809290B0",
 18594 => x"C0C0C0F980929099",
 18595 => x"C0C0C0F980929092",
 18596 => x"C0C0C0F980929082",
 18597 => x"C0C0C0F9809290F8",
 18598 => x"C0C0C0F980929080",
 18599 => x"C0C0C0F980929090",
 18600 => x"C0C0C0F98082C0C0",
 18601 => x"C0C0C0F98082C0F9",
 18602 => x"C0C0C0F98082C0A4",
 18603 => x"C0C0C0F98082C0B0",
 18604 => x"C0C0C0F98082C099",
 18605 => x"C0C0C0F98082C092",
 18606 => x"C0C0C0F98082C082",
 18607 => x"C0C0C0F98082C0F8",
 18608 => x"C0C0C0F98082C080",
 18609 => x"C0C0C0F98082C090",
 18610 => x"C0C0C0F98082F9C0",
 18611 => x"C0C0C0F98082F9F9",
 18612 => x"C0C0C0F98082F9A4",
 18613 => x"C0C0C0F98082F9B0",
 18614 => x"C0C0C0F98082F999",
 18615 => x"C0C0C0F98082F992",
 18616 => x"C0C0C0F98082F982",
 18617 => x"C0C0C0F98082F9F8",
 18618 => x"C0C0C0F98082F980",
 18619 => x"C0C0C0F98082F990",
 18620 => x"C0C0C0F98082A4C0",
 18621 => x"C0C0C0F98082A4F9",
 18622 => x"C0C0C0F98082A4A4",
 18623 => x"C0C0C0F98082A4B0",
 18624 => x"C0C0C0F98082A499",
 18625 => x"C0C0C0F98082A492",
 18626 => x"C0C0C0F98082A482",
 18627 => x"C0C0C0F98082A4F8",
 18628 => x"C0C0C0F98082A480",
 18629 => x"C0C0C0F98082A490",
 18630 => x"C0C0C0F98082B0C0",
 18631 => x"C0C0C0F98082B0F9",
 18632 => x"C0C0C0F98082B0A4",
 18633 => x"C0C0C0F98082B0B0",
 18634 => x"C0C0C0F98082B099",
 18635 => x"C0C0C0F98082B092",
 18636 => x"C0C0C0F98082B082",
 18637 => x"C0C0C0F98082B0F8",
 18638 => x"C0C0C0F98082B080",
 18639 => x"C0C0C0F98082B090",
 18640 => x"C0C0C0F9808299C0",
 18641 => x"C0C0C0F9808299F9",
 18642 => x"C0C0C0F9808299A4",
 18643 => x"C0C0C0F9808299B0",
 18644 => x"C0C0C0F980829999",
 18645 => x"C0C0C0F980829992",
 18646 => x"C0C0C0F980829982",
 18647 => x"C0C0C0F9808299F8",
 18648 => x"C0C0C0F980829980",
 18649 => x"C0C0C0F980829990",
 18650 => x"C0C0C0F9808292C0",
 18651 => x"C0C0C0F9808292F9",
 18652 => x"C0C0C0F9808292A4",
 18653 => x"C0C0C0F9808292B0",
 18654 => x"C0C0C0F980829299",
 18655 => x"C0C0C0F980829292",
 18656 => x"C0C0C0F980829282",
 18657 => x"C0C0C0F9808292F8",
 18658 => x"C0C0C0F980829280",
 18659 => x"C0C0C0F980829290",
 18660 => x"C0C0C0F9808282C0",
 18661 => x"C0C0C0F9808282F9",
 18662 => x"C0C0C0F9808282A4",
 18663 => x"C0C0C0F9808282B0",
 18664 => x"C0C0C0F980828299",
 18665 => x"C0C0C0F980828292",
 18666 => x"C0C0C0F980828282",
 18667 => x"C0C0C0F9808282F8",
 18668 => x"C0C0C0F980828280",
 18669 => x"C0C0C0F980828290",
 18670 => x"C0C0C0F98082F8C0",
 18671 => x"C0C0C0F98082F8F9",
 18672 => x"C0C0C0F98082F8A4",
 18673 => x"C0C0C0F98082F8B0",
 18674 => x"C0C0C0F98082F899",
 18675 => x"C0C0C0F98082F892",
 18676 => x"C0C0C0F98082F882",
 18677 => x"C0C0C0F98082F8F8",
 18678 => x"C0C0C0F98082F880",
 18679 => x"C0C0C0F98082F890",
 18680 => x"C0C0C0F9808280C0",
 18681 => x"C0C0C0F9808280F9",
 18682 => x"C0C0C0F9808280A4",
 18683 => x"C0C0C0F9808280B0",
 18684 => x"C0C0C0F980828099",
 18685 => x"C0C0C0F980828092",
 18686 => x"C0C0C0F980828082",
 18687 => x"C0C0C0F9808280F8",
 18688 => x"C0C0C0F980828080",
 18689 => x"C0C0C0F980828090",
 18690 => x"C0C0C0F9808290C0",
 18691 => x"C0C0C0F9808290F9",
 18692 => x"C0C0C0F9808290A4",
 18693 => x"C0C0C0F9808290B0",
 18694 => x"C0C0C0F980829099",
 18695 => x"C0C0C0F980829092",
 18696 => x"C0C0C0F980829082",
 18697 => x"C0C0C0F9808290F8",
 18698 => x"C0C0C0F980829080",
 18699 => x"C0C0C0F980829090",
 18700 => x"C0C0C0F980F8C0C0",
 18701 => x"C0C0C0F980F8C0F9",
 18702 => x"C0C0C0F980F8C0A4",
 18703 => x"C0C0C0F980F8C0B0",
 18704 => x"C0C0C0F980F8C099",
 18705 => x"C0C0C0F980F8C092",
 18706 => x"C0C0C0F980F8C082",
 18707 => x"C0C0C0F980F8C0F8",
 18708 => x"C0C0C0F980F8C080",
 18709 => x"C0C0C0F980F8C090",
 18710 => x"C0C0C0F980F8F9C0",
 18711 => x"C0C0C0F980F8F9F9",
 18712 => x"C0C0C0F980F8F9A4",
 18713 => x"C0C0C0F980F8F9B0",
 18714 => x"C0C0C0F980F8F999",
 18715 => x"C0C0C0F980F8F992",
 18716 => x"C0C0C0F980F8F982",
 18717 => x"C0C0C0F980F8F9F8",
 18718 => x"C0C0C0F980F8F980",
 18719 => x"C0C0C0F980F8F990",
 18720 => x"C0C0C0F980F8A4C0",
 18721 => x"C0C0C0F980F8A4F9",
 18722 => x"C0C0C0F980F8A4A4",
 18723 => x"C0C0C0F980F8A4B0",
 18724 => x"C0C0C0F980F8A499",
 18725 => x"C0C0C0F980F8A492",
 18726 => x"C0C0C0F980F8A482",
 18727 => x"C0C0C0F980F8A4F8",
 18728 => x"C0C0C0F980F8A480",
 18729 => x"C0C0C0F980F8A490",
 18730 => x"C0C0C0F980F8B0C0",
 18731 => x"C0C0C0F980F8B0F9",
 18732 => x"C0C0C0F980F8B0A4",
 18733 => x"C0C0C0F980F8B0B0",
 18734 => x"C0C0C0F980F8B099",
 18735 => x"C0C0C0F980F8B092",
 18736 => x"C0C0C0F980F8B082",
 18737 => x"C0C0C0F980F8B0F8",
 18738 => x"C0C0C0F980F8B080",
 18739 => x"C0C0C0F980F8B090",
 18740 => x"C0C0C0F980F899C0",
 18741 => x"C0C0C0F980F899F9",
 18742 => x"C0C0C0F980F899A4",
 18743 => x"C0C0C0F980F899B0",
 18744 => x"C0C0C0F980F89999",
 18745 => x"C0C0C0F980F89992",
 18746 => x"C0C0C0F980F89982",
 18747 => x"C0C0C0F980F899F8",
 18748 => x"C0C0C0F980F89980",
 18749 => x"C0C0C0F980F89990",
 18750 => x"C0C0C0F980F892C0",
 18751 => x"C0C0C0F980F892F9",
 18752 => x"C0C0C0F980F892A4",
 18753 => x"C0C0C0F980F892B0",
 18754 => x"C0C0C0F980F89299",
 18755 => x"C0C0C0F980F89292",
 18756 => x"C0C0C0F980F89282",
 18757 => x"C0C0C0F980F892F8",
 18758 => x"C0C0C0F980F89280",
 18759 => x"C0C0C0F980F89290",
 18760 => x"C0C0C0F980F882C0",
 18761 => x"C0C0C0F980F882F9",
 18762 => x"C0C0C0F980F882A4",
 18763 => x"C0C0C0F980F882B0",
 18764 => x"C0C0C0F980F88299",
 18765 => x"C0C0C0F980F88292",
 18766 => x"C0C0C0F980F88282",
 18767 => x"C0C0C0F980F882F8",
 18768 => x"C0C0C0F980F88280",
 18769 => x"C0C0C0F980F88290",
 18770 => x"C0C0C0F980F8F8C0",
 18771 => x"C0C0C0F980F8F8F9",
 18772 => x"C0C0C0F980F8F8A4",
 18773 => x"C0C0C0F980F8F8B0",
 18774 => x"C0C0C0F980F8F899",
 18775 => x"C0C0C0F980F8F892",
 18776 => x"C0C0C0F980F8F882",
 18777 => x"C0C0C0F980F8F8F8",
 18778 => x"C0C0C0F980F8F880",
 18779 => x"C0C0C0F980F8F890",
 18780 => x"C0C0C0F980F880C0",
 18781 => x"C0C0C0F980F880F9",
 18782 => x"C0C0C0F980F880A4",
 18783 => x"C0C0C0F980F880B0",
 18784 => x"C0C0C0F980F88099",
 18785 => x"C0C0C0F980F88092",
 18786 => x"C0C0C0F980F88082",
 18787 => x"C0C0C0F980F880F8",
 18788 => x"C0C0C0F980F88080",
 18789 => x"C0C0C0F980F88090",
 18790 => x"C0C0C0F980F890C0",
 18791 => x"C0C0C0F980F890F9",
 18792 => x"C0C0C0F980F890A4",
 18793 => x"C0C0C0F980F890B0",
 18794 => x"C0C0C0F980F89099",
 18795 => x"C0C0C0F980F89092",
 18796 => x"C0C0C0F980F89082",
 18797 => x"C0C0C0F980F890F8",
 18798 => x"C0C0C0F980F89080",
 18799 => x"C0C0C0F980F89090",
 18800 => x"C0C0C0F98080C0C0",
 18801 => x"C0C0C0F98080C0F9",
 18802 => x"C0C0C0F98080C0A4",
 18803 => x"C0C0C0F98080C0B0",
 18804 => x"C0C0C0F98080C099",
 18805 => x"C0C0C0F98080C092",
 18806 => x"C0C0C0F98080C082",
 18807 => x"C0C0C0F98080C0F8",
 18808 => x"C0C0C0F98080C080",
 18809 => x"C0C0C0F98080C090",
 18810 => x"C0C0C0F98080F9C0",
 18811 => x"C0C0C0F98080F9F9",
 18812 => x"C0C0C0F98080F9A4",
 18813 => x"C0C0C0F98080F9B0",
 18814 => x"C0C0C0F98080F999",
 18815 => x"C0C0C0F98080F992",
 18816 => x"C0C0C0F98080F982",
 18817 => x"C0C0C0F98080F9F8",
 18818 => x"C0C0C0F98080F980",
 18819 => x"C0C0C0F98080F990",
 18820 => x"C0C0C0F98080A4C0",
 18821 => x"C0C0C0F98080A4F9",
 18822 => x"C0C0C0F98080A4A4",
 18823 => x"C0C0C0F98080A4B0",
 18824 => x"C0C0C0F98080A499",
 18825 => x"C0C0C0F98080A492",
 18826 => x"C0C0C0F98080A482",
 18827 => x"C0C0C0F98080A4F8",
 18828 => x"C0C0C0F98080A480",
 18829 => x"C0C0C0F98080A490",
 18830 => x"C0C0C0F98080B0C0",
 18831 => x"C0C0C0F98080B0F9",
 18832 => x"C0C0C0F98080B0A4",
 18833 => x"C0C0C0F98080B0B0",
 18834 => x"C0C0C0F98080B099",
 18835 => x"C0C0C0F98080B092",
 18836 => x"C0C0C0F98080B082",
 18837 => x"C0C0C0F98080B0F8",
 18838 => x"C0C0C0F98080B080",
 18839 => x"C0C0C0F98080B090",
 18840 => x"C0C0C0F9808099C0",
 18841 => x"C0C0C0F9808099F9",
 18842 => x"C0C0C0F9808099A4",
 18843 => x"C0C0C0F9808099B0",
 18844 => x"C0C0C0F980809999",
 18845 => x"C0C0C0F980809992",
 18846 => x"C0C0C0F980809982",
 18847 => x"C0C0C0F9808099F8",
 18848 => x"C0C0C0F980809980",
 18849 => x"C0C0C0F980809990",
 18850 => x"C0C0C0F9808092C0",
 18851 => x"C0C0C0F9808092F9",
 18852 => x"C0C0C0F9808092A4",
 18853 => x"C0C0C0F9808092B0",
 18854 => x"C0C0C0F980809299",
 18855 => x"C0C0C0F980809292",
 18856 => x"C0C0C0F980809282",
 18857 => x"C0C0C0F9808092F8",
 18858 => x"C0C0C0F980809280",
 18859 => x"C0C0C0F980809290",
 18860 => x"C0C0C0F9808082C0",
 18861 => x"C0C0C0F9808082F9",
 18862 => x"C0C0C0F9808082A4",
 18863 => x"C0C0C0F9808082B0",
 18864 => x"C0C0C0F980808299",
 18865 => x"C0C0C0F980808292",
 18866 => x"C0C0C0F980808282",
 18867 => x"C0C0C0F9808082F8",
 18868 => x"C0C0C0F980808280",
 18869 => x"C0C0C0F980808290",
 18870 => x"C0C0C0F98080F8C0",
 18871 => x"C0C0C0F98080F8F9",
 18872 => x"C0C0C0F98080F8A4",
 18873 => x"C0C0C0F98080F8B0",
 18874 => x"C0C0C0F98080F899",
 18875 => x"C0C0C0F98080F892",
 18876 => x"C0C0C0F98080F882",
 18877 => x"C0C0C0F98080F8F8",
 18878 => x"C0C0C0F98080F880",
 18879 => x"C0C0C0F98080F890",
 18880 => x"C0C0C0F9808080C0",
 18881 => x"C0C0C0F9808080F9",
 18882 => x"C0C0C0F9808080A4",
 18883 => x"C0C0C0F9808080B0",
 18884 => x"C0C0C0F980808099",
 18885 => x"C0C0C0F980808092",
 18886 => x"C0C0C0F980808082",
 18887 => x"C0C0C0F9808080F8",
 18888 => x"C0C0C0F980808080",
 18889 => x"C0C0C0F980808090",
 18890 => x"C0C0C0F9808090C0",
 18891 => x"C0C0C0F9808090F9",
 18892 => x"C0C0C0F9808090A4",
 18893 => x"C0C0C0F9808090B0",
 18894 => x"C0C0C0F980809099",
 18895 => x"C0C0C0F980809092",
 18896 => x"C0C0C0F980809082",
 18897 => x"C0C0C0F9808090F8",
 18898 => x"C0C0C0F980809080",
 18899 => x"C0C0C0F980809090",
 18900 => x"C0C0C0F98090C0C0",
 18901 => x"C0C0C0F98090C0F9",
 18902 => x"C0C0C0F98090C0A4",
 18903 => x"C0C0C0F98090C0B0",
 18904 => x"C0C0C0F98090C099",
 18905 => x"C0C0C0F98090C092",
 18906 => x"C0C0C0F98090C082",
 18907 => x"C0C0C0F98090C0F8",
 18908 => x"C0C0C0F98090C080",
 18909 => x"C0C0C0F98090C090",
 18910 => x"C0C0C0F98090F9C0",
 18911 => x"C0C0C0F98090F9F9",
 18912 => x"C0C0C0F98090F9A4",
 18913 => x"C0C0C0F98090F9B0",
 18914 => x"C0C0C0F98090F999",
 18915 => x"C0C0C0F98090F992",
 18916 => x"C0C0C0F98090F982",
 18917 => x"C0C0C0F98090F9F8",
 18918 => x"C0C0C0F98090F980",
 18919 => x"C0C0C0F98090F990",
 18920 => x"C0C0C0F98090A4C0",
 18921 => x"C0C0C0F98090A4F9",
 18922 => x"C0C0C0F98090A4A4",
 18923 => x"C0C0C0F98090A4B0",
 18924 => x"C0C0C0F98090A499",
 18925 => x"C0C0C0F98090A492",
 18926 => x"C0C0C0F98090A482",
 18927 => x"C0C0C0F98090A4F8",
 18928 => x"C0C0C0F98090A480",
 18929 => x"C0C0C0F98090A490",
 18930 => x"C0C0C0F98090B0C0",
 18931 => x"C0C0C0F98090B0F9",
 18932 => x"C0C0C0F98090B0A4",
 18933 => x"C0C0C0F98090B0B0",
 18934 => x"C0C0C0F98090B099",
 18935 => x"C0C0C0F98090B092",
 18936 => x"C0C0C0F98090B082",
 18937 => x"C0C0C0F98090B0F8",
 18938 => x"C0C0C0F98090B080",
 18939 => x"C0C0C0F98090B090",
 18940 => x"C0C0C0F9809099C0",
 18941 => x"C0C0C0F9809099F9",
 18942 => x"C0C0C0F9809099A4",
 18943 => x"C0C0C0F9809099B0",
 18944 => x"C0C0C0F980909999",
 18945 => x"C0C0C0F980909992",
 18946 => x"C0C0C0F980909982",
 18947 => x"C0C0C0F9809099F8",
 18948 => x"C0C0C0F980909980",
 18949 => x"C0C0C0F980909990",
 18950 => x"C0C0C0F9809092C0",
 18951 => x"C0C0C0F9809092F9",
 18952 => x"C0C0C0F9809092A4",
 18953 => x"C0C0C0F9809092B0",
 18954 => x"C0C0C0F980909299",
 18955 => x"C0C0C0F980909292",
 18956 => x"C0C0C0F980909282",
 18957 => x"C0C0C0F9809092F8",
 18958 => x"C0C0C0F980909280",
 18959 => x"C0C0C0F980909290",
 18960 => x"C0C0C0F9809082C0",
 18961 => x"C0C0C0F9809082F9",
 18962 => x"C0C0C0F9809082A4",
 18963 => x"C0C0C0F9809082B0",
 18964 => x"C0C0C0F980908299",
 18965 => x"C0C0C0F980908292",
 18966 => x"C0C0C0F980908282",
 18967 => x"C0C0C0F9809082F8",
 18968 => x"C0C0C0F980908280",
 18969 => x"C0C0C0F980908290",
 18970 => x"C0C0C0F98090F8C0",
 18971 => x"C0C0C0F98090F8F9",
 18972 => x"C0C0C0F98090F8A4",
 18973 => x"C0C0C0F98090F8B0",
 18974 => x"C0C0C0F98090F899",
 18975 => x"C0C0C0F98090F892",
 18976 => x"C0C0C0F98090F882",
 18977 => x"C0C0C0F98090F8F8",
 18978 => x"C0C0C0F98090F880",
 18979 => x"C0C0C0F98090F890",
 18980 => x"C0C0C0F9809080C0",
 18981 => x"C0C0C0F9809080F9",
 18982 => x"C0C0C0F9809080A4",
 18983 => x"C0C0C0F9809080B0",
 18984 => x"C0C0C0F980908099",
 18985 => x"C0C0C0F980908092",
 18986 => x"C0C0C0F980908082",
 18987 => x"C0C0C0F9809080F8",
 18988 => x"C0C0C0F980908080",
 18989 => x"C0C0C0F980908090",
 18990 => x"C0C0C0F9809090C0",
 18991 => x"C0C0C0F9809090F9",
 18992 => x"C0C0C0F9809090A4",
 18993 => x"C0C0C0F9809090B0",
 18994 => x"C0C0C0F980909099",
 18995 => x"C0C0C0F980909092",
 18996 => x"C0C0C0F980909082",
 18997 => x"C0C0C0F9809090F8",
 18998 => x"C0C0C0F980909080",
 18999 => x"C0C0C0F980909090",
 19000 => x"C0C0C0F990C0C0C0",
 19001 => x"C0C0C0F990C0C0F9",
 19002 => x"C0C0C0F990C0C0A4",
 19003 => x"C0C0C0F990C0C0B0",
 19004 => x"C0C0C0F990C0C099",
 19005 => x"C0C0C0F990C0C092",
 19006 => x"C0C0C0F990C0C082",
 19007 => x"C0C0C0F990C0C0F8",
 19008 => x"C0C0C0F990C0C080",
 19009 => x"C0C0C0F990C0C090",
 19010 => x"C0C0C0F990C0F9C0",
 19011 => x"C0C0C0F990C0F9F9",
 19012 => x"C0C0C0F990C0F9A4",
 19013 => x"C0C0C0F990C0F9B0",
 19014 => x"C0C0C0F990C0F999",
 19015 => x"C0C0C0F990C0F992",
 19016 => x"C0C0C0F990C0F982",
 19017 => x"C0C0C0F990C0F9F8",
 19018 => x"C0C0C0F990C0F980",
 19019 => x"C0C0C0F990C0F990",
 19020 => x"C0C0C0F990C0A4C0",
 19021 => x"C0C0C0F990C0A4F9",
 19022 => x"C0C0C0F990C0A4A4",
 19023 => x"C0C0C0F990C0A4B0",
 19024 => x"C0C0C0F990C0A499",
 19025 => x"C0C0C0F990C0A492",
 19026 => x"C0C0C0F990C0A482",
 19027 => x"C0C0C0F990C0A4F8",
 19028 => x"C0C0C0F990C0A480",
 19029 => x"C0C0C0F990C0A490",
 19030 => x"C0C0C0F990C0B0C0",
 19031 => x"C0C0C0F990C0B0F9",
 19032 => x"C0C0C0F990C0B0A4",
 19033 => x"C0C0C0F990C0B0B0",
 19034 => x"C0C0C0F990C0B099",
 19035 => x"C0C0C0F990C0B092",
 19036 => x"C0C0C0F990C0B082",
 19037 => x"C0C0C0F990C0B0F8",
 19038 => x"C0C0C0F990C0B080",
 19039 => x"C0C0C0F990C0B090",
 19040 => x"C0C0C0F990C099C0",
 19041 => x"C0C0C0F990C099F9",
 19042 => x"C0C0C0F990C099A4",
 19043 => x"C0C0C0F990C099B0",
 19044 => x"C0C0C0F990C09999",
 19045 => x"C0C0C0F990C09992",
 19046 => x"C0C0C0F990C09982",
 19047 => x"C0C0C0F990C099F8",
 19048 => x"C0C0C0F990C09980",
 19049 => x"C0C0C0F990C09990",
 19050 => x"C0C0C0F990C092C0",
 19051 => x"C0C0C0F990C092F9",
 19052 => x"C0C0C0F990C092A4",
 19053 => x"C0C0C0F990C092B0",
 19054 => x"C0C0C0F990C09299",
 19055 => x"C0C0C0F990C09292",
 19056 => x"C0C0C0F990C09282",
 19057 => x"C0C0C0F990C092F8",
 19058 => x"C0C0C0F990C09280",
 19059 => x"C0C0C0F990C09290",
 19060 => x"C0C0C0F990C082C0",
 19061 => x"C0C0C0F990C082F9",
 19062 => x"C0C0C0F990C082A4",
 19063 => x"C0C0C0F990C082B0",
 19064 => x"C0C0C0F990C08299",
 19065 => x"C0C0C0F990C08292",
 19066 => x"C0C0C0F990C08282",
 19067 => x"C0C0C0F990C082F8",
 19068 => x"C0C0C0F990C08280",
 19069 => x"C0C0C0F990C08290",
 19070 => x"C0C0C0F990C0F8C0",
 19071 => x"C0C0C0F990C0F8F9",
 19072 => x"C0C0C0F990C0F8A4",
 19073 => x"C0C0C0F990C0F8B0",
 19074 => x"C0C0C0F990C0F899",
 19075 => x"C0C0C0F990C0F892",
 19076 => x"C0C0C0F990C0F882",
 19077 => x"C0C0C0F990C0F8F8",
 19078 => x"C0C0C0F990C0F880",
 19079 => x"C0C0C0F990C0F890",
 19080 => x"C0C0C0F990C080C0",
 19081 => x"C0C0C0F990C080F9",
 19082 => x"C0C0C0F990C080A4",
 19083 => x"C0C0C0F990C080B0",
 19084 => x"C0C0C0F990C08099",
 19085 => x"C0C0C0F990C08092",
 19086 => x"C0C0C0F990C08082",
 19087 => x"C0C0C0F990C080F8",
 19088 => x"C0C0C0F990C08080",
 19089 => x"C0C0C0F990C08090",
 19090 => x"C0C0C0F990C090C0",
 19091 => x"C0C0C0F990C090F9",
 19092 => x"C0C0C0F990C090A4",
 19093 => x"C0C0C0F990C090B0",
 19094 => x"C0C0C0F990C09099",
 19095 => x"C0C0C0F990C09092",
 19096 => x"C0C0C0F990C09082",
 19097 => x"C0C0C0F990C090F8",
 19098 => x"C0C0C0F990C09080",
 19099 => x"C0C0C0F990C09090",
 19100 => x"C0C0C0F990F9C0C0",
 19101 => x"C0C0C0F990F9C0F9",
 19102 => x"C0C0C0F990F9C0A4",
 19103 => x"C0C0C0F990F9C0B0",
 19104 => x"C0C0C0F990F9C099",
 19105 => x"C0C0C0F990F9C092",
 19106 => x"C0C0C0F990F9C082",
 19107 => x"C0C0C0F990F9C0F8",
 19108 => x"C0C0C0F990F9C080",
 19109 => x"C0C0C0F990F9C090",
 19110 => x"C0C0C0F990F9F9C0",
 19111 => x"C0C0C0F990F9F9F9",
 19112 => x"C0C0C0F990F9F9A4",
 19113 => x"C0C0C0F990F9F9B0",
 19114 => x"C0C0C0F990F9F999",
 19115 => x"C0C0C0F990F9F992",
 19116 => x"C0C0C0F990F9F982",
 19117 => x"C0C0C0F990F9F9F8",
 19118 => x"C0C0C0F990F9F980",
 19119 => x"C0C0C0F990F9F990",
 19120 => x"C0C0C0F990F9A4C0",
 19121 => x"C0C0C0F990F9A4F9",
 19122 => x"C0C0C0F990F9A4A4",
 19123 => x"C0C0C0F990F9A4B0",
 19124 => x"C0C0C0F990F9A499",
 19125 => x"C0C0C0F990F9A492",
 19126 => x"C0C0C0F990F9A482",
 19127 => x"C0C0C0F990F9A4F8",
 19128 => x"C0C0C0F990F9A480",
 19129 => x"C0C0C0F990F9A490",
 19130 => x"C0C0C0F990F9B0C0",
 19131 => x"C0C0C0F990F9B0F9",
 19132 => x"C0C0C0F990F9B0A4",
 19133 => x"C0C0C0F990F9B0B0",
 19134 => x"C0C0C0F990F9B099",
 19135 => x"C0C0C0F990F9B092",
 19136 => x"C0C0C0F990F9B082",
 19137 => x"C0C0C0F990F9B0F8",
 19138 => x"C0C0C0F990F9B080",
 19139 => x"C0C0C0F990F9B090",
 19140 => x"C0C0C0F990F999C0",
 19141 => x"C0C0C0F990F999F9",
 19142 => x"C0C0C0F990F999A4",
 19143 => x"C0C0C0F990F999B0",
 19144 => x"C0C0C0F990F99999",
 19145 => x"C0C0C0F990F99992",
 19146 => x"C0C0C0F990F99982",
 19147 => x"C0C0C0F990F999F8",
 19148 => x"C0C0C0F990F99980",
 19149 => x"C0C0C0F990F99990",
 19150 => x"C0C0C0F990F992C0",
 19151 => x"C0C0C0F990F992F9",
 19152 => x"C0C0C0F990F992A4",
 19153 => x"C0C0C0F990F992B0",
 19154 => x"C0C0C0F990F99299",
 19155 => x"C0C0C0F990F99292",
 19156 => x"C0C0C0F990F99282",
 19157 => x"C0C0C0F990F992F8",
 19158 => x"C0C0C0F990F99280",
 19159 => x"C0C0C0F990F99290",
 19160 => x"C0C0C0F990F982C0",
 19161 => x"C0C0C0F990F982F9",
 19162 => x"C0C0C0F990F982A4",
 19163 => x"C0C0C0F990F982B0",
 19164 => x"C0C0C0F990F98299",
 19165 => x"C0C0C0F990F98292",
 19166 => x"C0C0C0F990F98282",
 19167 => x"C0C0C0F990F982F8",
 19168 => x"C0C0C0F990F98280",
 19169 => x"C0C0C0F990F98290",
 19170 => x"C0C0C0F990F9F8C0",
 19171 => x"C0C0C0F990F9F8F9",
 19172 => x"C0C0C0F990F9F8A4",
 19173 => x"C0C0C0F990F9F8B0",
 19174 => x"C0C0C0F990F9F899",
 19175 => x"C0C0C0F990F9F892",
 19176 => x"C0C0C0F990F9F882",
 19177 => x"C0C0C0F990F9F8F8",
 19178 => x"C0C0C0F990F9F880",
 19179 => x"C0C0C0F990F9F890",
 19180 => x"C0C0C0F990F980C0",
 19181 => x"C0C0C0F990F980F9",
 19182 => x"C0C0C0F990F980A4",
 19183 => x"C0C0C0F990F980B0",
 19184 => x"C0C0C0F990F98099",
 19185 => x"C0C0C0F990F98092",
 19186 => x"C0C0C0F990F98082",
 19187 => x"C0C0C0F990F980F8",
 19188 => x"C0C0C0F990F98080",
 19189 => x"C0C0C0F990F98090",
 19190 => x"C0C0C0F990F990C0",
 19191 => x"C0C0C0F990F990F9",
 19192 => x"C0C0C0F990F990A4",
 19193 => x"C0C0C0F990F990B0",
 19194 => x"C0C0C0F990F99099",
 19195 => x"C0C0C0F990F99092",
 19196 => x"C0C0C0F990F99082",
 19197 => x"C0C0C0F990F990F8",
 19198 => x"C0C0C0F990F99080",
 19199 => x"C0C0C0F990F99090",
 19200 => x"C0C0C0F990A4C0C0",
 19201 => x"C0C0C0F990A4C0F9",
 19202 => x"C0C0C0F990A4C0A4",
 19203 => x"C0C0C0F990A4C0B0",
 19204 => x"C0C0C0F990A4C099",
 19205 => x"C0C0C0F990A4C092",
 19206 => x"C0C0C0F990A4C082",
 19207 => x"C0C0C0F990A4C0F8",
 19208 => x"C0C0C0F990A4C080",
 19209 => x"C0C0C0F990A4C090",
 19210 => x"C0C0C0F990A4F9C0",
 19211 => x"C0C0C0F990A4F9F9",
 19212 => x"C0C0C0F990A4F9A4",
 19213 => x"C0C0C0F990A4F9B0",
 19214 => x"C0C0C0F990A4F999",
 19215 => x"C0C0C0F990A4F992",
 19216 => x"C0C0C0F990A4F982",
 19217 => x"C0C0C0F990A4F9F8",
 19218 => x"C0C0C0F990A4F980",
 19219 => x"C0C0C0F990A4F990",
 19220 => x"C0C0C0F990A4A4C0",
 19221 => x"C0C0C0F990A4A4F9",
 19222 => x"C0C0C0F990A4A4A4",
 19223 => x"C0C0C0F990A4A4B0",
 19224 => x"C0C0C0F990A4A499",
 19225 => x"C0C0C0F990A4A492",
 19226 => x"C0C0C0F990A4A482",
 19227 => x"C0C0C0F990A4A4F8",
 19228 => x"C0C0C0F990A4A480",
 19229 => x"C0C0C0F990A4A490",
 19230 => x"C0C0C0F990A4B0C0",
 19231 => x"C0C0C0F990A4B0F9",
 19232 => x"C0C0C0F990A4B0A4",
 19233 => x"C0C0C0F990A4B0B0",
 19234 => x"C0C0C0F990A4B099",
 19235 => x"C0C0C0F990A4B092",
 19236 => x"C0C0C0F990A4B082",
 19237 => x"C0C0C0F990A4B0F8",
 19238 => x"C0C0C0F990A4B080",
 19239 => x"C0C0C0F990A4B090",
 19240 => x"C0C0C0F990A499C0",
 19241 => x"C0C0C0F990A499F9",
 19242 => x"C0C0C0F990A499A4",
 19243 => x"C0C0C0F990A499B0",
 19244 => x"C0C0C0F990A49999",
 19245 => x"C0C0C0F990A49992",
 19246 => x"C0C0C0F990A49982",
 19247 => x"C0C0C0F990A499F8",
 19248 => x"C0C0C0F990A49980",
 19249 => x"C0C0C0F990A49990",
 19250 => x"C0C0C0F990A492C0",
 19251 => x"C0C0C0F990A492F9",
 19252 => x"C0C0C0F990A492A4",
 19253 => x"C0C0C0F990A492B0",
 19254 => x"C0C0C0F990A49299",
 19255 => x"C0C0C0F990A49292",
 19256 => x"C0C0C0F990A49282",
 19257 => x"C0C0C0F990A492F8",
 19258 => x"C0C0C0F990A49280",
 19259 => x"C0C0C0F990A49290",
 19260 => x"C0C0C0F990A482C0",
 19261 => x"C0C0C0F990A482F9",
 19262 => x"C0C0C0F990A482A4",
 19263 => x"C0C0C0F990A482B0",
 19264 => x"C0C0C0F990A48299",
 19265 => x"C0C0C0F990A48292",
 19266 => x"C0C0C0F990A48282",
 19267 => x"C0C0C0F990A482F8",
 19268 => x"C0C0C0F990A48280",
 19269 => x"C0C0C0F990A48290",
 19270 => x"C0C0C0F990A4F8C0",
 19271 => x"C0C0C0F990A4F8F9",
 19272 => x"C0C0C0F990A4F8A4",
 19273 => x"C0C0C0F990A4F8B0",
 19274 => x"C0C0C0F990A4F899",
 19275 => x"C0C0C0F990A4F892",
 19276 => x"C0C0C0F990A4F882",
 19277 => x"C0C0C0F990A4F8F8",
 19278 => x"C0C0C0F990A4F880",
 19279 => x"C0C0C0F990A4F890",
 19280 => x"C0C0C0F990A480C0",
 19281 => x"C0C0C0F990A480F9",
 19282 => x"C0C0C0F990A480A4",
 19283 => x"C0C0C0F990A480B0",
 19284 => x"C0C0C0F990A48099",
 19285 => x"C0C0C0F990A48092",
 19286 => x"C0C0C0F990A48082",
 19287 => x"C0C0C0F990A480F8",
 19288 => x"C0C0C0F990A48080",
 19289 => x"C0C0C0F990A48090",
 19290 => x"C0C0C0F990A490C0",
 19291 => x"C0C0C0F990A490F9",
 19292 => x"C0C0C0F990A490A4",
 19293 => x"C0C0C0F990A490B0",
 19294 => x"C0C0C0F990A49099",
 19295 => x"C0C0C0F990A49092",
 19296 => x"C0C0C0F990A49082",
 19297 => x"C0C0C0F990A490F8",
 19298 => x"C0C0C0F990A49080",
 19299 => x"C0C0C0F990A49090",
 19300 => x"C0C0C0F990B0C0C0",
 19301 => x"C0C0C0F990B0C0F9",
 19302 => x"C0C0C0F990B0C0A4",
 19303 => x"C0C0C0F990B0C0B0",
 19304 => x"C0C0C0F990B0C099",
 19305 => x"C0C0C0F990B0C092",
 19306 => x"C0C0C0F990B0C082",
 19307 => x"C0C0C0F990B0C0F8",
 19308 => x"C0C0C0F990B0C080",
 19309 => x"C0C0C0F990B0C090",
 19310 => x"C0C0C0F990B0F9C0",
 19311 => x"C0C0C0F990B0F9F9",
 19312 => x"C0C0C0F990B0F9A4",
 19313 => x"C0C0C0F990B0F9B0",
 19314 => x"C0C0C0F990B0F999",
 19315 => x"C0C0C0F990B0F992",
 19316 => x"C0C0C0F990B0F982",
 19317 => x"C0C0C0F990B0F9F8",
 19318 => x"C0C0C0F990B0F980",
 19319 => x"C0C0C0F990B0F990",
 19320 => x"C0C0C0F990B0A4C0",
 19321 => x"C0C0C0F990B0A4F9",
 19322 => x"C0C0C0F990B0A4A4",
 19323 => x"C0C0C0F990B0A4B0",
 19324 => x"C0C0C0F990B0A499",
 19325 => x"C0C0C0F990B0A492",
 19326 => x"C0C0C0F990B0A482",
 19327 => x"C0C0C0F990B0A4F8",
 19328 => x"C0C0C0F990B0A480",
 19329 => x"C0C0C0F990B0A490",
 19330 => x"C0C0C0F990B0B0C0",
 19331 => x"C0C0C0F990B0B0F9",
 19332 => x"C0C0C0F990B0B0A4",
 19333 => x"C0C0C0F990B0B0B0",
 19334 => x"C0C0C0F990B0B099",
 19335 => x"C0C0C0F990B0B092",
 19336 => x"C0C0C0F990B0B082",
 19337 => x"C0C0C0F990B0B0F8",
 19338 => x"C0C0C0F990B0B080",
 19339 => x"C0C0C0F990B0B090",
 19340 => x"C0C0C0F990B099C0",
 19341 => x"C0C0C0F990B099F9",
 19342 => x"C0C0C0F990B099A4",
 19343 => x"C0C0C0F990B099B0",
 19344 => x"C0C0C0F990B09999",
 19345 => x"C0C0C0F990B09992",
 19346 => x"C0C0C0F990B09982",
 19347 => x"C0C0C0F990B099F8",
 19348 => x"C0C0C0F990B09980",
 19349 => x"C0C0C0F990B09990",
 19350 => x"C0C0C0F990B092C0",
 19351 => x"C0C0C0F990B092F9",
 19352 => x"C0C0C0F990B092A4",
 19353 => x"C0C0C0F990B092B0",
 19354 => x"C0C0C0F990B09299",
 19355 => x"C0C0C0F990B09292",
 19356 => x"C0C0C0F990B09282",
 19357 => x"C0C0C0F990B092F8",
 19358 => x"C0C0C0F990B09280",
 19359 => x"C0C0C0F990B09290",
 19360 => x"C0C0C0F990B082C0",
 19361 => x"C0C0C0F990B082F9",
 19362 => x"C0C0C0F990B082A4",
 19363 => x"C0C0C0F990B082B0",
 19364 => x"C0C0C0F990B08299",
 19365 => x"C0C0C0F990B08292",
 19366 => x"C0C0C0F990B08282",
 19367 => x"C0C0C0F990B082F8",
 19368 => x"C0C0C0F990B08280",
 19369 => x"C0C0C0F990B08290",
 19370 => x"C0C0C0F990B0F8C0",
 19371 => x"C0C0C0F990B0F8F9",
 19372 => x"C0C0C0F990B0F8A4",
 19373 => x"C0C0C0F990B0F8B0",
 19374 => x"C0C0C0F990B0F899",
 19375 => x"C0C0C0F990B0F892",
 19376 => x"C0C0C0F990B0F882",
 19377 => x"C0C0C0F990B0F8F8",
 19378 => x"C0C0C0F990B0F880",
 19379 => x"C0C0C0F990B0F890",
 19380 => x"C0C0C0F990B080C0",
 19381 => x"C0C0C0F990B080F9",
 19382 => x"C0C0C0F990B080A4",
 19383 => x"C0C0C0F990B080B0",
 19384 => x"C0C0C0F990B08099",
 19385 => x"C0C0C0F990B08092",
 19386 => x"C0C0C0F990B08082",
 19387 => x"C0C0C0F990B080F8",
 19388 => x"C0C0C0F990B08080",
 19389 => x"C0C0C0F990B08090",
 19390 => x"C0C0C0F990B090C0",
 19391 => x"C0C0C0F990B090F9",
 19392 => x"C0C0C0F990B090A4",
 19393 => x"C0C0C0F990B090B0",
 19394 => x"C0C0C0F990B09099",
 19395 => x"C0C0C0F990B09092",
 19396 => x"C0C0C0F990B09082",
 19397 => x"C0C0C0F990B090F8",
 19398 => x"C0C0C0F990B09080",
 19399 => x"C0C0C0F990B09090",
 19400 => x"C0C0C0F99099C0C0",
 19401 => x"C0C0C0F99099C0F9",
 19402 => x"C0C0C0F99099C0A4",
 19403 => x"C0C0C0F99099C0B0",
 19404 => x"C0C0C0F99099C099",
 19405 => x"C0C0C0F99099C092",
 19406 => x"C0C0C0F99099C082",
 19407 => x"C0C0C0F99099C0F8",
 19408 => x"C0C0C0F99099C080",
 19409 => x"C0C0C0F99099C090",
 19410 => x"C0C0C0F99099F9C0",
 19411 => x"C0C0C0F99099F9F9",
 19412 => x"C0C0C0F99099F9A4",
 19413 => x"C0C0C0F99099F9B0",
 19414 => x"C0C0C0F99099F999",
 19415 => x"C0C0C0F99099F992",
 19416 => x"C0C0C0F99099F982",
 19417 => x"C0C0C0F99099F9F8",
 19418 => x"C0C0C0F99099F980",
 19419 => x"C0C0C0F99099F990",
 19420 => x"C0C0C0F99099A4C0",
 19421 => x"C0C0C0F99099A4F9",
 19422 => x"C0C0C0F99099A4A4",
 19423 => x"C0C0C0F99099A4B0",
 19424 => x"C0C0C0F99099A499",
 19425 => x"C0C0C0F99099A492",
 19426 => x"C0C0C0F99099A482",
 19427 => x"C0C0C0F99099A4F8",
 19428 => x"C0C0C0F99099A480",
 19429 => x"C0C0C0F99099A490",
 19430 => x"C0C0C0F99099B0C0",
 19431 => x"C0C0C0F99099B0F9",
 19432 => x"C0C0C0F99099B0A4",
 19433 => x"C0C0C0F99099B0B0",
 19434 => x"C0C0C0F99099B099",
 19435 => x"C0C0C0F99099B092",
 19436 => x"C0C0C0F99099B082",
 19437 => x"C0C0C0F99099B0F8",
 19438 => x"C0C0C0F99099B080",
 19439 => x"C0C0C0F99099B090",
 19440 => x"C0C0C0F9909999C0",
 19441 => x"C0C0C0F9909999F9",
 19442 => x"C0C0C0F9909999A4",
 19443 => x"C0C0C0F9909999B0",
 19444 => x"C0C0C0F990999999",
 19445 => x"C0C0C0F990999992",
 19446 => x"C0C0C0F990999982",
 19447 => x"C0C0C0F9909999F8",
 19448 => x"C0C0C0F990999980",
 19449 => x"C0C0C0F990999990",
 19450 => x"C0C0C0F9909992C0",
 19451 => x"C0C0C0F9909992F9",
 19452 => x"C0C0C0F9909992A4",
 19453 => x"C0C0C0F9909992B0",
 19454 => x"C0C0C0F990999299",
 19455 => x"C0C0C0F990999292",
 19456 => x"C0C0C0F990999282",
 19457 => x"C0C0C0F9909992F8",
 19458 => x"C0C0C0F990999280",
 19459 => x"C0C0C0F990999290",
 19460 => x"C0C0C0F9909982C0",
 19461 => x"C0C0C0F9909982F9",
 19462 => x"C0C0C0F9909982A4",
 19463 => x"C0C0C0F9909982B0",
 19464 => x"C0C0C0F990998299",
 19465 => x"C0C0C0F990998292",
 19466 => x"C0C0C0F990998282",
 19467 => x"C0C0C0F9909982F8",
 19468 => x"C0C0C0F990998280",
 19469 => x"C0C0C0F990998290",
 19470 => x"C0C0C0F99099F8C0",
 19471 => x"C0C0C0F99099F8F9",
 19472 => x"C0C0C0F99099F8A4",
 19473 => x"C0C0C0F99099F8B0",
 19474 => x"C0C0C0F99099F899",
 19475 => x"C0C0C0F99099F892",
 19476 => x"C0C0C0F99099F882",
 19477 => x"C0C0C0F99099F8F8",
 19478 => x"C0C0C0F99099F880",
 19479 => x"C0C0C0F99099F890",
 19480 => x"C0C0C0F9909980C0",
 19481 => x"C0C0C0F9909980F9",
 19482 => x"C0C0C0F9909980A4",
 19483 => x"C0C0C0F9909980B0",
 19484 => x"C0C0C0F990998099",
 19485 => x"C0C0C0F990998092",
 19486 => x"C0C0C0F990998082",
 19487 => x"C0C0C0F9909980F8",
 19488 => x"C0C0C0F990998080",
 19489 => x"C0C0C0F990998090",
 19490 => x"C0C0C0F9909990C0",
 19491 => x"C0C0C0F9909990F9",
 19492 => x"C0C0C0F9909990A4",
 19493 => x"C0C0C0F9909990B0",
 19494 => x"C0C0C0F990999099",
 19495 => x"C0C0C0F990999092",
 19496 => x"C0C0C0F990999082",
 19497 => x"C0C0C0F9909990F8",
 19498 => x"C0C0C0F990999080",
 19499 => x"C0C0C0F990999090",
 19500 => x"C0C0C0F99092C0C0",
 19501 => x"C0C0C0F99092C0F9",
 19502 => x"C0C0C0F99092C0A4",
 19503 => x"C0C0C0F99092C0B0",
 19504 => x"C0C0C0F99092C099",
 19505 => x"C0C0C0F99092C092",
 19506 => x"C0C0C0F99092C082",
 19507 => x"C0C0C0F99092C0F8",
 19508 => x"C0C0C0F99092C080",
 19509 => x"C0C0C0F99092C090",
 19510 => x"C0C0C0F99092F9C0",
 19511 => x"C0C0C0F99092F9F9",
 19512 => x"C0C0C0F99092F9A4",
 19513 => x"C0C0C0F99092F9B0",
 19514 => x"C0C0C0F99092F999",
 19515 => x"C0C0C0F99092F992",
 19516 => x"C0C0C0F99092F982",
 19517 => x"C0C0C0F99092F9F8",
 19518 => x"C0C0C0F99092F980",
 19519 => x"C0C0C0F99092F990",
 19520 => x"C0C0C0F99092A4C0",
 19521 => x"C0C0C0F99092A4F9",
 19522 => x"C0C0C0F99092A4A4",
 19523 => x"C0C0C0F99092A4B0",
 19524 => x"C0C0C0F99092A499",
 19525 => x"C0C0C0F99092A492",
 19526 => x"C0C0C0F99092A482",
 19527 => x"C0C0C0F99092A4F8",
 19528 => x"C0C0C0F99092A480",
 19529 => x"C0C0C0F99092A490",
 19530 => x"C0C0C0F99092B0C0",
 19531 => x"C0C0C0F99092B0F9",
 19532 => x"C0C0C0F99092B0A4",
 19533 => x"C0C0C0F99092B0B0",
 19534 => x"C0C0C0F99092B099",
 19535 => x"C0C0C0F99092B092",
 19536 => x"C0C0C0F99092B082",
 19537 => x"C0C0C0F99092B0F8",
 19538 => x"C0C0C0F99092B080",
 19539 => x"C0C0C0F99092B090",
 19540 => x"C0C0C0F9909299C0",
 19541 => x"C0C0C0F9909299F9",
 19542 => x"C0C0C0F9909299A4",
 19543 => x"C0C0C0F9909299B0",
 19544 => x"C0C0C0F990929999",
 19545 => x"C0C0C0F990929992",
 19546 => x"C0C0C0F990929982",
 19547 => x"C0C0C0F9909299F8",
 19548 => x"C0C0C0F990929980",
 19549 => x"C0C0C0F990929990",
 19550 => x"C0C0C0F9909292C0",
 19551 => x"C0C0C0F9909292F9",
 19552 => x"C0C0C0F9909292A4",
 19553 => x"C0C0C0F9909292B0",
 19554 => x"C0C0C0F990929299",
 19555 => x"C0C0C0F990929292",
 19556 => x"C0C0C0F990929282",
 19557 => x"C0C0C0F9909292F8",
 19558 => x"C0C0C0F990929280",
 19559 => x"C0C0C0F990929290",
 19560 => x"C0C0C0F9909282C0",
 19561 => x"C0C0C0F9909282F9",
 19562 => x"C0C0C0F9909282A4",
 19563 => x"C0C0C0F9909282B0",
 19564 => x"C0C0C0F990928299",
 19565 => x"C0C0C0F990928292",
 19566 => x"C0C0C0F990928282",
 19567 => x"C0C0C0F9909282F8",
 19568 => x"C0C0C0F990928280",
 19569 => x"C0C0C0F990928290",
 19570 => x"C0C0C0F99092F8C0",
 19571 => x"C0C0C0F99092F8F9",
 19572 => x"C0C0C0F99092F8A4",
 19573 => x"C0C0C0F99092F8B0",
 19574 => x"C0C0C0F99092F899",
 19575 => x"C0C0C0F99092F892",
 19576 => x"C0C0C0F99092F882",
 19577 => x"C0C0C0F99092F8F8",
 19578 => x"C0C0C0F99092F880",
 19579 => x"C0C0C0F99092F890",
 19580 => x"C0C0C0F9909280C0",
 19581 => x"C0C0C0F9909280F9",
 19582 => x"C0C0C0F9909280A4",
 19583 => x"C0C0C0F9909280B0",
 19584 => x"C0C0C0F990928099",
 19585 => x"C0C0C0F990928092",
 19586 => x"C0C0C0F990928082",
 19587 => x"C0C0C0F9909280F8",
 19588 => x"C0C0C0F990928080",
 19589 => x"C0C0C0F990928090",
 19590 => x"C0C0C0F9909290C0",
 19591 => x"C0C0C0F9909290F9",
 19592 => x"C0C0C0F9909290A4",
 19593 => x"C0C0C0F9909290B0",
 19594 => x"C0C0C0F990929099",
 19595 => x"C0C0C0F990929092",
 19596 => x"C0C0C0F990929082",
 19597 => x"C0C0C0F9909290F8",
 19598 => x"C0C0C0F990929080",
 19599 => x"C0C0C0F990929090",
 19600 => x"C0C0C0F99082C0C0",
 19601 => x"C0C0C0F99082C0F9",
 19602 => x"C0C0C0F99082C0A4",
 19603 => x"C0C0C0F99082C0B0",
 19604 => x"C0C0C0F99082C099",
 19605 => x"C0C0C0F99082C092",
 19606 => x"C0C0C0F99082C082",
 19607 => x"C0C0C0F99082C0F8",
 19608 => x"C0C0C0F99082C080",
 19609 => x"C0C0C0F99082C090",
 19610 => x"C0C0C0F99082F9C0",
 19611 => x"C0C0C0F99082F9F9",
 19612 => x"C0C0C0F99082F9A4",
 19613 => x"C0C0C0F99082F9B0",
 19614 => x"C0C0C0F99082F999",
 19615 => x"C0C0C0F99082F992",
 19616 => x"C0C0C0F99082F982",
 19617 => x"C0C0C0F99082F9F8",
 19618 => x"C0C0C0F99082F980",
 19619 => x"C0C0C0F99082F990",
 19620 => x"C0C0C0F99082A4C0",
 19621 => x"C0C0C0F99082A4F9",
 19622 => x"C0C0C0F99082A4A4",
 19623 => x"C0C0C0F99082A4B0",
 19624 => x"C0C0C0F99082A499",
 19625 => x"C0C0C0F99082A492",
 19626 => x"C0C0C0F99082A482",
 19627 => x"C0C0C0F99082A4F8",
 19628 => x"C0C0C0F99082A480",
 19629 => x"C0C0C0F99082A490",
 19630 => x"C0C0C0F99082B0C0",
 19631 => x"C0C0C0F99082B0F9",
 19632 => x"C0C0C0F99082B0A4",
 19633 => x"C0C0C0F99082B0B0",
 19634 => x"C0C0C0F99082B099",
 19635 => x"C0C0C0F99082B092",
 19636 => x"C0C0C0F99082B082",
 19637 => x"C0C0C0F99082B0F8",
 19638 => x"C0C0C0F99082B080",
 19639 => x"C0C0C0F99082B090",
 19640 => x"C0C0C0F9908299C0",
 19641 => x"C0C0C0F9908299F9",
 19642 => x"C0C0C0F9908299A4",
 19643 => x"C0C0C0F9908299B0",
 19644 => x"C0C0C0F990829999",
 19645 => x"C0C0C0F990829992",
 19646 => x"C0C0C0F990829982",
 19647 => x"C0C0C0F9908299F8",
 19648 => x"C0C0C0F990829980",
 19649 => x"C0C0C0F990829990",
 19650 => x"C0C0C0F9908292C0",
 19651 => x"C0C0C0F9908292F9",
 19652 => x"C0C0C0F9908292A4",
 19653 => x"C0C0C0F9908292B0",
 19654 => x"C0C0C0F990829299",
 19655 => x"C0C0C0F990829292",
 19656 => x"C0C0C0F990829282",
 19657 => x"C0C0C0F9908292F8",
 19658 => x"C0C0C0F990829280",
 19659 => x"C0C0C0F990829290",
 19660 => x"C0C0C0F9908282C0",
 19661 => x"C0C0C0F9908282F9",
 19662 => x"C0C0C0F9908282A4",
 19663 => x"C0C0C0F9908282B0",
 19664 => x"C0C0C0F990828299",
 19665 => x"C0C0C0F990828292",
 19666 => x"C0C0C0F990828282",
 19667 => x"C0C0C0F9908282F8",
 19668 => x"C0C0C0F990828280",
 19669 => x"C0C0C0F990828290",
 19670 => x"C0C0C0F99082F8C0",
 19671 => x"C0C0C0F99082F8F9",
 19672 => x"C0C0C0F99082F8A4",
 19673 => x"C0C0C0F99082F8B0",
 19674 => x"C0C0C0F99082F899",
 19675 => x"C0C0C0F99082F892",
 19676 => x"C0C0C0F99082F882",
 19677 => x"C0C0C0F99082F8F8",
 19678 => x"C0C0C0F99082F880",
 19679 => x"C0C0C0F99082F890",
 19680 => x"C0C0C0F9908280C0",
 19681 => x"C0C0C0F9908280F9",
 19682 => x"C0C0C0F9908280A4",
 19683 => x"C0C0C0F9908280B0",
 19684 => x"C0C0C0F990828099",
 19685 => x"C0C0C0F990828092",
 19686 => x"C0C0C0F990828082",
 19687 => x"C0C0C0F9908280F8",
 19688 => x"C0C0C0F990828080",
 19689 => x"C0C0C0F990828090",
 19690 => x"C0C0C0F9908290C0",
 19691 => x"C0C0C0F9908290F9",
 19692 => x"C0C0C0F9908290A4",
 19693 => x"C0C0C0F9908290B0",
 19694 => x"C0C0C0F990829099",
 19695 => x"C0C0C0F990829092",
 19696 => x"C0C0C0F990829082",
 19697 => x"C0C0C0F9908290F8",
 19698 => x"C0C0C0F990829080",
 19699 => x"C0C0C0F990829090",
 19700 => x"C0C0C0F990F8C0C0",
 19701 => x"C0C0C0F990F8C0F9",
 19702 => x"C0C0C0F990F8C0A4",
 19703 => x"C0C0C0F990F8C0B0",
 19704 => x"C0C0C0F990F8C099",
 19705 => x"C0C0C0F990F8C092",
 19706 => x"C0C0C0F990F8C082",
 19707 => x"C0C0C0F990F8C0F8",
 19708 => x"C0C0C0F990F8C080",
 19709 => x"C0C0C0F990F8C090",
 19710 => x"C0C0C0F990F8F9C0",
 19711 => x"C0C0C0F990F8F9F9",
 19712 => x"C0C0C0F990F8F9A4",
 19713 => x"C0C0C0F990F8F9B0",
 19714 => x"C0C0C0F990F8F999",
 19715 => x"C0C0C0F990F8F992",
 19716 => x"C0C0C0F990F8F982",
 19717 => x"C0C0C0F990F8F9F8",
 19718 => x"C0C0C0F990F8F980",
 19719 => x"C0C0C0F990F8F990",
 19720 => x"C0C0C0F990F8A4C0",
 19721 => x"C0C0C0F990F8A4F9",
 19722 => x"C0C0C0F990F8A4A4",
 19723 => x"C0C0C0F990F8A4B0",
 19724 => x"C0C0C0F990F8A499",
 19725 => x"C0C0C0F990F8A492",
 19726 => x"C0C0C0F990F8A482",
 19727 => x"C0C0C0F990F8A4F8",
 19728 => x"C0C0C0F990F8A480",
 19729 => x"C0C0C0F990F8A490",
 19730 => x"C0C0C0F990F8B0C0",
 19731 => x"C0C0C0F990F8B0F9",
 19732 => x"C0C0C0F990F8B0A4",
 19733 => x"C0C0C0F990F8B0B0",
 19734 => x"C0C0C0F990F8B099",
 19735 => x"C0C0C0F990F8B092",
 19736 => x"C0C0C0F990F8B082",
 19737 => x"C0C0C0F990F8B0F8",
 19738 => x"C0C0C0F990F8B080",
 19739 => x"C0C0C0F990F8B090",
 19740 => x"C0C0C0F990F899C0",
 19741 => x"C0C0C0F990F899F9",
 19742 => x"C0C0C0F990F899A4",
 19743 => x"C0C0C0F990F899B0",
 19744 => x"C0C0C0F990F89999",
 19745 => x"C0C0C0F990F89992",
 19746 => x"C0C0C0F990F89982",
 19747 => x"C0C0C0F990F899F8",
 19748 => x"C0C0C0F990F89980",
 19749 => x"C0C0C0F990F89990",
 19750 => x"C0C0C0F990F892C0",
 19751 => x"C0C0C0F990F892F9",
 19752 => x"C0C0C0F990F892A4",
 19753 => x"C0C0C0F990F892B0",
 19754 => x"C0C0C0F990F89299",
 19755 => x"C0C0C0F990F89292",
 19756 => x"C0C0C0F990F89282",
 19757 => x"C0C0C0F990F892F8",
 19758 => x"C0C0C0F990F89280",
 19759 => x"C0C0C0F990F89290",
 19760 => x"C0C0C0F990F882C0",
 19761 => x"C0C0C0F990F882F9",
 19762 => x"C0C0C0F990F882A4",
 19763 => x"C0C0C0F990F882B0",
 19764 => x"C0C0C0F990F88299",
 19765 => x"C0C0C0F990F88292",
 19766 => x"C0C0C0F990F88282",
 19767 => x"C0C0C0F990F882F8",
 19768 => x"C0C0C0F990F88280",
 19769 => x"C0C0C0F990F88290",
 19770 => x"C0C0C0F990F8F8C0",
 19771 => x"C0C0C0F990F8F8F9",
 19772 => x"C0C0C0F990F8F8A4",
 19773 => x"C0C0C0F990F8F8B0",
 19774 => x"C0C0C0F990F8F899",
 19775 => x"C0C0C0F990F8F892",
 19776 => x"C0C0C0F990F8F882",
 19777 => x"C0C0C0F990F8F8F8",
 19778 => x"C0C0C0F990F8F880",
 19779 => x"C0C0C0F990F8F890",
 19780 => x"C0C0C0F990F880C0",
 19781 => x"C0C0C0F990F880F9",
 19782 => x"C0C0C0F990F880A4",
 19783 => x"C0C0C0F990F880B0",
 19784 => x"C0C0C0F990F88099",
 19785 => x"C0C0C0F990F88092",
 19786 => x"C0C0C0F990F88082",
 19787 => x"C0C0C0F990F880F8",
 19788 => x"C0C0C0F990F88080",
 19789 => x"C0C0C0F990F88090",
 19790 => x"C0C0C0F990F890C0",
 19791 => x"C0C0C0F990F890F9",
 19792 => x"C0C0C0F990F890A4",
 19793 => x"C0C0C0F990F890B0",
 19794 => x"C0C0C0F990F89099",
 19795 => x"C0C0C0F990F89092",
 19796 => x"C0C0C0F990F89082",
 19797 => x"C0C0C0F990F890F8",
 19798 => x"C0C0C0F990F89080",
 19799 => x"C0C0C0F990F89090",
 19800 => x"C0C0C0F99080C0C0",
 19801 => x"C0C0C0F99080C0F9",
 19802 => x"C0C0C0F99080C0A4",
 19803 => x"C0C0C0F99080C0B0",
 19804 => x"C0C0C0F99080C099",
 19805 => x"C0C0C0F99080C092",
 19806 => x"C0C0C0F99080C082",
 19807 => x"C0C0C0F99080C0F8",
 19808 => x"C0C0C0F99080C080",
 19809 => x"C0C0C0F99080C090",
 19810 => x"C0C0C0F99080F9C0",
 19811 => x"C0C0C0F99080F9F9",
 19812 => x"C0C0C0F99080F9A4",
 19813 => x"C0C0C0F99080F9B0",
 19814 => x"C0C0C0F99080F999",
 19815 => x"C0C0C0F99080F992",
 19816 => x"C0C0C0F99080F982",
 19817 => x"C0C0C0F99080F9F8",
 19818 => x"C0C0C0F99080F980",
 19819 => x"C0C0C0F99080F990",
 19820 => x"C0C0C0F99080A4C0",
 19821 => x"C0C0C0F99080A4F9",
 19822 => x"C0C0C0F99080A4A4",
 19823 => x"C0C0C0F99080A4B0",
 19824 => x"C0C0C0F99080A499",
 19825 => x"C0C0C0F99080A492",
 19826 => x"C0C0C0F99080A482",
 19827 => x"C0C0C0F99080A4F8",
 19828 => x"C0C0C0F99080A480",
 19829 => x"C0C0C0F99080A490",
 19830 => x"C0C0C0F99080B0C0",
 19831 => x"C0C0C0F99080B0F9",
 19832 => x"C0C0C0F99080B0A4",
 19833 => x"C0C0C0F99080B0B0",
 19834 => x"C0C0C0F99080B099",
 19835 => x"C0C0C0F99080B092",
 19836 => x"C0C0C0F99080B082",
 19837 => x"C0C0C0F99080B0F8",
 19838 => x"C0C0C0F99080B080",
 19839 => x"C0C0C0F99080B090",
 19840 => x"C0C0C0F9908099C0",
 19841 => x"C0C0C0F9908099F9",
 19842 => x"C0C0C0F9908099A4",
 19843 => x"C0C0C0F9908099B0",
 19844 => x"C0C0C0F990809999",
 19845 => x"C0C0C0F990809992",
 19846 => x"C0C0C0F990809982",
 19847 => x"C0C0C0F9908099F8",
 19848 => x"C0C0C0F990809980",
 19849 => x"C0C0C0F990809990",
 19850 => x"C0C0C0F9908092C0",
 19851 => x"C0C0C0F9908092F9",
 19852 => x"C0C0C0F9908092A4",
 19853 => x"C0C0C0F9908092B0",
 19854 => x"C0C0C0F990809299",
 19855 => x"C0C0C0F990809292",
 19856 => x"C0C0C0F990809282",
 19857 => x"C0C0C0F9908092F8",
 19858 => x"C0C0C0F990809280",
 19859 => x"C0C0C0F990809290",
 19860 => x"C0C0C0F9908082C0",
 19861 => x"C0C0C0F9908082F9",
 19862 => x"C0C0C0F9908082A4",
 19863 => x"C0C0C0F9908082B0",
 19864 => x"C0C0C0F990808299",
 19865 => x"C0C0C0F990808292",
 19866 => x"C0C0C0F990808282",
 19867 => x"C0C0C0F9908082F8",
 19868 => x"C0C0C0F990808280",
 19869 => x"C0C0C0F990808290",
 19870 => x"C0C0C0F99080F8C0",
 19871 => x"C0C0C0F99080F8F9",
 19872 => x"C0C0C0F99080F8A4",
 19873 => x"C0C0C0F99080F8B0",
 19874 => x"C0C0C0F99080F899",
 19875 => x"C0C0C0F99080F892",
 19876 => x"C0C0C0F99080F882",
 19877 => x"C0C0C0F99080F8F8",
 19878 => x"C0C0C0F99080F880",
 19879 => x"C0C0C0F99080F890",
 19880 => x"C0C0C0F9908080C0",
 19881 => x"C0C0C0F9908080F9",
 19882 => x"C0C0C0F9908080A4",
 19883 => x"C0C0C0F9908080B0",
 19884 => x"C0C0C0F990808099",
 19885 => x"C0C0C0F990808092",
 19886 => x"C0C0C0F990808082",
 19887 => x"C0C0C0F9908080F8",
 19888 => x"C0C0C0F990808080",
 19889 => x"C0C0C0F990808090",
 19890 => x"C0C0C0F9908090C0",
 19891 => x"C0C0C0F9908090F9",
 19892 => x"C0C0C0F9908090A4",
 19893 => x"C0C0C0F9908090B0",
 19894 => x"C0C0C0F990809099",
 19895 => x"C0C0C0F990809092",
 19896 => x"C0C0C0F990809082",
 19897 => x"C0C0C0F9908090F8",
 19898 => x"C0C0C0F990809080",
 19899 => x"C0C0C0F990809090",
 19900 => x"C0C0C0F99090C0C0",
 19901 => x"C0C0C0F99090C0F9",
 19902 => x"C0C0C0F99090C0A4",
 19903 => x"C0C0C0F99090C0B0",
 19904 => x"C0C0C0F99090C099",
 19905 => x"C0C0C0F99090C092",
 19906 => x"C0C0C0F99090C082",
 19907 => x"C0C0C0F99090C0F8",
 19908 => x"C0C0C0F99090C080",
 19909 => x"C0C0C0F99090C090",
 19910 => x"C0C0C0F99090F9C0",
 19911 => x"C0C0C0F99090F9F9",
 19912 => x"C0C0C0F99090F9A4",
 19913 => x"C0C0C0F99090F9B0",
 19914 => x"C0C0C0F99090F999",
 19915 => x"C0C0C0F99090F992",
 19916 => x"C0C0C0F99090F982",
 19917 => x"C0C0C0F99090F9F8",
 19918 => x"C0C0C0F99090F980",
 19919 => x"C0C0C0F99090F990",
 19920 => x"C0C0C0F99090A4C0",
 19921 => x"C0C0C0F99090A4F9",
 19922 => x"C0C0C0F99090A4A4",
 19923 => x"C0C0C0F99090A4B0",
 19924 => x"C0C0C0F99090A499",
 19925 => x"C0C0C0F99090A492",
 19926 => x"C0C0C0F99090A482",
 19927 => x"C0C0C0F99090A4F8",
 19928 => x"C0C0C0F99090A480",
 19929 => x"C0C0C0F99090A490",
 19930 => x"C0C0C0F99090B0C0",
 19931 => x"C0C0C0F99090B0F9",
 19932 => x"C0C0C0F99090B0A4",
 19933 => x"C0C0C0F99090B0B0",
 19934 => x"C0C0C0F99090B099",
 19935 => x"C0C0C0F99090B092",
 19936 => x"C0C0C0F99090B082",
 19937 => x"C0C0C0F99090B0F8",
 19938 => x"C0C0C0F99090B080",
 19939 => x"C0C0C0F99090B090",
 19940 => x"C0C0C0F9909099C0",
 19941 => x"C0C0C0F9909099F9",
 19942 => x"C0C0C0F9909099A4",
 19943 => x"C0C0C0F9909099B0",
 19944 => x"C0C0C0F990909999",
 19945 => x"C0C0C0F990909992",
 19946 => x"C0C0C0F990909982",
 19947 => x"C0C0C0F9909099F8",
 19948 => x"C0C0C0F990909980",
 19949 => x"C0C0C0F990909990",
 19950 => x"C0C0C0F9909092C0",
 19951 => x"C0C0C0F9909092F9",
 19952 => x"C0C0C0F9909092A4",
 19953 => x"C0C0C0F9909092B0",
 19954 => x"C0C0C0F990909299",
 19955 => x"C0C0C0F990909292",
 19956 => x"C0C0C0F990909282",
 19957 => x"C0C0C0F9909092F8",
 19958 => x"C0C0C0F990909280",
 19959 => x"C0C0C0F990909290",
 19960 => x"C0C0C0F9909082C0",
 19961 => x"C0C0C0F9909082F9",
 19962 => x"C0C0C0F9909082A4",
 19963 => x"C0C0C0F9909082B0",
 19964 => x"C0C0C0F990908299",
 19965 => x"C0C0C0F990908292",
 19966 => x"C0C0C0F990908282",
 19967 => x"C0C0C0F9909082F8",
 19968 => x"C0C0C0F990908280",
 19969 => x"C0C0C0F990908290",
 19970 => x"C0C0C0F99090F8C0",
 19971 => x"C0C0C0F99090F8F9",
 19972 => x"C0C0C0F99090F8A4",
 19973 => x"C0C0C0F99090F8B0",
 19974 => x"C0C0C0F99090F899",
 19975 => x"C0C0C0F99090F892",
 19976 => x"C0C0C0F99090F882",
 19977 => x"C0C0C0F99090F8F8",
 19978 => x"C0C0C0F99090F880",
 19979 => x"C0C0C0F99090F890",
 19980 => x"C0C0C0F9909080C0",
 19981 => x"C0C0C0F9909080F9",
 19982 => x"C0C0C0F9909080A4",
 19983 => x"C0C0C0F9909080B0",
 19984 => x"C0C0C0F990908099",
 19985 => x"C0C0C0F990908092",
 19986 => x"C0C0C0F990908082",
 19987 => x"C0C0C0F9909080F8",
 19988 => x"C0C0C0F990908080",
 19989 => x"C0C0C0F990908090",
 19990 => x"C0C0C0F9909090C0",
 19991 => x"C0C0C0F9909090F9",
 19992 => x"C0C0C0F9909090A4",
 19993 => x"C0C0C0F9909090B0",
 19994 => x"C0C0C0F990909099",
 19995 => x"C0C0C0F990909092",
 19996 => x"C0C0C0F990909082",
 19997 => x"C0C0C0F9909090F8",
 19998 => x"C0C0C0F990909080",
 19999 => x"C0C0C0F990909090",
 20000 => x"C0C0C0A4C0C0C0C0",
 20001 => x"C0C0C0A4C0C0C0F9",
 20002 => x"C0C0C0A4C0C0C0A4",
 20003 => x"C0C0C0A4C0C0C0B0",
 20004 => x"C0C0C0A4C0C0C099",
 20005 => x"C0C0C0A4C0C0C092",
 20006 => x"C0C0C0A4C0C0C082",
 20007 => x"C0C0C0A4C0C0C0F8",
 20008 => x"C0C0C0A4C0C0C080",
 20009 => x"C0C0C0A4C0C0C090",
 20010 => x"C0C0C0A4C0C0F9C0",
 20011 => x"C0C0C0A4C0C0F9F9",
 20012 => x"C0C0C0A4C0C0F9A4",
 20013 => x"C0C0C0A4C0C0F9B0",
 20014 => x"C0C0C0A4C0C0F999",
 20015 => x"C0C0C0A4C0C0F992",
 20016 => x"C0C0C0A4C0C0F982",
 20017 => x"C0C0C0A4C0C0F9F8",
 20018 => x"C0C0C0A4C0C0F980",
 20019 => x"C0C0C0A4C0C0F990",
 20020 => x"C0C0C0A4C0C0A4C0",
 20021 => x"C0C0C0A4C0C0A4F9",
 20022 => x"C0C0C0A4C0C0A4A4",
 20023 => x"C0C0C0A4C0C0A4B0",
 20024 => x"C0C0C0A4C0C0A499",
 20025 => x"C0C0C0A4C0C0A492",
 20026 => x"C0C0C0A4C0C0A482",
 20027 => x"C0C0C0A4C0C0A4F8",
 20028 => x"C0C0C0A4C0C0A480",
 20029 => x"C0C0C0A4C0C0A490",
 20030 => x"C0C0C0A4C0C0B0C0",
 20031 => x"C0C0C0A4C0C0B0F9",
 20032 => x"C0C0C0A4C0C0B0A4",
 20033 => x"C0C0C0A4C0C0B0B0",
 20034 => x"C0C0C0A4C0C0B099",
 20035 => x"C0C0C0A4C0C0B092",
 20036 => x"C0C0C0A4C0C0B082",
 20037 => x"C0C0C0A4C0C0B0F8",
 20038 => x"C0C0C0A4C0C0B080",
 20039 => x"C0C0C0A4C0C0B090",
 20040 => x"C0C0C0A4C0C099C0",
 20041 => x"C0C0C0A4C0C099F9",
 20042 => x"C0C0C0A4C0C099A4",
 20043 => x"C0C0C0A4C0C099B0",
 20044 => x"C0C0C0A4C0C09999",
 20045 => x"C0C0C0A4C0C09992",
 20046 => x"C0C0C0A4C0C09982",
 20047 => x"C0C0C0A4C0C099F8",
 20048 => x"C0C0C0A4C0C09980",
 20049 => x"C0C0C0A4C0C09990",
 20050 => x"C0C0C0A4C0C092C0",
 20051 => x"C0C0C0A4C0C092F9",
 20052 => x"C0C0C0A4C0C092A4",
 20053 => x"C0C0C0A4C0C092B0",
 20054 => x"C0C0C0A4C0C09299",
 20055 => x"C0C0C0A4C0C09292",
 20056 => x"C0C0C0A4C0C09282",
 20057 => x"C0C0C0A4C0C092F8",
 20058 => x"C0C0C0A4C0C09280",
 20059 => x"C0C0C0A4C0C09290",
 20060 => x"C0C0C0A4C0C082C0",
 20061 => x"C0C0C0A4C0C082F9",
 20062 => x"C0C0C0A4C0C082A4",
 20063 => x"C0C0C0A4C0C082B0",
 20064 => x"C0C0C0A4C0C08299",
 20065 => x"C0C0C0A4C0C08292",
 20066 => x"C0C0C0A4C0C08282",
 20067 => x"C0C0C0A4C0C082F8",
 20068 => x"C0C0C0A4C0C08280",
 20069 => x"C0C0C0A4C0C08290",
 20070 => x"C0C0C0A4C0C0F8C0",
 20071 => x"C0C0C0A4C0C0F8F9",
 20072 => x"C0C0C0A4C0C0F8A4",
 20073 => x"C0C0C0A4C0C0F8B0",
 20074 => x"C0C0C0A4C0C0F899",
 20075 => x"C0C0C0A4C0C0F892",
 20076 => x"C0C0C0A4C0C0F882",
 20077 => x"C0C0C0A4C0C0F8F8",
 20078 => x"C0C0C0A4C0C0F880",
 20079 => x"C0C0C0A4C0C0F890",
 20080 => x"C0C0C0A4C0C080C0",
 20081 => x"C0C0C0A4C0C080F9",
 20082 => x"C0C0C0A4C0C080A4",
 20083 => x"C0C0C0A4C0C080B0",
 20084 => x"C0C0C0A4C0C08099",
 20085 => x"C0C0C0A4C0C08092",
 20086 => x"C0C0C0A4C0C08082",
 20087 => x"C0C0C0A4C0C080F8",
 20088 => x"C0C0C0A4C0C08080",
 20089 => x"C0C0C0A4C0C08090",
 20090 => x"C0C0C0A4C0C090C0",
 20091 => x"C0C0C0A4C0C090F9",
 20092 => x"C0C0C0A4C0C090A4",
 20093 => x"C0C0C0A4C0C090B0",
 20094 => x"C0C0C0A4C0C09099",
 20095 => x"C0C0C0A4C0C09092",
 20096 => x"C0C0C0A4C0C09082",
 20097 => x"C0C0C0A4C0C090F8",
 20098 => x"C0C0C0A4C0C09080",
 20099 => x"C0C0C0A4C0C09090",
 20100 => x"C0C0C0A4C0F9C0C0",
 20101 => x"C0C0C0A4C0F9C0F9",
 20102 => x"C0C0C0A4C0F9C0A4",
 20103 => x"C0C0C0A4C0F9C0B0",
 20104 => x"C0C0C0A4C0F9C099",
 20105 => x"C0C0C0A4C0F9C092",
 20106 => x"C0C0C0A4C0F9C082",
 20107 => x"C0C0C0A4C0F9C0F8",
 20108 => x"C0C0C0A4C0F9C080",
 20109 => x"C0C0C0A4C0F9C090",
 20110 => x"C0C0C0A4C0F9F9C0",
 20111 => x"C0C0C0A4C0F9F9F9",
 20112 => x"C0C0C0A4C0F9F9A4",
 20113 => x"C0C0C0A4C0F9F9B0",
 20114 => x"C0C0C0A4C0F9F999",
 20115 => x"C0C0C0A4C0F9F992",
 20116 => x"C0C0C0A4C0F9F982",
 20117 => x"C0C0C0A4C0F9F9F8",
 20118 => x"C0C0C0A4C0F9F980",
 20119 => x"C0C0C0A4C0F9F990",
 20120 => x"C0C0C0A4C0F9A4C0",
 20121 => x"C0C0C0A4C0F9A4F9",
 20122 => x"C0C0C0A4C0F9A4A4",
 20123 => x"C0C0C0A4C0F9A4B0",
 20124 => x"C0C0C0A4C0F9A499",
 20125 => x"C0C0C0A4C0F9A492",
 20126 => x"C0C0C0A4C0F9A482",
 20127 => x"C0C0C0A4C0F9A4F8",
 20128 => x"C0C0C0A4C0F9A480",
 20129 => x"C0C0C0A4C0F9A490",
 20130 => x"C0C0C0A4C0F9B0C0",
 20131 => x"C0C0C0A4C0F9B0F9",
 20132 => x"C0C0C0A4C0F9B0A4",
 20133 => x"C0C0C0A4C0F9B0B0",
 20134 => x"C0C0C0A4C0F9B099",
 20135 => x"C0C0C0A4C0F9B092",
 20136 => x"C0C0C0A4C0F9B082",
 20137 => x"C0C0C0A4C0F9B0F8",
 20138 => x"C0C0C0A4C0F9B080",
 20139 => x"C0C0C0A4C0F9B090",
 20140 => x"C0C0C0A4C0F999C0",
 20141 => x"C0C0C0A4C0F999F9",
 20142 => x"C0C0C0A4C0F999A4",
 20143 => x"C0C0C0A4C0F999B0",
 20144 => x"C0C0C0A4C0F99999",
 20145 => x"C0C0C0A4C0F99992",
 20146 => x"C0C0C0A4C0F99982",
 20147 => x"C0C0C0A4C0F999F8",
 20148 => x"C0C0C0A4C0F99980",
 20149 => x"C0C0C0A4C0F99990",
 20150 => x"C0C0C0A4C0F992C0",
 20151 => x"C0C0C0A4C0F992F9",
 20152 => x"C0C0C0A4C0F992A4",
 20153 => x"C0C0C0A4C0F992B0",
 20154 => x"C0C0C0A4C0F99299",
 20155 => x"C0C0C0A4C0F99292",
 20156 => x"C0C0C0A4C0F99282",
 20157 => x"C0C0C0A4C0F992F8",
 20158 => x"C0C0C0A4C0F99280",
 20159 => x"C0C0C0A4C0F99290",
 20160 => x"C0C0C0A4C0F982C0",
 20161 => x"C0C0C0A4C0F982F9",
 20162 => x"C0C0C0A4C0F982A4",
 20163 => x"C0C0C0A4C0F982B0",
 20164 => x"C0C0C0A4C0F98299",
 20165 => x"C0C0C0A4C0F98292",
 20166 => x"C0C0C0A4C0F98282",
 20167 => x"C0C0C0A4C0F982F8",
 20168 => x"C0C0C0A4C0F98280",
 20169 => x"C0C0C0A4C0F98290",
 20170 => x"C0C0C0A4C0F9F8C0",
 20171 => x"C0C0C0A4C0F9F8F9",
 20172 => x"C0C0C0A4C0F9F8A4",
 20173 => x"C0C0C0A4C0F9F8B0",
 20174 => x"C0C0C0A4C0F9F899",
 20175 => x"C0C0C0A4C0F9F892",
 20176 => x"C0C0C0A4C0F9F882",
 20177 => x"C0C0C0A4C0F9F8F8",
 20178 => x"C0C0C0A4C0F9F880",
 20179 => x"C0C0C0A4C0F9F890",
 20180 => x"C0C0C0A4C0F980C0",
 20181 => x"C0C0C0A4C0F980F9",
 20182 => x"C0C0C0A4C0F980A4",
 20183 => x"C0C0C0A4C0F980B0",
 20184 => x"C0C0C0A4C0F98099",
 20185 => x"C0C0C0A4C0F98092",
 20186 => x"C0C0C0A4C0F98082",
 20187 => x"C0C0C0A4C0F980F8",
 20188 => x"C0C0C0A4C0F98080",
 20189 => x"C0C0C0A4C0F98090",
 20190 => x"C0C0C0A4C0F990C0",
 20191 => x"C0C0C0A4C0F990F9",
 20192 => x"C0C0C0A4C0F990A4",
 20193 => x"C0C0C0A4C0F990B0",
 20194 => x"C0C0C0A4C0F99099",
 20195 => x"C0C0C0A4C0F99092",
 20196 => x"C0C0C0A4C0F99082",
 20197 => x"C0C0C0A4C0F990F8",
 20198 => x"C0C0C0A4C0F99080",
 20199 => x"C0C0C0A4C0F99090",
 20200 => x"C0C0C0A4C0A4C0C0",
 20201 => x"C0C0C0A4C0A4C0F9",
 20202 => x"C0C0C0A4C0A4C0A4",
 20203 => x"C0C0C0A4C0A4C0B0",
 20204 => x"C0C0C0A4C0A4C099",
 20205 => x"C0C0C0A4C0A4C092",
 20206 => x"C0C0C0A4C0A4C082",
 20207 => x"C0C0C0A4C0A4C0F8",
 20208 => x"C0C0C0A4C0A4C080",
 20209 => x"C0C0C0A4C0A4C090",
 20210 => x"C0C0C0A4C0A4F9C0",
 20211 => x"C0C0C0A4C0A4F9F9",
 20212 => x"C0C0C0A4C0A4F9A4",
 20213 => x"C0C0C0A4C0A4F9B0",
 20214 => x"C0C0C0A4C0A4F999",
 20215 => x"C0C0C0A4C0A4F992",
 20216 => x"C0C0C0A4C0A4F982",
 20217 => x"C0C0C0A4C0A4F9F8",
 20218 => x"C0C0C0A4C0A4F980",
 20219 => x"C0C0C0A4C0A4F990",
 20220 => x"C0C0C0A4C0A4A4C0",
 20221 => x"C0C0C0A4C0A4A4F9",
 20222 => x"C0C0C0A4C0A4A4A4",
 20223 => x"C0C0C0A4C0A4A4B0",
 20224 => x"C0C0C0A4C0A4A499",
 20225 => x"C0C0C0A4C0A4A492",
 20226 => x"C0C0C0A4C0A4A482",
 20227 => x"C0C0C0A4C0A4A4F8",
 20228 => x"C0C0C0A4C0A4A480",
 20229 => x"C0C0C0A4C0A4A490",
 20230 => x"C0C0C0A4C0A4B0C0",
 20231 => x"C0C0C0A4C0A4B0F9",
 20232 => x"C0C0C0A4C0A4B0A4",
 20233 => x"C0C0C0A4C0A4B0B0",
 20234 => x"C0C0C0A4C0A4B099",
 20235 => x"C0C0C0A4C0A4B092",
 20236 => x"C0C0C0A4C0A4B082",
 20237 => x"C0C0C0A4C0A4B0F8",
 20238 => x"C0C0C0A4C0A4B080",
 20239 => x"C0C0C0A4C0A4B090",
 20240 => x"C0C0C0A4C0A499C0",
 20241 => x"C0C0C0A4C0A499F9",
 20242 => x"C0C0C0A4C0A499A4",
 20243 => x"C0C0C0A4C0A499B0",
 20244 => x"C0C0C0A4C0A49999",
 20245 => x"C0C0C0A4C0A49992",
 20246 => x"C0C0C0A4C0A49982",
 20247 => x"C0C0C0A4C0A499F8",
 20248 => x"C0C0C0A4C0A49980",
 20249 => x"C0C0C0A4C0A49990",
 20250 => x"C0C0C0A4C0A492C0",
 20251 => x"C0C0C0A4C0A492F9",
 20252 => x"C0C0C0A4C0A492A4",
 20253 => x"C0C0C0A4C0A492B0",
 20254 => x"C0C0C0A4C0A49299",
 20255 => x"C0C0C0A4C0A49292",
 20256 => x"C0C0C0A4C0A49282",
 20257 => x"C0C0C0A4C0A492F8",
 20258 => x"C0C0C0A4C0A49280",
 20259 => x"C0C0C0A4C0A49290",
 20260 => x"C0C0C0A4C0A482C0",
 20261 => x"C0C0C0A4C0A482F9",
 20262 => x"C0C0C0A4C0A482A4",
 20263 => x"C0C0C0A4C0A482B0",
 20264 => x"C0C0C0A4C0A48299",
 20265 => x"C0C0C0A4C0A48292",
 20266 => x"C0C0C0A4C0A48282",
 20267 => x"C0C0C0A4C0A482F8",
 20268 => x"C0C0C0A4C0A48280",
 20269 => x"C0C0C0A4C0A48290",
 20270 => x"C0C0C0A4C0A4F8C0",
 20271 => x"C0C0C0A4C0A4F8F9",
 20272 => x"C0C0C0A4C0A4F8A4",
 20273 => x"C0C0C0A4C0A4F8B0",
 20274 => x"C0C0C0A4C0A4F899",
 20275 => x"C0C0C0A4C0A4F892",
 20276 => x"C0C0C0A4C0A4F882",
 20277 => x"C0C0C0A4C0A4F8F8",
 20278 => x"C0C0C0A4C0A4F880",
 20279 => x"C0C0C0A4C0A4F890",
 20280 => x"C0C0C0A4C0A480C0",
 20281 => x"C0C0C0A4C0A480F9",
 20282 => x"C0C0C0A4C0A480A4",
 20283 => x"C0C0C0A4C0A480B0",
 20284 => x"C0C0C0A4C0A48099",
 20285 => x"C0C0C0A4C0A48092",
 20286 => x"C0C0C0A4C0A48082",
 20287 => x"C0C0C0A4C0A480F8",
 20288 => x"C0C0C0A4C0A48080",
 20289 => x"C0C0C0A4C0A48090",
 20290 => x"C0C0C0A4C0A490C0",
 20291 => x"C0C0C0A4C0A490F9",
 20292 => x"C0C0C0A4C0A490A4",
 20293 => x"C0C0C0A4C0A490B0",
 20294 => x"C0C0C0A4C0A49099",
 20295 => x"C0C0C0A4C0A49092",
 20296 => x"C0C0C0A4C0A49082",
 20297 => x"C0C0C0A4C0A490F8",
 20298 => x"C0C0C0A4C0A49080",
 20299 => x"C0C0C0A4C0A49090",
 20300 => x"C0C0C0A4C0B0C0C0",
 20301 => x"C0C0C0A4C0B0C0F9",
 20302 => x"C0C0C0A4C0B0C0A4",
 20303 => x"C0C0C0A4C0B0C0B0",
 20304 => x"C0C0C0A4C0B0C099",
 20305 => x"C0C0C0A4C0B0C092",
 20306 => x"C0C0C0A4C0B0C082",
 20307 => x"C0C0C0A4C0B0C0F8",
 20308 => x"C0C0C0A4C0B0C080",
 20309 => x"C0C0C0A4C0B0C090",
 20310 => x"C0C0C0A4C0B0F9C0",
 20311 => x"C0C0C0A4C0B0F9F9",
 20312 => x"C0C0C0A4C0B0F9A4",
 20313 => x"C0C0C0A4C0B0F9B0",
 20314 => x"C0C0C0A4C0B0F999",
 20315 => x"C0C0C0A4C0B0F992",
 20316 => x"C0C0C0A4C0B0F982",
 20317 => x"C0C0C0A4C0B0F9F8",
 20318 => x"C0C0C0A4C0B0F980",
 20319 => x"C0C0C0A4C0B0F990",
 20320 => x"C0C0C0A4C0B0A4C0",
 20321 => x"C0C0C0A4C0B0A4F9",
 20322 => x"C0C0C0A4C0B0A4A4",
 20323 => x"C0C0C0A4C0B0A4B0",
 20324 => x"C0C0C0A4C0B0A499",
 20325 => x"C0C0C0A4C0B0A492",
 20326 => x"C0C0C0A4C0B0A482",
 20327 => x"C0C0C0A4C0B0A4F8",
 20328 => x"C0C0C0A4C0B0A480",
 20329 => x"C0C0C0A4C0B0A490",
 20330 => x"C0C0C0A4C0B0B0C0",
 20331 => x"C0C0C0A4C0B0B0F9",
 20332 => x"C0C0C0A4C0B0B0A4",
 20333 => x"C0C0C0A4C0B0B0B0",
 20334 => x"C0C0C0A4C0B0B099",
 20335 => x"C0C0C0A4C0B0B092",
 20336 => x"C0C0C0A4C0B0B082",
 20337 => x"C0C0C0A4C0B0B0F8",
 20338 => x"C0C0C0A4C0B0B080",
 20339 => x"C0C0C0A4C0B0B090",
 20340 => x"C0C0C0A4C0B099C0",
 20341 => x"C0C0C0A4C0B099F9",
 20342 => x"C0C0C0A4C0B099A4",
 20343 => x"C0C0C0A4C0B099B0",
 20344 => x"C0C0C0A4C0B09999",
 20345 => x"C0C0C0A4C0B09992",
 20346 => x"C0C0C0A4C0B09982",
 20347 => x"C0C0C0A4C0B099F8",
 20348 => x"C0C0C0A4C0B09980",
 20349 => x"C0C0C0A4C0B09990",
 20350 => x"C0C0C0A4C0B092C0",
 20351 => x"C0C0C0A4C0B092F9",
 20352 => x"C0C0C0A4C0B092A4",
 20353 => x"C0C0C0A4C0B092B0",
 20354 => x"C0C0C0A4C0B09299",
 20355 => x"C0C0C0A4C0B09292",
 20356 => x"C0C0C0A4C0B09282",
 20357 => x"C0C0C0A4C0B092F8",
 20358 => x"C0C0C0A4C0B09280",
 20359 => x"C0C0C0A4C0B09290",
 20360 => x"C0C0C0A4C0B082C0",
 20361 => x"C0C0C0A4C0B082F9",
 20362 => x"C0C0C0A4C0B082A4",
 20363 => x"C0C0C0A4C0B082B0",
 20364 => x"C0C0C0A4C0B08299",
 20365 => x"C0C0C0A4C0B08292",
 20366 => x"C0C0C0A4C0B08282",
 20367 => x"C0C0C0A4C0B082F8",
 20368 => x"C0C0C0A4C0B08280",
 20369 => x"C0C0C0A4C0B08290",
 20370 => x"C0C0C0A4C0B0F8C0",
 20371 => x"C0C0C0A4C0B0F8F9",
 20372 => x"C0C0C0A4C0B0F8A4",
 20373 => x"C0C0C0A4C0B0F8B0",
 20374 => x"C0C0C0A4C0B0F899",
 20375 => x"C0C0C0A4C0B0F892",
 20376 => x"C0C0C0A4C0B0F882",
 20377 => x"C0C0C0A4C0B0F8F8",
 20378 => x"C0C0C0A4C0B0F880",
 20379 => x"C0C0C0A4C0B0F890",
 20380 => x"C0C0C0A4C0B080C0",
 20381 => x"C0C0C0A4C0B080F9",
 20382 => x"C0C0C0A4C0B080A4",
 20383 => x"C0C0C0A4C0B080B0",
 20384 => x"C0C0C0A4C0B08099",
 20385 => x"C0C0C0A4C0B08092",
 20386 => x"C0C0C0A4C0B08082",
 20387 => x"C0C0C0A4C0B080F8",
 20388 => x"C0C0C0A4C0B08080",
 20389 => x"C0C0C0A4C0B08090",
 20390 => x"C0C0C0A4C0B090C0",
 20391 => x"C0C0C0A4C0B090F9",
 20392 => x"C0C0C0A4C0B090A4",
 20393 => x"C0C0C0A4C0B090B0",
 20394 => x"C0C0C0A4C0B09099",
 20395 => x"C0C0C0A4C0B09092",
 20396 => x"C0C0C0A4C0B09082",
 20397 => x"C0C0C0A4C0B090F8",
 20398 => x"C0C0C0A4C0B09080",
 20399 => x"C0C0C0A4C0B09090",
 20400 => x"C0C0C0A4C099C0C0",
 20401 => x"C0C0C0A4C099C0F9",
 20402 => x"C0C0C0A4C099C0A4",
 20403 => x"C0C0C0A4C099C0B0",
 20404 => x"C0C0C0A4C099C099",
 20405 => x"C0C0C0A4C099C092",
 20406 => x"C0C0C0A4C099C082",
 20407 => x"C0C0C0A4C099C0F8",
 20408 => x"C0C0C0A4C099C080",
 20409 => x"C0C0C0A4C099C090",
 20410 => x"C0C0C0A4C099F9C0",
 20411 => x"C0C0C0A4C099F9F9",
 20412 => x"C0C0C0A4C099F9A4",
 20413 => x"C0C0C0A4C099F9B0",
 20414 => x"C0C0C0A4C099F999",
 20415 => x"C0C0C0A4C099F992",
 20416 => x"C0C0C0A4C099F982",
 20417 => x"C0C0C0A4C099F9F8",
 20418 => x"C0C0C0A4C099F980",
 20419 => x"C0C0C0A4C099F990",
 20420 => x"C0C0C0A4C099A4C0",
 20421 => x"C0C0C0A4C099A4F9",
 20422 => x"C0C0C0A4C099A4A4",
 20423 => x"C0C0C0A4C099A4B0",
 20424 => x"C0C0C0A4C099A499",
 20425 => x"C0C0C0A4C099A492",
 20426 => x"C0C0C0A4C099A482",
 20427 => x"C0C0C0A4C099A4F8",
 20428 => x"C0C0C0A4C099A480",
 20429 => x"C0C0C0A4C099A490",
 20430 => x"C0C0C0A4C099B0C0",
 20431 => x"C0C0C0A4C099B0F9",
 20432 => x"C0C0C0A4C099B0A4",
 20433 => x"C0C0C0A4C099B0B0",
 20434 => x"C0C0C0A4C099B099",
 20435 => x"C0C0C0A4C099B092",
 20436 => x"C0C0C0A4C099B082",
 20437 => x"C0C0C0A4C099B0F8",
 20438 => x"C0C0C0A4C099B080",
 20439 => x"C0C0C0A4C099B090",
 20440 => x"C0C0C0A4C09999C0",
 20441 => x"C0C0C0A4C09999F9",
 20442 => x"C0C0C0A4C09999A4",
 20443 => x"C0C0C0A4C09999B0",
 20444 => x"C0C0C0A4C0999999",
 20445 => x"C0C0C0A4C0999992",
 20446 => x"C0C0C0A4C0999982",
 20447 => x"C0C0C0A4C09999F8",
 20448 => x"C0C0C0A4C0999980",
 20449 => x"C0C0C0A4C0999990",
 20450 => x"C0C0C0A4C09992C0",
 20451 => x"C0C0C0A4C09992F9",
 20452 => x"C0C0C0A4C09992A4",
 20453 => x"C0C0C0A4C09992B0",
 20454 => x"C0C0C0A4C0999299",
 20455 => x"C0C0C0A4C0999292",
 20456 => x"C0C0C0A4C0999282",
 20457 => x"C0C0C0A4C09992F8",
 20458 => x"C0C0C0A4C0999280",
 20459 => x"C0C0C0A4C0999290",
 20460 => x"C0C0C0A4C09982C0",
 20461 => x"C0C0C0A4C09982F9",
 20462 => x"C0C0C0A4C09982A4",
 20463 => x"C0C0C0A4C09982B0",
 20464 => x"C0C0C0A4C0998299",
 20465 => x"C0C0C0A4C0998292",
 20466 => x"C0C0C0A4C0998282",
 20467 => x"C0C0C0A4C09982F8",
 20468 => x"C0C0C0A4C0998280",
 20469 => x"C0C0C0A4C0998290",
 20470 => x"C0C0C0A4C099F8C0",
 20471 => x"C0C0C0A4C099F8F9",
 20472 => x"C0C0C0A4C099F8A4",
 20473 => x"C0C0C0A4C099F8B0",
 20474 => x"C0C0C0A4C099F899",
 20475 => x"C0C0C0A4C099F892",
 20476 => x"C0C0C0A4C099F882",
 20477 => x"C0C0C0A4C099F8F8",
 20478 => x"C0C0C0A4C099F880",
 20479 => x"C0C0C0A4C099F890",
 20480 => x"C0C0C0A4C09980C0",
 20481 => x"C0C0C0A4C09980F9",
 20482 => x"C0C0C0A4C09980A4",
 20483 => x"C0C0C0A4C09980B0",
 20484 => x"C0C0C0A4C0998099",
 20485 => x"C0C0C0A4C0998092",
 20486 => x"C0C0C0A4C0998082",
 20487 => x"C0C0C0A4C09980F8",
 20488 => x"C0C0C0A4C0998080",
 20489 => x"C0C0C0A4C0998090",
 20490 => x"C0C0C0A4C09990C0",
 20491 => x"C0C0C0A4C09990F9",
 20492 => x"C0C0C0A4C09990A4",
 20493 => x"C0C0C0A4C09990B0",
 20494 => x"C0C0C0A4C0999099",
 20495 => x"C0C0C0A4C0999092",
 20496 => x"C0C0C0A4C0999082",
 20497 => x"C0C0C0A4C09990F8",
 20498 => x"C0C0C0A4C0999080",
 20499 => x"C0C0C0A4C0999090",
 20500 => x"C0C0C0A4C092C0C0",
 20501 => x"C0C0C0A4C092C0F9",
 20502 => x"C0C0C0A4C092C0A4",
 20503 => x"C0C0C0A4C092C0B0",
 20504 => x"C0C0C0A4C092C099",
 20505 => x"C0C0C0A4C092C092",
 20506 => x"C0C0C0A4C092C082",
 20507 => x"C0C0C0A4C092C0F8",
 20508 => x"C0C0C0A4C092C080",
 20509 => x"C0C0C0A4C092C090",
 20510 => x"C0C0C0A4C092F9C0",
 20511 => x"C0C0C0A4C092F9F9",
 20512 => x"C0C0C0A4C092F9A4",
 20513 => x"C0C0C0A4C092F9B0",
 20514 => x"C0C0C0A4C092F999",
 20515 => x"C0C0C0A4C092F992",
 20516 => x"C0C0C0A4C092F982",
 20517 => x"C0C0C0A4C092F9F8",
 20518 => x"C0C0C0A4C092F980",
 20519 => x"C0C0C0A4C092F990",
 20520 => x"C0C0C0A4C092A4C0",
 20521 => x"C0C0C0A4C092A4F9",
 20522 => x"C0C0C0A4C092A4A4",
 20523 => x"C0C0C0A4C092A4B0",
 20524 => x"C0C0C0A4C092A499",
 20525 => x"C0C0C0A4C092A492",
 20526 => x"C0C0C0A4C092A482",
 20527 => x"C0C0C0A4C092A4F8",
 20528 => x"C0C0C0A4C092A480",
 20529 => x"C0C0C0A4C092A490",
 20530 => x"C0C0C0A4C092B0C0",
 20531 => x"C0C0C0A4C092B0F9",
 20532 => x"C0C0C0A4C092B0A4",
 20533 => x"C0C0C0A4C092B0B0",
 20534 => x"C0C0C0A4C092B099",
 20535 => x"C0C0C0A4C092B092",
 20536 => x"C0C0C0A4C092B082",
 20537 => x"C0C0C0A4C092B0F8",
 20538 => x"C0C0C0A4C092B080",
 20539 => x"C0C0C0A4C092B090",
 20540 => x"C0C0C0A4C09299C0",
 20541 => x"C0C0C0A4C09299F9",
 20542 => x"C0C0C0A4C09299A4",
 20543 => x"C0C0C0A4C09299B0",
 20544 => x"C0C0C0A4C0929999",
 20545 => x"C0C0C0A4C0929992",
 20546 => x"C0C0C0A4C0929982",
 20547 => x"C0C0C0A4C09299F8",
 20548 => x"C0C0C0A4C0929980",
 20549 => x"C0C0C0A4C0929990",
 20550 => x"C0C0C0A4C09292C0",
 20551 => x"C0C0C0A4C09292F9",
 20552 => x"C0C0C0A4C09292A4",
 20553 => x"C0C0C0A4C09292B0",
 20554 => x"C0C0C0A4C0929299",
 20555 => x"C0C0C0A4C0929292",
 20556 => x"C0C0C0A4C0929282",
 20557 => x"C0C0C0A4C09292F8",
 20558 => x"C0C0C0A4C0929280",
 20559 => x"C0C0C0A4C0929290",
 20560 => x"C0C0C0A4C09282C0",
 20561 => x"C0C0C0A4C09282F9",
 20562 => x"C0C0C0A4C09282A4",
 20563 => x"C0C0C0A4C09282B0",
 20564 => x"C0C0C0A4C0928299",
 20565 => x"C0C0C0A4C0928292",
 20566 => x"C0C0C0A4C0928282",
 20567 => x"C0C0C0A4C09282F8",
 20568 => x"C0C0C0A4C0928280",
 20569 => x"C0C0C0A4C0928290",
 20570 => x"C0C0C0A4C092F8C0",
 20571 => x"C0C0C0A4C092F8F9",
 20572 => x"C0C0C0A4C092F8A4",
 20573 => x"C0C0C0A4C092F8B0",
 20574 => x"C0C0C0A4C092F899",
 20575 => x"C0C0C0A4C092F892",
 20576 => x"C0C0C0A4C092F882",
 20577 => x"C0C0C0A4C092F8F8",
 20578 => x"C0C0C0A4C092F880",
 20579 => x"C0C0C0A4C092F890",
 20580 => x"C0C0C0A4C09280C0",
 20581 => x"C0C0C0A4C09280F9",
 20582 => x"C0C0C0A4C09280A4",
 20583 => x"C0C0C0A4C09280B0",
 20584 => x"C0C0C0A4C0928099",
 20585 => x"C0C0C0A4C0928092",
 20586 => x"C0C0C0A4C0928082",
 20587 => x"C0C0C0A4C09280F8",
 20588 => x"C0C0C0A4C0928080",
 20589 => x"C0C0C0A4C0928090",
 20590 => x"C0C0C0A4C09290C0",
 20591 => x"C0C0C0A4C09290F9",
 20592 => x"C0C0C0A4C09290A4",
 20593 => x"C0C0C0A4C09290B0",
 20594 => x"C0C0C0A4C0929099",
 20595 => x"C0C0C0A4C0929092",
 20596 => x"C0C0C0A4C0929082",
 20597 => x"C0C0C0A4C09290F8",
 20598 => x"C0C0C0A4C0929080",
 20599 => x"C0C0C0A4C0929090",
 20600 => x"C0C0C0A4C082C0C0",
 20601 => x"C0C0C0A4C082C0F9",
 20602 => x"C0C0C0A4C082C0A4",
 20603 => x"C0C0C0A4C082C0B0",
 20604 => x"C0C0C0A4C082C099",
 20605 => x"C0C0C0A4C082C092",
 20606 => x"C0C0C0A4C082C082",
 20607 => x"C0C0C0A4C082C0F8",
 20608 => x"C0C0C0A4C082C080",
 20609 => x"C0C0C0A4C082C090",
 20610 => x"C0C0C0A4C082F9C0",
 20611 => x"C0C0C0A4C082F9F9",
 20612 => x"C0C0C0A4C082F9A4",
 20613 => x"C0C0C0A4C082F9B0",
 20614 => x"C0C0C0A4C082F999",
 20615 => x"C0C0C0A4C082F992",
 20616 => x"C0C0C0A4C082F982",
 20617 => x"C0C0C0A4C082F9F8",
 20618 => x"C0C0C0A4C082F980",
 20619 => x"C0C0C0A4C082F990",
 20620 => x"C0C0C0A4C082A4C0",
 20621 => x"C0C0C0A4C082A4F9",
 20622 => x"C0C0C0A4C082A4A4",
 20623 => x"C0C0C0A4C082A4B0",
 20624 => x"C0C0C0A4C082A499",
 20625 => x"C0C0C0A4C082A492",
 20626 => x"C0C0C0A4C082A482",
 20627 => x"C0C0C0A4C082A4F8",
 20628 => x"C0C0C0A4C082A480",
 20629 => x"C0C0C0A4C082A490",
 20630 => x"C0C0C0A4C082B0C0",
 20631 => x"C0C0C0A4C082B0F9",
 20632 => x"C0C0C0A4C082B0A4",
 20633 => x"C0C0C0A4C082B0B0",
 20634 => x"C0C0C0A4C082B099",
 20635 => x"C0C0C0A4C082B092",
 20636 => x"C0C0C0A4C082B082",
 20637 => x"C0C0C0A4C082B0F8",
 20638 => x"C0C0C0A4C082B080",
 20639 => x"C0C0C0A4C082B090",
 20640 => x"C0C0C0A4C08299C0",
 20641 => x"C0C0C0A4C08299F9",
 20642 => x"C0C0C0A4C08299A4",
 20643 => x"C0C0C0A4C08299B0",
 20644 => x"C0C0C0A4C0829999",
 20645 => x"C0C0C0A4C0829992",
 20646 => x"C0C0C0A4C0829982",
 20647 => x"C0C0C0A4C08299F8",
 20648 => x"C0C0C0A4C0829980",
 20649 => x"C0C0C0A4C0829990",
 20650 => x"C0C0C0A4C08292C0",
 20651 => x"C0C0C0A4C08292F9",
 20652 => x"C0C0C0A4C08292A4",
 20653 => x"C0C0C0A4C08292B0",
 20654 => x"C0C0C0A4C0829299",
 20655 => x"C0C0C0A4C0829292",
 20656 => x"C0C0C0A4C0829282",
 20657 => x"C0C0C0A4C08292F8",
 20658 => x"C0C0C0A4C0829280",
 20659 => x"C0C0C0A4C0829290",
 20660 => x"C0C0C0A4C08282C0",
 20661 => x"C0C0C0A4C08282F9",
 20662 => x"C0C0C0A4C08282A4",
 20663 => x"C0C0C0A4C08282B0",
 20664 => x"C0C0C0A4C0828299",
 20665 => x"C0C0C0A4C0828292",
 20666 => x"C0C0C0A4C0828282",
 20667 => x"C0C0C0A4C08282F8",
 20668 => x"C0C0C0A4C0828280",
 20669 => x"C0C0C0A4C0828290",
 20670 => x"C0C0C0A4C082F8C0",
 20671 => x"C0C0C0A4C082F8F9",
 20672 => x"C0C0C0A4C082F8A4",
 20673 => x"C0C0C0A4C082F8B0",
 20674 => x"C0C0C0A4C082F899",
 20675 => x"C0C0C0A4C082F892",
 20676 => x"C0C0C0A4C082F882",
 20677 => x"C0C0C0A4C082F8F8",
 20678 => x"C0C0C0A4C082F880",
 20679 => x"C0C0C0A4C082F890",
 20680 => x"C0C0C0A4C08280C0",
 20681 => x"C0C0C0A4C08280F9",
 20682 => x"C0C0C0A4C08280A4",
 20683 => x"C0C0C0A4C08280B0",
 20684 => x"C0C0C0A4C0828099",
 20685 => x"C0C0C0A4C0828092",
 20686 => x"C0C0C0A4C0828082",
 20687 => x"C0C0C0A4C08280F8",
 20688 => x"C0C0C0A4C0828080",
 20689 => x"C0C0C0A4C0828090",
 20690 => x"C0C0C0A4C08290C0",
 20691 => x"C0C0C0A4C08290F9",
 20692 => x"C0C0C0A4C08290A4",
 20693 => x"C0C0C0A4C08290B0",
 20694 => x"C0C0C0A4C0829099",
 20695 => x"C0C0C0A4C0829092",
 20696 => x"C0C0C0A4C0829082",
 20697 => x"C0C0C0A4C08290F8",
 20698 => x"C0C0C0A4C0829080",
 20699 => x"C0C0C0A4C0829090",
 20700 => x"C0C0C0A4C0F8C0C0",
 20701 => x"C0C0C0A4C0F8C0F9",
 20702 => x"C0C0C0A4C0F8C0A4",
 20703 => x"C0C0C0A4C0F8C0B0",
 20704 => x"C0C0C0A4C0F8C099",
 20705 => x"C0C0C0A4C0F8C092",
 20706 => x"C0C0C0A4C0F8C082",
 20707 => x"C0C0C0A4C0F8C0F8",
 20708 => x"C0C0C0A4C0F8C080",
 20709 => x"C0C0C0A4C0F8C090",
 20710 => x"C0C0C0A4C0F8F9C0",
 20711 => x"C0C0C0A4C0F8F9F9",
 20712 => x"C0C0C0A4C0F8F9A4",
 20713 => x"C0C0C0A4C0F8F9B0",
 20714 => x"C0C0C0A4C0F8F999",
 20715 => x"C0C0C0A4C0F8F992",
 20716 => x"C0C0C0A4C0F8F982",
 20717 => x"C0C0C0A4C0F8F9F8",
 20718 => x"C0C0C0A4C0F8F980",
 20719 => x"C0C0C0A4C0F8F990",
 20720 => x"C0C0C0A4C0F8A4C0",
 20721 => x"C0C0C0A4C0F8A4F9",
 20722 => x"C0C0C0A4C0F8A4A4",
 20723 => x"C0C0C0A4C0F8A4B0",
 20724 => x"C0C0C0A4C0F8A499",
 20725 => x"C0C0C0A4C0F8A492",
 20726 => x"C0C0C0A4C0F8A482",
 20727 => x"C0C0C0A4C0F8A4F8",
 20728 => x"C0C0C0A4C0F8A480",
 20729 => x"C0C0C0A4C0F8A490",
 20730 => x"C0C0C0A4C0F8B0C0",
 20731 => x"C0C0C0A4C0F8B0F9",
 20732 => x"C0C0C0A4C0F8B0A4",
 20733 => x"C0C0C0A4C0F8B0B0",
 20734 => x"C0C0C0A4C0F8B099",
 20735 => x"C0C0C0A4C0F8B092",
 20736 => x"C0C0C0A4C0F8B082",
 20737 => x"C0C0C0A4C0F8B0F8",
 20738 => x"C0C0C0A4C0F8B080",
 20739 => x"C0C0C0A4C0F8B090",
 20740 => x"C0C0C0A4C0F899C0",
 20741 => x"C0C0C0A4C0F899F9",
 20742 => x"C0C0C0A4C0F899A4",
 20743 => x"C0C0C0A4C0F899B0",
 20744 => x"C0C0C0A4C0F89999",
 20745 => x"C0C0C0A4C0F89992",
 20746 => x"C0C0C0A4C0F89982",
 20747 => x"C0C0C0A4C0F899F8",
 20748 => x"C0C0C0A4C0F89980",
 20749 => x"C0C0C0A4C0F89990",
 20750 => x"C0C0C0A4C0F892C0",
 20751 => x"C0C0C0A4C0F892F9",
 20752 => x"C0C0C0A4C0F892A4",
 20753 => x"C0C0C0A4C0F892B0",
 20754 => x"C0C0C0A4C0F89299",
 20755 => x"C0C0C0A4C0F89292",
 20756 => x"C0C0C0A4C0F89282",
 20757 => x"C0C0C0A4C0F892F8",
 20758 => x"C0C0C0A4C0F89280",
 20759 => x"C0C0C0A4C0F89290",
 20760 => x"C0C0C0A4C0F882C0",
 20761 => x"C0C0C0A4C0F882F9",
 20762 => x"C0C0C0A4C0F882A4",
 20763 => x"C0C0C0A4C0F882B0",
 20764 => x"C0C0C0A4C0F88299",
 20765 => x"C0C0C0A4C0F88292",
 20766 => x"C0C0C0A4C0F88282",
 20767 => x"C0C0C0A4C0F882F8",
 20768 => x"C0C0C0A4C0F88280",
 20769 => x"C0C0C0A4C0F88290",
 20770 => x"C0C0C0A4C0F8F8C0",
 20771 => x"C0C0C0A4C0F8F8F9",
 20772 => x"C0C0C0A4C0F8F8A4",
 20773 => x"C0C0C0A4C0F8F8B0",
 20774 => x"C0C0C0A4C0F8F899",
 20775 => x"C0C0C0A4C0F8F892",
 20776 => x"C0C0C0A4C0F8F882",
 20777 => x"C0C0C0A4C0F8F8F8",
 20778 => x"C0C0C0A4C0F8F880",
 20779 => x"C0C0C0A4C0F8F890",
 20780 => x"C0C0C0A4C0F880C0",
 20781 => x"C0C0C0A4C0F880F9",
 20782 => x"C0C0C0A4C0F880A4",
 20783 => x"C0C0C0A4C0F880B0",
 20784 => x"C0C0C0A4C0F88099",
 20785 => x"C0C0C0A4C0F88092",
 20786 => x"C0C0C0A4C0F88082",
 20787 => x"C0C0C0A4C0F880F8",
 20788 => x"C0C0C0A4C0F88080",
 20789 => x"C0C0C0A4C0F88090",
 20790 => x"C0C0C0A4C0F890C0",
 20791 => x"C0C0C0A4C0F890F9",
 20792 => x"C0C0C0A4C0F890A4",
 20793 => x"C0C0C0A4C0F890B0",
 20794 => x"C0C0C0A4C0F89099",
 20795 => x"C0C0C0A4C0F89092",
 20796 => x"C0C0C0A4C0F89082",
 20797 => x"C0C0C0A4C0F890F8",
 20798 => x"C0C0C0A4C0F89080",
 20799 => x"C0C0C0A4C0F89090",
 20800 => x"C0C0C0A4C080C0C0",
 20801 => x"C0C0C0A4C080C0F9",
 20802 => x"C0C0C0A4C080C0A4",
 20803 => x"C0C0C0A4C080C0B0",
 20804 => x"C0C0C0A4C080C099",
 20805 => x"C0C0C0A4C080C092",
 20806 => x"C0C0C0A4C080C082",
 20807 => x"C0C0C0A4C080C0F8",
 20808 => x"C0C0C0A4C080C080",
 20809 => x"C0C0C0A4C080C090",
 20810 => x"C0C0C0A4C080F9C0",
 20811 => x"C0C0C0A4C080F9F9",
 20812 => x"C0C0C0A4C080F9A4",
 20813 => x"C0C0C0A4C080F9B0",
 20814 => x"C0C0C0A4C080F999",
 20815 => x"C0C0C0A4C080F992",
 20816 => x"C0C0C0A4C080F982",
 20817 => x"C0C0C0A4C080F9F8",
 20818 => x"C0C0C0A4C080F980",
 20819 => x"C0C0C0A4C080F990",
 20820 => x"C0C0C0A4C080A4C0",
 20821 => x"C0C0C0A4C080A4F9",
 20822 => x"C0C0C0A4C080A4A4",
 20823 => x"C0C0C0A4C080A4B0",
 20824 => x"C0C0C0A4C080A499",
 20825 => x"C0C0C0A4C080A492",
 20826 => x"C0C0C0A4C080A482",
 20827 => x"C0C0C0A4C080A4F8",
 20828 => x"C0C0C0A4C080A480",
 20829 => x"C0C0C0A4C080A490",
 20830 => x"C0C0C0A4C080B0C0",
 20831 => x"C0C0C0A4C080B0F9",
 20832 => x"C0C0C0A4C080B0A4",
 20833 => x"C0C0C0A4C080B0B0",
 20834 => x"C0C0C0A4C080B099",
 20835 => x"C0C0C0A4C080B092",
 20836 => x"C0C0C0A4C080B082",
 20837 => x"C0C0C0A4C080B0F8",
 20838 => x"C0C0C0A4C080B080",
 20839 => x"C0C0C0A4C080B090",
 20840 => x"C0C0C0A4C08099C0",
 20841 => x"C0C0C0A4C08099F9",
 20842 => x"C0C0C0A4C08099A4",
 20843 => x"C0C0C0A4C08099B0",
 20844 => x"C0C0C0A4C0809999",
 20845 => x"C0C0C0A4C0809992",
 20846 => x"C0C0C0A4C0809982",
 20847 => x"C0C0C0A4C08099F8",
 20848 => x"C0C0C0A4C0809980",
 20849 => x"C0C0C0A4C0809990",
 20850 => x"C0C0C0A4C08092C0",
 20851 => x"C0C0C0A4C08092F9",
 20852 => x"C0C0C0A4C08092A4",
 20853 => x"C0C0C0A4C08092B0",
 20854 => x"C0C0C0A4C0809299",
 20855 => x"C0C0C0A4C0809292",
 20856 => x"C0C0C0A4C0809282",
 20857 => x"C0C0C0A4C08092F8",
 20858 => x"C0C0C0A4C0809280",
 20859 => x"C0C0C0A4C0809290",
 20860 => x"C0C0C0A4C08082C0",
 20861 => x"C0C0C0A4C08082F9",
 20862 => x"C0C0C0A4C08082A4",
 20863 => x"C0C0C0A4C08082B0",
 20864 => x"C0C0C0A4C0808299",
 20865 => x"C0C0C0A4C0808292",
 20866 => x"C0C0C0A4C0808282",
 20867 => x"C0C0C0A4C08082F8",
 20868 => x"C0C0C0A4C0808280",
 20869 => x"C0C0C0A4C0808290",
 20870 => x"C0C0C0A4C080F8C0",
 20871 => x"C0C0C0A4C080F8F9",
 20872 => x"C0C0C0A4C080F8A4",
 20873 => x"C0C0C0A4C080F8B0",
 20874 => x"C0C0C0A4C080F899",
 20875 => x"C0C0C0A4C080F892",
 20876 => x"C0C0C0A4C080F882",
 20877 => x"C0C0C0A4C080F8F8",
 20878 => x"C0C0C0A4C080F880",
 20879 => x"C0C0C0A4C080F890",
 20880 => x"C0C0C0A4C08080C0",
 20881 => x"C0C0C0A4C08080F9",
 20882 => x"C0C0C0A4C08080A4",
 20883 => x"C0C0C0A4C08080B0",
 20884 => x"C0C0C0A4C0808099",
 20885 => x"C0C0C0A4C0808092",
 20886 => x"C0C0C0A4C0808082",
 20887 => x"C0C0C0A4C08080F8",
 20888 => x"C0C0C0A4C0808080",
 20889 => x"C0C0C0A4C0808090",
 20890 => x"C0C0C0A4C08090C0",
 20891 => x"C0C0C0A4C08090F9",
 20892 => x"C0C0C0A4C08090A4",
 20893 => x"C0C0C0A4C08090B0",
 20894 => x"C0C0C0A4C0809099",
 20895 => x"C0C0C0A4C0809092",
 20896 => x"C0C0C0A4C0809082",
 20897 => x"C0C0C0A4C08090F8",
 20898 => x"C0C0C0A4C0809080",
 20899 => x"C0C0C0A4C0809090",
 20900 => x"C0C0C0A4C090C0C0",
 20901 => x"C0C0C0A4C090C0F9",
 20902 => x"C0C0C0A4C090C0A4",
 20903 => x"C0C0C0A4C090C0B0",
 20904 => x"C0C0C0A4C090C099",
 20905 => x"C0C0C0A4C090C092",
 20906 => x"C0C0C0A4C090C082",
 20907 => x"C0C0C0A4C090C0F8",
 20908 => x"C0C0C0A4C090C080",
 20909 => x"C0C0C0A4C090C090",
 20910 => x"C0C0C0A4C090F9C0",
 20911 => x"C0C0C0A4C090F9F9",
 20912 => x"C0C0C0A4C090F9A4",
 20913 => x"C0C0C0A4C090F9B0",
 20914 => x"C0C0C0A4C090F999",
 20915 => x"C0C0C0A4C090F992",
 20916 => x"C0C0C0A4C090F982",
 20917 => x"C0C0C0A4C090F9F8",
 20918 => x"C0C0C0A4C090F980",
 20919 => x"C0C0C0A4C090F990",
 20920 => x"C0C0C0A4C090A4C0",
 20921 => x"C0C0C0A4C090A4F9",
 20922 => x"C0C0C0A4C090A4A4",
 20923 => x"C0C0C0A4C090A4B0",
 20924 => x"C0C0C0A4C090A499",
 20925 => x"C0C0C0A4C090A492",
 20926 => x"C0C0C0A4C090A482",
 20927 => x"C0C0C0A4C090A4F8",
 20928 => x"C0C0C0A4C090A480",
 20929 => x"C0C0C0A4C090A490",
 20930 => x"C0C0C0A4C090B0C0",
 20931 => x"C0C0C0A4C090B0F9",
 20932 => x"C0C0C0A4C090B0A4",
 20933 => x"C0C0C0A4C090B0B0",
 20934 => x"C0C0C0A4C090B099",
 20935 => x"C0C0C0A4C090B092",
 20936 => x"C0C0C0A4C090B082",
 20937 => x"C0C0C0A4C090B0F8",
 20938 => x"C0C0C0A4C090B080",
 20939 => x"C0C0C0A4C090B090",
 20940 => x"C0C0C0A4C09099C0",
 20941 => x"C0C0C0A4C09099F9",
 20942 => x"C0C0C0A4C09099A4",
 20943 => x"C0C0C0A4C09099B0",
 20944 => x"C0C0C0A4C0909999",
 20945 => x"C0C0C0A4C0909992",
 20946 => x"C0C0C0A4C0909982",
 20947 => x"C0C0C0A4C09099F8",
 20948 => x"C0C0C0A4C0909980",
 20949 => x"C0C0C0A4C0909990",
 20950 => x"C0C0C0A4C09092C0",
 20951 => x"C0C0C0A4C09092F9",
 20952 => x"C0C0C0A4C09092A4",
 20953 => x"C0C0C0A4C09092B0",
 20954 => x"C0C0C0A4C0909299",
 20955 => x"C0C0C0A4C0909292",
 20956 => x"C0C0C0A4C0909282",
 20957 => x"C0C0C0A4C09092F8",
 20958 => x"C0C0C0A4C0909280",
 20959 => x"C0C0C0A4C0909290",
 20960 => x"C0C0C0A4C09082C0",
 20961 => x"C0C0C0A4C09082F9",
 20962 => x"C0C0C0A4C09082A4",
 20963 => x"C0C0C0A4C09082B0",
 20964 => x"C0C0C0A4C0908299",
 20965 => x"C0C0C0A4C0908292",
 20966 => x"C0C0C0A4C0908282",
 20967 => x"C0C0C0A4C09082F8",
 20968 => x"C0C0C0A4C0908280",
 20969 => x"C0C0C0A4C0908290",
 20970 => x"C0C0C0A4C090F8C0",
 20971 => x"C0C0C0A4C090F8F9",
 20972 => x"C0C0C0A4C090F8A4",
 20973 => x"C0C0C0A4C090F8B0",
 20974 => x"C0C0C0A4C090F899",
 20975 => x"C0C0C0A4C090F892",
 20976 => x"C0C0C0A4C090F882",
 20977 => x"C0C0C0A4C090F8F8",
 20978 => x"C0C0C0A4C090F880",
 20979 => x"C0C0C0A4C090F890",
 20980 => x"C0C0C0A4C09080C0",
 20981 => x"C0C0C0A4C09080F9",
 20982 => x"C0C0C0A4C09080A4",
 20983 => x"C0C0C0A4C09080B0",
 20984 => x"C0C0C0A4C0908099",
 20985 => x"C0C0C0A4C0908092",
 20986 => x"C0C0C0A4C0908082",
 20987 => x"C0C0C0A4C09080F8",
 20988 => x"C0C0C0A4C0908080",
 20989 => x"C0C0C0A4C0908090",
 20990 => x"C0C0C0A4C09090C0",
 20991 => x"C0C0C0A4C09090F9",
 20992 => x"C0C0C0A4C09090A4",
 20993 => x"C0C0C0A4C09090B0",
 20994 => x"C0C0C0A4C0909099",
 20995 => x"C0C0C0A4C0909092",
 20996 => x"C0C0C0A4C0909082",
 20997 => x"C0C0C0A4C09090F8",
 20998 => x"C0C0C0A4C0909080",
 20999 => x"C0C0C0A4C0909090",
 21000 => x"C0C0C0A4F9C0C0C0",
 21001 => x"C0C0C0A4F9C0C0F9",
 21002 => x"C0C0C0A4F9C0C0A4",
 21003 => x"C0C0C0A4F9C0C0B0",
 21004 => x"C0C0C0A4F9C0C099",
 21005 => x"C0C0C0A4F9C0C092",
 21006 => x"C0C0C0A4F9C0C082",
 21007 => x"C0C0C0A4F9C0C0F8",
 21008 => x"C0C0C0A4F9C0C080",
 21009 => x"C0C0C0A4F9C0C090",
 21010 => x"C0C0C0A4F9C0F9C0",
 21011 => x"C0C0C0A4F9C0F9F9",
 21012 => x"C0C0C0A4F9C0F9A4",
 21013 => x"C0C0C0A4F9C0F9B0",
 21014 => x"C0C0C0A4F9C0F999",
 21015 => x"C0C0C0A4F9C0F992",
 21016 => x"C0C0C0A4F9C0F982",
 21017 => x"C0C0C0A4F9C0F9F8",
 21018 => x"C0C0C0A4F9C0F980",
 21019 => x"C0C0C0A4F9C0F990",
 21020 => x"C0C0C0A4F9C0A4C0",
 21021 => x"C0C0C0A4F9C0A4F9",
 21022 => x"C0C0C0A4F9C0A4A4",
 21023 => x"C0C0C0A4F9C0A4B0",
 21024 => x"C0C0C0A4F9C0A499",
 21025 => x"C0C0C0A4F9C0A492",
 21026 => x"C0C0C0A4F9C0A482",
 21027 => x"C0C0C0A4F9C0A4F8",
 21028 => x"C0C0C0A4F9C0A480",
 21029 => x"C0C0C0A4F9C0A490",
 21030 => x"C0C0C0A4F9C0B0C0",
 21031 => x"C0C0C0A4F9C0B0F9",
 21032 => x"C0C0C0A4F9C0B0A4",
 21033 => x"C0C0C0A4F9C0B0B0",
 21034 => x"C0C0C0A4F9C0B099",
 21035 => x"C0C0C0A4F9C0B092",
 21036 => x"C0C0C0A4F9C0B082",
 21037 => x"C0C0C0A4F9C0B0F8",
 21038 => x"C0C0C0A4F9C0B080",
 21039 => x"C0C0C0A4F9C0B090",
 21040 => x"C0C0C0A4F9C099C0",
 21041 => x"C0C0C0A4F9C099F9",
 21042 => x"C0C0C0A4F9C099A4",
 21043 => x"C0C0C0A4F9C099B0",
 21044 => x"C0C0C0A4F9C09999",
 21045 => x"C0C0C0A4F9C09992",
 21046 => x"C0C0C0A4F9C09982",
 21047 => x"C0C0C0A4F9C099F8",
 21048 => x"C0C0C0A4F9C09980",
 21049 => x"C0C0C0A4F9C09990",
 21050 => x"C0C0C0A4F9C092C0",
 21051 => x"C0C0C0A4F9C092F9",
 21052 => x"C0C0C0A4F9C092A4",
 21053 => x"C0C0C0A4F9C092B0",
 21054 => x"C0C0C0A4F9C09299",
 21055 => x"C0C0C0A4F9C09292",
 21056 => x"C0C0C0A4F9C09282",
 21057 => x"C0C0C0A4F9C092F8",
 21058 => x"C0C0C0A4F9C09280",
 21059 => x"C0C0C0A4F9C09290",
 21060 => x"C0C0C0A4F9C082C0",
 21061 => x"C0C0C0A4F9C082F9",
 21062 => x"C0C0C0A4F9C082A4",
 21063 => x"C0C0C0A4F9C082B0",
 21064 => x"C0C0C0A4F9C08299",
 21065 => x"C0C0C0A4F9C08292",
 21066 => x"C0C0C0A4F9C08282",
 21067 => x"C0C0C0A4F9C082F8",
 21068 => x"C0C0C0A4F9C08280",
 21069 => x"C0C0C0A4F9C08290",
 21070 => x"C0C0C0A4F9C0F8C0",
 21071 => x"C0C0C0A4F9C0F8F9",
 21072 => x"C0C0C0A4F9C0F8A4",
 21073 => x"C0C0C0A4F9C0F8B0",
 21074 => x"C0C0C0A4F9C0F899",
 21075 => x"C0C0C0A4F9C0F892",
 21076 => x"C0C0C0A4F9C0F882",
 21077 => x"C0C0C0A4F9C0F8F8",
 21078 => x"C0C0C0A4F9C0F880",
 21079 => x"C0C0C0A4F9C0F890",
 21080 => x"C0C0C0A4F9C080C0",
 21081 => x"C0C0C0A4F9C080F9",
 21082 => x"C0C0C0A4F9C080A4",
 21083 => x"C0C0C0A4F9C080B0",
 21084 => x"C0C0C0A4F9C08099",
 21085 => x"C0C0C0A4F9C08092",
 21086 => x"C0C0C0A4F9C08082",
 21087 => x"C0C0C0A4F9C080F8",
 21088 => x"C0C0C0A4F9C08080",
 21089 => x"C0C0C0A4F9C08090",
 21090 => x"C0C0C0A4F9C090C0",
 21091 => x"C0C0C0A4F9C090F9",
 21092 => x"C0C0C0A4F9C090A4",
 21093 => x"C0C0C0A4F9C090B0",
 21094 => x"C0C0C0A4F9C09099",
 21095 => x"C0C0C0A4F9C09092",
 21096 => x"C0C0C0A4F9C09082",
 21097 => x"C0C0C0A4F9C090F8",
 21098 => x"C0C0C0A4F9C09080",
 21099 => x"C0C0C0A4F9C09090",
 21100 => x"C0C0C0A4F9F9C0C0",
 21101 => x"C0C0C0A4F9F9C0F9",
 21102 => x"C0C0C0A4F9F9C0A4",
 21103 => x"C0C0C0A4F9F9C0B0",
 21104 => x"C0C0C0A4F9F9C099",
 21105 => x"C0C0C0A4F9F9C092",
 21106 => x"C0C0C0A4F9F9C082",
 21107 => x"C0C0C0A4F9F9C0F8",
 21108 => x"C0C0C0A4F9F9C080",
 21109 => x"C0C0C0A4F9F9C090",
 21110 => x"C0C0C0A4F9F9F9C0",
 21111 => x"C0C0C0A4F9F9F9F9",
 21112 => x"C0C0C0A4F9F9F9A4",
 21113 => x"C0C0C0A4F9F9F9B0",
 21114 => x"C0C0C0A4F9F9F999",
 21115 => x"C0C0C0A4F9F9F992",
 21116 => x"C0C0C0A4F9F9F982",
 21117 => x"C0C0C0A4F9F9F9F8",
 21118 => x"C0C0C0A4F9F9F980",
 21119 => x"C0C0C0A4F9F9F990",
 21120 => x"C0C0C0A4F9F9A4C0",
 21121 => x"C0C0C0A4F9F9A4F9",
 21122 => x"C0C0C0A4F9F9A4A4",
 21123 => x"C0C0C0A4F9F9A4B0",
 21124 => x"C0C0C0A4F9F9A499",
 21125 => x"C0C0C0A4F9F9A492",
 21126 => x"C0C0C0A4F9F9A482",
 21127 => x"C0C0C0A4F9F9A4F8",
 21128 => x"C0C0C0A4F9F9A480",
 21129 => x"C0C0C0A4F9F9A490",
 21130 => x"C0C0C0A4F9F9B0C0",
 21131 => x"C0C0C0A4F9F9B0F9",
 21132 => x"C0C0C0A4F9F9B0A4",
 21133 => x"C0C0C0A4F9F9B0B0",
 21134 => x"C0C0C0A4F9F9B099",
 21135 => x"C0C0C0A4F9F9B092",
 21136 => x"C0C0C0A4F9F9B082",
 21137 => x"C0C0C0A4F9F9B0F8",
 21138 => x"C0C0C0A4F9F9B080",
 21139 => x"C0C0C0A4F9F9B090",
 21140 => x"C0C0C0A4F9F999C0",
 21141 => x"C0C0C0A4F9F999F9",
 21142 => x"C0C0C0A4F9F999A4",
 21143 => x"C0C0C0A4F9F999B0",
 21144 => x"C0C0C0A4F9F99999",
 21145 => x"C0C0C0A4F9F99992",
 21146 => x"C0C0C0A4F9F99982",
 21147 => x"C0C0C0A4F9F999F8",
 21148 => x"C0C0C0A4F9F99980",
 21149 => x"C0C0C0A4F9F99990",
 21150 => x"C0C0C0A4F9F992C0",
 21151 => x"C0C0C0A4F9F992F9",
 21152 => x"C0C0C0A4F9F992A4",
 21153 => x"C0C0C0A4F9F992B0",
 21154 => x"C0C0C0A4F9F99299",
 21155 => x"C0C0C0A4F9F99292",
 21156 => x"C0C0C0A4F9F99282",
 21157 => x"C0C0C0A4F9F992F8",
 21158 => x"C0C0C0A4F9F99280",
 21159 => x"C0C0C0A4F9F99290",
 21160 => x"C0C0C0A4F9F982C0",
 21161 => x"C0C0C0A4F9F982F9",
 21162 => x"C0C0C0A4F9F982A4",
 21163 => x"C0C0C0A4F9F982B0",
 21164 => x"C0C0C0A4F9F98299",
 21165 => x"C0C0C0A4F9F98292",
 21166 => x"C0C0C0A4F9F98282",
 21167 => x"C0C0C0A4F9F982F8",
 21168 => x"C0C0C0A4F9F98280",
 21169 => x"C0C0C0A4F9F98290",
 21170 => x"C0C0C0A4F9F9F8C0",
 21171 => x"C0C0C0A4F9F9F8F9",
 21172 => x"C0C0C0A4F9F9F8A4",
 21173 => x"C0C0C0A4F9F9F8B0",
 21174 => x"C0C0C0A4F9F9F899",
 21175 => x"C0C0C0A4F9F9F892",
 21176 => x"C0C0C0A4F9F9F882",
 21177 => x"C0C0C0A4F9F9F8F8",
 21178 => x"C0C0C0A4F9F9F880",
 21179 => x"C0C0C0A4F9F9F890",
 21180 => x"C0C0C0A4F9F980C0",
 21181 => x"C0C0C0A4F9F980F9",
 21182 => x"C0C0C0A4F9F980A4",
 21183 => x"C0C0C0A4F9F980B0",
 21184 => x"C0C0C0A4F9F98099",
 21185 => x"C0C0C0A4F9F98092",
 21186 => x"C0C0C0A4F9F98082",
 21187 => x"C0C0C0A4F9F980F8",
 21188 => x"C0C0C0A4F9F98080",
 21189 => x"C0C0C0A4F9F98090",
 21190 => x"C0C0C0A4F9F990C0",
 21191 => x"C0C0C0A4F9F990F9",
 21192 => x"C0C0C0A4F9F990A4",
 21193 => x"C0C0C0A4F9F990B0",
 21194 => x"C0C0C0A4F9F99099",
 21195 => x"C0C0C0A4F9F99092",
 21196 => x"C0C0C0A4F9F99082",
 21197 => x"C0C0C0A4F9F990F8",
 21198 => x"C0C0C0A4F9F99080",
 21199 => x"C0C0C0A4F9F99090",
 21200 => x"C0C0C0A4F9A4C0C0",
 21201 => x"C0C0C0A4F9A4C0F9",
 21202 => x"C0C0C0A4F9A4C0A4",
 21203 => x"C0C0C0A4F9A4C0B0",
 21204 => x"C0C0C0A4F9A4C099",
 21205 => x"C0C0C0A4F9A4C092",
 21206 => x"C0C0C0A4F9A4C082",
 21207 => x"C0C0C0A4F9A4C0F8",
 21208 => x"C0C0C0A4F9A4C080",
 21209 => x"C0C0C0A4F9A4C090",
 21210 => x"C0C0C0A4F9A4F9C0",
 21211 => x"C0C0C0A4F9A4F9F9",
 21212 => x"C0C0C0A4F9A4F9A4",
 21213 => x"C0C0C0A4F9A4F9B0",
 21214 => x"C0C0C0A4F9A4F999",
 21215 => x"C0C0C0A4F9A4F992",
 21216 => x"C0C0C0A4F9A4F982",
 21217 => x"C0C0C0A4F9A4F9F8",
 21218 => x"C0C0C0A4F9A4F980",
 21219 => x"C0C0C0A4F9A4F990",
 21220 => x"C0C0C0A4F9A4A4C0",
 21221 => x"C0C0C0A4F9A4A4F9",
 21222 => x"C0C0C0A4F9A4A4A4",
 21223 => x"C0C0C0A4F9A4A4B0",
 21224 => x"C0C0C0A4F9A4A499",
 21225 => x"C0C0C0A4F9A4A492",
 21226 => x"C0C0C0A4F9A4A482",
 21227 => x"C0C0C0A4F9A4A4F8",
 21228 => x"C0C0C0A4F9A4A480",
 21229 => x"C0C0C0A4F9A4A490",
 21230 => x"C0C0C0A4F9A4B0C0",
 21231 => x"C0C0C0A4F9A4B0F9",
 21232 => x"C0C0C0A4F9A4B0A4",
 21233 => x"C0C0C0A4F9A4B0B0",
 21234 => x"C0C0C0A4F9A4B099",
 21235 => x"C0C0C0A4F9A4B092",
 21236 => x"C0C0C0A4F9A4B082",
 21237 => x"C0C0C0A4F9A4B0F8",
 21238 => x"C0C0C0A4F9A4B080",
 21239 => x"C0C0C0A4F9A4B090",
 21240 => x"C0C0C0A4F9A499C0",
 21241 => x"C0C0C0A4F9A499F9",
 21242 => x"C0C0C0A4F9A499A4",
 21243 => x"C0C0C0A4F9A499B0",
 21244 => x"C0C0C0A4F9A49999",
 21245 => x"C0C0C0A4F9A49992",
 21246 => x"C0C0C0A4F9A49982",
 21247 => x"C0C0C0A4F9A499F8",
 21248 => x"C0C0C0A4F9A49980",
 21249 => x"C0C0C0A4F9A49990",
 21250 => x"C0C0C0A4F9A492C0",
 21251 => x"C0C0C0A4F9A492F9",
 21252 => x"C0C0C0A4F9A492A4",
 21253 => x"C0C0C0A4F9A492B0",
 21254 => x"C0C0C0A4F9A49299",
 21255 => x"C0C0C0A4F9A49292",
 21256 => x"C0C0C0A4F9A49282",
 21257 => x"C0C0C0A4F9A492F8",
 21258 => x"C0C0C0A4F9A49280",
 21259 => x"C0C0C0A4F9A49290",
 21260 => x"C0C0C0A4F9A482C0",
 21261 => x"C0C0C0A4F9A482F9",
 21262 => x"C0C0C0A4F9A482A4",
 21263 => x"C0C0C0A4F9A482B0",
 21264 => x"C0C0C0A4F9A48299",
 21265 => x"C0C0C0A4F9A48292",
 21266 => x"C0C0C0A4F9A48282",
 21267 => x"C0C0C0A4F9A482F8",
 21268 => x"C0C0C0A4F9A48280",
 21269 => x"C0C0C0A4F9A48290",
 21270 => x"C0C0C0A4F9A4F8C0",
 21271 => x"C0C0C0A4F9A4F8F9",
 21272 => x"C0C0C0A4F9A4F8A4",
 21273 => x"C0C0C0A4F9A4F8B0",
 21274 => x"C0C0C0A4F9A4F899",
 21275 => x"C0C0C0A4F9A4F892",
 21276 => x"C0C0C0A4F9A4F882",
 21277 => x"C0C0C0A4F9A4F8F8",
 21278 => x"C0C0C0A4F9A4F880",
 21279 => x"C0C0C0A4F9A4F890",
 21280 => x"C0C0C0A4F9A480C0",
 21281 => x"C0C0C0A4F9A480F9",
 21282 => x"C0C0C0A4F9A480A4",
 21283 => x"C0C0C0A4F9A480B0",
 21284 => x"C0C0C0A4F9A48099",
 21285 => x"C0C0C0A4F9A48092",
 21286 => x"C0C0C0A4F9A48082",
 21287 => x"C0C0C0A4F9A480F8",
 21288 => x"C0C0C0A4F9A48080",
 21289 => x"C0C0C0A4F9A48090",
 21290 => x"C0C0C0A4F9A490C0",
 21291 => x"C0C0C0A4F9A490F9",
 21292 => x"C0C0C0A4F9A490A4",
 21293 => x"C0C0C0A4F9A490B0",
 21294 => x"C0C0C0A4F9A49099",
 21295 => x"C0C0C0A4F9A49092",
 21296 => x"C0C0C0A4F9A49082",
 21297 => x"C0C0C0A4F9A490F8",
 21298 => x"C0C0C0A4F9A49080",
 21299 => x"C0C0C0A4F9A49090",
 21300 => x"C0C0C0A4F9B0C0C0",
 21301 => x"C0C0C0A4F9B0C0F9",
 21302 => x"C0C0C0A4F9B0C0A4",
 21303 => x"C0C0C0A4F9B0C0B0",
 21304 => x"C0C0C0A4F9B0C099",
 21305 => x"C0C0C0A4F9B0C092",
 21306 => x"C0C0C0A4F9B0C082",
 21307 => x"C0C0C0A4F9B0C0F8",
 21308 => x"C0C0C0A4F9B0C080",
 21309 => x"C0C0C0A4F9B0C090",
 21310 => x"C0C0C0A4F9B0F9C0",
 21311 => x"C0C0C0A4F9B0F9F9",
 21312 => x"C0C0C0A4F9B0F9A4",
 21313 => x"C0C0C0A4F9B0F9B0",
 21314 => x"C0C0C0A4F9B0F999",
 21315 => x"C0C0C0A4F9B0F992",
 21316 => x"C0C0C0A4F9B0F982",
 21317 => x"C0C0C0A4F9B0F9F8",
 21318 => x"C0C0C0A4F9B0F980",
 21319 => x"C0C0C0A4F9B0F990",
 21320 => x"C0C0C0A4F9B0A4C0",
 21321 => x"C0C0C0A4F9B0A4F9",
 21322 => x"C0C0C0A4F9B0A4A4",
 21323 => x"C0C0C0A4F9B0A4B0",
 21324 => x"C0C0C0A4F9B0A499",
 21325 => x"C0C0C0A4F9B0A492",
 21326 => x"C0C0C0A4F9B0A482",
 21327 => x"C0C0C0A4F9B0A4F8",
 21328 => x"C0C0C0A4F9B0A480",
 21329 => x"C0C0C0A4F9B0A490",
 21330 => x"C0C0C0A4F9B0B0C0",
 21331 => x"C0C0C0A4F9B0B0F9",
 21332 => x"C0C0C0A4F9B0B0A4",
 21333 => x"C0C0C0A4F9B0B0B0",
 21334 => x"C0C0C0A4F9B0B099",
 21335 => x"C0C0C0A4F9B0B092",
 21336 => x"C0C0C0A4F9B0B082",
 21337 => x"C0C0C0A4F9B0B0F8",
 21338 => x"C0C0C0A4F9B0B080",
 21339 => x"C0C0C0A4F9B0B090",
 21340 => x"C0C0C0A4F9B099C0",
 21341 => x"C0C0C0A4F9B099F9",
 21342 => x"C0C0C0A4F9B099A4",
 21343 => x"C0C0C0A4F9B099B0",
 21344 => x"C0C0C0A4F9B09999",
 21345 => x"C0C0C0A4F9B09992",
 21346 => x"C0C0C0A4F9B09982",
 21347 => x"C0C0C0A4F9B099F8",
 21348 => x"C0C0C0A4F9B09980",
 21349 => x"C0C0C0A4F9B09990",
 21350 => x"C0C0C0A4F9B092C0",
 21351 => x"C0C0C0A4F9B092F9",
 21352 => x"C0C0C0A4F9B092A4",
 21353 => x"C0C0C0A4F9B092B0",
 21354 => x"C0C0C0A4F9B09299",
 21355 => x"C0C0C0A4F9B09292",
 21356 => x"C0C0C0A4F9B09282",
 21357 => x"C0C0C0A4F9B092F8",
 21358 => x"C0C0C0A4F9B09280",
 21359 => x"C0C0C0A4F9B09290",
 21360 => x"C0C0C0A4F9B082C0",
 21361 => x"C0C0C0A4F9B082F9",
 21362 => x"C0C0C0A4F9B082A4",
 21363 => x"C0C0C0A4F9B082B0",
 21364 => x"C0C0C0A4F9B08299",
 21365 => x"C0C0C0A4F9B08292",
 21366 => x"C0C0C0A4F9B08282",
 21367 => x"C0C0C0A4F9B082F8",
 21368 => x"C0C0C0A4F9B08280",
 21369 => x"C0C0C0A4F9B08290",
 21370 => x"C0C0C0A4F9B0F8C0",
 21371 => x"C0C0C0A4F9B0F8F9",
 21372 => x"C0C0C0A4F9B0F8A4",
 21373 => x"C0C0C0A4F9B0F8B0",
 21374 => x"C0C0C0A4F9B0F899",
 21375 => x"C0C0C0A4F9B0F892",
 21376 => x"C0C0C0A4F9B0F882",
 21377 => x"C0C0C0A4F9B0F8F8",
 21378 => x"C0C0C0A4F9B0F880",
 21379 => x"C0C0C0A4F9B0F890",
 21380 => x"C0C0C0A4F9B080C0",
 21381 => x"C0C0C0A4F9B080F9",
 21382 => x"C0C0C0A4F9B080A4",
 21383 => x"C0C0C0A4F9B080B0",
 21384 => x"C0C0C0A4F9B08099",
 21385 => x"C0C0C0A4F9B08092",
 21386 => x"C0C0C0A4F9B08082",
 21387 => x"C0C0C0A4F9B080F8",
 21388 => x"C0C0C0A4F9B08080",
 21389 => x"C0C0C0A4F9B08090",
 21390 => x"C0C0C0A4F9B090C0",
 21391 => x"C0C0C0A4F9B090F9",
 21392 => x"C0C0C0A4F9B090A4",
 21393 => x"C0C0C0A4F9B090B0",
 21394 => x"C0C0C0A4F9B09099",
 21395 => x"C0C0C0A4F9B09092",
 21396 => x"C0C0C0A4F9B09082",
 21397 => x"C0C0C0A4F9B090F8",
 21398 => x"C0C0C0A4F9B09080",
 21399 => x"C0C0C0A4F9B09090",
 21400 => x"C0C0C0A4F999C0C0",
 21401 => x"C0C0C0A4F999C0F9",
 21402 => x"C0C0C0A4F999C0A4",
 21403 => x"C0C0C0A4F999C0B0",
 21404 => x"C0C0C0A4F999C099",
 21405 => x"C0C0C0A4F999C092",
 21406 => x"C0C0C0A4F999C082",
 21407 => x"C0C0C0A4F999C0F8",
 21408 => x"C0C0C0A4F999C080",
 21409 => x"C0C0C0A4F999C090",
 21410 => x"C0C0C0A4F999F9C0",
 21411 => x"C0C0C0A4F999F9F9",
 21412 => x"C0C0C0A4F999F9A4",
 21413 => x"C0C0C0A4F999F9B0",
 21414 => x"C0C0C0A4F999F999",
 21415 => x"C0C0C0A4F999F992",
 21416 => x"C0C0C0A4F999F982",
 21417 => x"C0C0C0A4F999F9F8",
 21418 => x"C0C0C0A4F999F980",
 21419 => x"C0C0C0A4F999F990",
 21420 => x"C0C0C0A4F999A4C0",
 21421 => x"C0C0C0A4F999A4F9",
 21422 => x"C0C0C0A4F999A4A4",
 21423 => x"C0C0C0A4F999A4B0",
 21424 => x"C0C0C0A4F999A499",
 21425 => x"C0C0C0A4F999A492",
 21426 => x"C0C0C0A4F999A482",
 21427 => x"C0C0C0A4F999A4F8",
 21428 => x"C0C0C0A4F999A480",
 21429 => x"C0C0C0A4F999A490",
 21430 => x"C0C0C0A4F999B0C0",
 21431 => x"C0C0C0A4F999B0F9",
 21432 => x"C0C0C0A4F999B0A4",
 21433 => x"C0C0C0A4F999B0B0",
 21434 => x"C0C0C0A4F999B099",
 21435 => x"C0C0C0A4F999B092",
 21436 => x"C0C0C0A4F999B082",
 21437 => x"C0C0C0A4F999B0F8",
 21438 => x"C0C0C0A4F999B080",
 21439 => x"C0C0C0A4F999B090",
 21440 => x"C0C0C0A4F99999C0",
 21441 => x"C0C0C0A4F99999F9",
 21442 => x"C0C0C0A4F99999A4",
 21443 => x"C0C0C0A4F99999B0",
 21444 => x"C0C0C0A4F9999999",
 21445 => x"C0C0C0A4F9999992",
 21446 => x"C0C0C0A4F9999982",
 21447 => x"C0C0C0A4F99999F8",
 21448 => x"C0C0C0A4F9999980",
 21449 => x"C0C0C0A4F9999990",
 21450 => x"C0C0C0A4F99992C0",
 21451 => x"C0C0C0A4F99992F9",
 21452 => x"C0C0C0A4F99992A4",
 21453 => x"C0C0C0A4F99992B0",
 21454 => x"C0C0C0A4F9999299",
 21455 => x"C0C0C0A4F9999292",
 21456 => x"C0C0C0A4F9999282",
 21457 => x"C0C0C0A4F99992F8",
 21458 => x"C0C0C0A4F9999280",
 21459 => x"C0C0C0A4F9999290",
 21460 => x"C0C0C0A4F99982C0",
 21461 => x"C0C0C0A4F99982F9",
 21462 => x"C0C0C0A4F99982A4",
 21463 => x"C0C0C0A4F99982B0",
 21464 => x"C0C0C0A4F9998299",
 21465 => x"C0C0C0A4F9998292",
 21466 => x"C0C0C0A4F9998282",
 21467 => x"C0C0C0A4F99982F8",
 21468 => x"C0C0C0A4F9998280",
 21469 => x"C0C0C0A4F9998290",
 21470 => x"C0C0C0A4F999F8C0",
 21471 => x"C0C0C0A4F999F8F9",
 21472 => x"C0C0C0A4F999F8A4",
 21473 => x"C0C0C0A4F999F8B0",
 21474 => x"C0C0C0A4F999F899",
 21475 => x"C0C0C0A4F999F892",
 21476 => x"C0C0C0A4F999F882",
 21477 => x"C0C0C0A4F999F8F8",
 21478 => x"C0C0C0A4F999F880",
 21479 => x"C0C0C0A4F999F890",
 21480 => x"C0C0C0A4F99980C0",
 21481 => x"C0C0C0A4F99980F9",
 21482 => x"C0C0C0A4F99980A4",
 21483 => x"C0C0C0A4F99980B0",
 21484 => x"C0C0C0A4F9998099",
 21485 => x"C0C0C0A4F9998092",
 21486 => x"C0C0C0A4F9998082",
 21487 => x"C0C0C0A4F99980F8",
 21488 => x"C0C0C0A4F9998080",
 21489 => x"C0C0C0A4F9998090",
 21490 => x"C0C0C0A4F99990C0",
 21491 => x"C0C0C0A4F99990F9",
 21492 => x"C0C0C0A4F99990A4",
 21493 => x"C0C0C0A4F99990B0",
 21494 => x"C0C0C0A4F9999099",
 21495 => x"C0C0C0A4F9999092",
 21496 => x"C0C0C0A4F9999082",
 21497 => x"C0C0C0A4F99990F8",
 21498 => x"C0C0C0A4F9999080",
 21499 => x"C0C0C0A4F9999090",
 21500 => x"C0C0C0A4F992C0C0",
 21501 => x"C0C0C0A4F992C0F9",
 21502 => x"C0C0C0A4F992C0A4",
 21503 => x"C0C0C0A4F992C0B0",
 21504 => x"C0C0C0A4F992C099",
 21505 => x"C0C0C0A4F992C092",
 21506 => x"C0C0C0A4F992C082",
 21507 => x"C0C0C0A4F992C0F8",
 21508 => x"C0C0C0A4F992C080",
 21509 => x"C0C0C0A4F992C090",
 21510 => x"C0C0C0A4F992F9C0",
 21511 => x"C0C0C0A4F992F9F9",
 21512 => x"C0C0C0A4F992F9A4",
 21513 => x"C0C0C0A4F992F9B0",
 21514 => x"C0C0C0A4F992F999",
 21515 => x"C0C0C0A4F992F992",
 21516 => x"C0C0C0A4F992F982",
 21517 => x"C0C0C0A4F992F9F8",
 21518 => x"C0C0C0A4F992F980",
 21519 => x"C0C0C0A4F992F990",
 21520 => x"C0C0C0A4F992A4C0",
 21521 => x"C0C0C0A4F992A4F9",
 21522 => x"C0C0C0A4F992A4A4",
 21523 => x"C0C0C0A4F992A4B0",
 21524 => x"C0C0C0A4F992A499",
 21525 => x"C0C0C0A4F992A492",
 21526 => x"C0C0C0A4F992A482",
 21527 => x"C0C0C0A4F992A4F8",
 21528 => x"C0C0C0A4F992A480",
 21529 => x"C0C0C0A4F992A490",
 21530 => x"C0C0C0A4F992B0C0",
 21531 => x"C0C0C0A4F992B0F9",
 21532 => x"C0C0C0A4F992B0A4",
 21533 => x"C0C0C0A4F992B0B0",
 21534 => x"C0C0C0A4F992B099",
 21535 => x"C0C0C0A4F992B092",
 21536 => x"C0C0C0A4F992B082",
 21537 => x"C0C0C0A4F992B0F8",
 21538 => x"C0C0C0A4F992B080",
 21539 => x"C0C0C0A4F992B090",
 21540 => x"C0C0C0A4F99299C0",
 21541 => x"C0C0C0A4F99299F9",
 21542 => x"C0C0C0A4F99299A4",
 21543 => x"C0C0C0A4F99299B0",
 21544 => x"C0C0C0A4F9929999",
 21545 => x"C0C0C0A4F9929992",
 21546 => x"C0C0C0A4F9929982",
 21547 => x"C0C0C0A4F99299F8",
 21548 => x"C0C0C0A4F9929980",
 21549 => x"C0C0C0A4F9929990",
 21550 => x"C0C0C0A4F99292C0",
 21551 => x"C0C0C0A4F99292F9",
 21552 => x"C0C0C0A4F99292A4",
 21553 => x"C0C0C0A4F99292B0",
 21554 => x"C0C0C0A4F9929299",
 21555 => x"C0C0C0A4F9929292",
 21556 => x"C0C0C0A4F9929282",
 21557 => x"C0C0C0A4F99292F8",
 21558 => x"C0C0C0A4F9929280",
 21559 => x"C0C0C0A4F9929290",
 21560 => x"C0C0C0A4F99282C0",
 21561 => x"C0C0C0A4F99282F9",
 21562 => x"C0C0C0A4F99282A4",
 21563 => x"C0C0C0A4F99282B0",
 21564 => x"C0C0C0A4F9928299",
 21565 => x"C0C0C0A4F9928292",
 21566 => x"C0C0C0A4F9928282",
 21567 => x"C0C0C0A4F99282F8",
 21568 => x"C0C0C0A4F9928280",
 21569 => x"C0C0C0A4F9928290",
 21570 => x"C0C0C0A4F992F8C0",
 21571 => x"C0C0C0A4F992F8F9",
 21572 => x"C0C0C0A4F992F8A4",
 21573 => x"C0C0C0A4F992F8B0",
 21574 => x"C0C0C0A4F992F899",
 21575 => x"C0C0C0A4F992F892",
 21576 => x"C0C0C0A4F992F882",
 21577 => x"C0C0C0A4F992F8F8",
 21578 => x"C0C0C0A4F992F880",
 21579 => x"C0C0C0A4F992F890",
 21580 => x"C0C0C0A4F99280C0",
 21581 => x"C0C0C0A4F99280F9",
 21582 => x"C0C0C0A4F99280A4",
 21583 => x"C0C0C0A4F99280B0",
 21584 => x"C0C0C0A4F9928099",
 21585 => x"C0C0C0A4F9928092",
 21586 => x"C0C0C0A4F9928082",
 21587 => x"C0C0C0A4F99280F8",
 21588 => x"C0C0C0A4F9928080",
 21589 => x"C0C0C0A4F9928090",
 21590 => x"C0C0C0A4F99290C0",
 21591 => x"C0C0C0A4F99290F9",
 21592 => x"C0C0C0A4F99290A4",
 21593 => x"C0C0C0A4F99290B0",
 21594 => x"C0C0C0A4F9929099",
 21595 => x"C0C0C0A4F9929092",
 21596 => x"C0C0C0A4F9929082",
 21597 => x"C0C0C0A4F99290F8",
 21598 => x"C0C0C0A4F9929080",
 21599 => x"C0C0C0A4F9929090",
 21600 => x"C0C0C0A4F982C0C0",
 21601 => x"C0C0C0A4F982C0F9",
 21602 => x"C0C0C0A4F982C0A4",
 21603 => x"C0C0C0A4F982C0B0",
 21604 => x"C0C0C0A4F982C099",
 21605 => x"C0C0C0A4F982C092",
 21606 => x"C0C0C0A4F982C082",
 21607 => x"C0C0C0A4F982C0F8",
 21608 => x"C0C0C0A4F982C080",
 21609 => x"C0C0C0A4F982C090",
 21610 => x"C0C0C0A4F982F9C0",
 21611 => x"C0C0C0A4F982F9F9",
 21612 => x"C0C0C0A4F982F9A4",
 21613 => x"C0C0C0A4F982F9B0",
 21614 => x"C0C0C0A4F982F999",
 21615 => x"C0C0C0A4F982F992",
 21616 => x"C0C0C0A4F982F982",
 21617 => x"C0C0C0A4F982F9F8",
 21618 => x"C0C0C0A4F982F980",
 21619 => x"C0C0C0A4F982F990",
 21620 => x"C0C0C0A4F982A4C0",
 21621 => x"C0C0C0A4F982A4F9",
 21622 => x"C0C0C0A4F982A4A4",
 21623 => x"C0C0C0A4F982A4B0",
 21624 => x"C0C0C0A4F982A499",
 21625 => x"C0C0C0A4F982A492",
 21626 => x"C0C0C0A4F982A482",
 21627 => x"C0C0C0A4F982A4F8",
 21628 => x"C0C0C0A4F982A480",
 21629 => x"C0C0C0A4F982A490",
 21630 => x"C0C0C0A4F982B0C0",
 21631 => x"C0C0C0A4F982B0F9",
 21632 => x"C0C0C0A4F982B0A4",
 21633 => x"C0C0C0A4F982B0B0",
 21634 => x"C0C0C0A4F982B099",
 21635 => x"C0C0C0A4F982B092",
 21636 => x"C0C0C0A4F982B082",
 21637 => x"C0C0C0A4F982B0F8",
 21638 => x"C0C0C0A4F982B080",
 21639 => x"C0C0C0A4F982B090",
 21640 => x"C0C0C0A4F98299C0",
 21641 => x"C0C0C0A4F98299F9",
 21642 => x"C0C0C0A4F98299A4",
 21643 => x"C0C0C0A4F98299B0",
 21644 => x"C0C0C0A4F9829999",
 21645 => x"C0C0C0A4F9829992",
 21646 => x"C0C0C0A4F9829982",
 21647 => x"C0C0C0A4F98299F8",
 21648 => x"C0C0C0A4F9829980",
 21649 => x"C0C0C0A4F9829990",
 21650 => x"C0C0C0A4F98292C0",
 21651 => x"C0C0C0A4F98292F9",
 21652 => x"C0C0C0A4F98292A4",
 21653 => x"C0C0C0A4F98292B0",
 21654 => x"C0C0C0A4F9829299",
 21655 => x"C0C0C0A4F9829292",
 21656 => x"C0C0C0A4F9829282",
 21657 => x"C0C0C0A4F98292F8",
 21658 => x"C0C0C0A4F9829280",
 21659 => x"C0C0C0A4F9829290",
 21660 => x"C0C0C0A4F98282C0",
 21661 => x"C0C0C0A4F98282F9",
 21662 => x"C0C0C0A4F98282A4",
 21663 => x"C0C0C0A4F98282B0",
 21664 => x"C0C0C0A4F9828299",
 21665 => x"C0C0C0A4F9828292",
 21666 => x"C0C0C0A4F9828282",
 21667 => x"C0C0C0A4F98282F8",
 21668 => x"C0C0C0A4F9828280",
 21669 => x"C0C0C0A4F9828290",
 21670 => x"C0C0C0A4F982F8C0",
 21671 => x"C0C0C0A4F982F8F9",
 21672 => x"C0C0C0A4F982F8A4",
 21673 => x"C0C0C0A4F982F8B0",
 21674 => x"C0C0C0A4F982F899",
 21675 => x"C0C0C0A4F982F892",
 21676 => x"C0C0C0A4F982F882",
 21677 => x"C0C0C0A4F982F8F8",
 21678 => x"C0C0C0A4F982F880",
 21679 => x"C0C0C0A4F982F890",
 21680 => x"C0C0C0A4F98280C0",
 21681 => x"C0C0C0A4F98280F9",
 21682 => x"C0C0C0A4F98280A4",
 21683 => x"C0C0C0A4F98280B0",
 21684 => x"C0C0C0A4F9828099",
 21685 => x"C0C0C0A4F9828092",
 21686 => x"C0C0C0A4F9828082",
 21687 => x"C0C0C0A4F98280F8",
 21688 => x"C0C0C0A4F9828080",
 21689 => x"C0C0C0A4F9828090",
 21690 => x"C0C0C0A4F98290C0",
 21691 => x"C0C0C0A4F98290F9",
 21692 => x"C0C0C0A4F98290A4",
 21693 => x"C0C0C0A4F98290B0",
 21694 => x"C0C0C0A4F9829099",
 21695 => x"C0C0C0A4F9829092",
 21696 => x"C0C0C0A4F9829082",
 21697 => x"C0C0C0A4F98290F8",
 21698 => x"C0C0C0A4F9829080",
 21699 => x"C0C0C0A4F9829090",
 21700 => x"C0C0C0A4F9F8C0C0",
 21701 => x"C0C0C0A4F9F8C0F9",
 21702 => x"C0C0C0A4F9F8C0A4",
 21703 => x"C0C0C0A4F9F8C0B0",
 21704 => x"C0C0C0A4F9F8C099",
 21705 => x"C0C0C0A4F9F8C092",
 21706 => x"C0C0C0A4F9F8C082",
 21707 => x"C0C0C0A4F9F8C0F8",
 21708 => x"C0C0C0A4F9F8C080",
 21709 => x"C0C0C0A4F9F8C090",
 21710 => x"C0C0C0A4F9F8F9C0",
 21711 => x"C0C0C0A4F9F8F9F9",
 21712 => x"C0C0C0A4F9F8F9A4",
 21713 => x"C0C0C0A4F9F8F9B0",
 21714 => x"C0C0C0A4F9F8F999",
 21715 => x"C0C0C0A4F9F8F992",
 21716 => x"C0C0C0A4F9F8F982",
 21717 => x"C0C0C0A4F9F8F9F8",
 21718 => x"C0C0C0A4F9F8F980",
 21719 => x"C0C0C0A4F9F8F990",
 21720 => x"C0C0C0A4F9F8A4C0",
 21721 => x"C0C0C0A4F9F8A4F9",
 21722 => x"C0C0C0A4F9F8A4A4",
 21723 => x"C0C0C0A4F9F8A4B0",
 21724 => x"C0C0C0A4F9F8A499",
 21725 => x"C0C0C0A4F9F8A492",
 21726 => x"C0C0C0A4F9F8A482",
 21727 => x"C0C0C0A4F9F8A4F8",
 21728 => x"C0C0C0A4F9F8A480",
 21729 => x"C0C0C0A4F9F8A490",
 21730 => x"C0C0C0A4F9F8B0C0",
 21731 => x"C0C0C0A4F9F8B0F9",
 21732 => x"C0C0C0A4F9F8B0A4",
 21733 => x"C0C0C0A4F9F8B0B0",
 21734 => x"C0C0C0A4F9F8B099",
 21735 => x"C0C0C0A4F9F8B092",
 21736 => x"C0C0C0A4F9F8B082",
 21737 => x"C0C0C0A4F9F8B0F8",
 21738 => x"C0C0C0A4F9F8B080",
 21739 => x"C0C0C0A4F9F8B090",
 21740 => x"C0C0C0A4F9F899C0",
 21741 => x"C0C0C0A4F9F899F9",
 21742 => x"C0C0C0A4F9F899A4",
 21743 => x"C0C0C0A4F9F899B0",
 21744 => x"C0C0C0A4F9F89999",
 21745 => x"C0C0C0A4F9F89992",
 21746 => x"C0C0C0A4F9F89982",
 21747 => x"C0C0C0A4F9F899F8",
 21748 => x"C0C0C0A4F9F89980",
 21749 => x"C0C0C0A4F9F89990",
 21750 => x"C0C0C0A4F9F892C0",
 21751 => x"C0C0C0A4F9F892F9",
 21752 => x"C0C0C0A4F9F892A4",
 21753 => x"C0C0C0A4F9F892B0",
 21754 => x"C0C0C0A4F9F89299",
 21755 => x"C0C0C0A4F9F89292",
 21756 => x"C0C0C0A4F9F89282",
 21757 => x"C0C0C0A4F9F892F8",
 21758 => x"C0C0C0A4F9F89280",
 21759 => x"C0C0C0A4F9F89290",
 21760 => x"C0C0C0A4F9F882C0",
 21761 => x"C0C0C0A4F9F882F9",
 21762 => x"C0C0C0A4F9F882A4",
 21763 => x"C0C0C0A4F9F882B0",
 21764 => x"C0C0C0A4F9F88299",
 21765 => x"C0C0C0A4F9F88292",
 21766 => x"C0C0C0A4F9F88282",
 21767 => x"C0C0C0A4F9F882F8",
 21768 => x"C0C0C0A4F9F88280",
 21769 => x"C0C0C0A4F9F88290",
 21770 => x"C0C0C0A4F9F8F8C0",
 21771 => x"C0C0C0A4F9F8F8F9",
 21772 => x"C0C0C0A4F9F8F8A4",
 21773 => x"C0C0C0A4F9F8F8B0",
 21774 => x"C0C0C0A4F9F8F899",
 21775 => x"C0C0C0A4F9F8F892",
 21776 => x"C0C0C0A4F9F8F882",
 21777 => x"C0C0C0A4F9F8F8F8",
 21778 => x"C0C0C0A4F9F8F880",
 21779 => x"C0C0C0A4F9F8F890",
 21780 => x"C0C0C0A4F9F880C0",
 21781 => x"C0C0C0A4F9F880F9",
 21782 => x"C0C0C0A4F9F880A4",
 21783 => x"C0C0C0A4F9F880B0",
 21784 => x"C0C0C0A4F9F88099",
 21785 => x"C0C0C0A4F9F88092",
 21786 => x"C0C0C0A4F9F88082",
 21787 => x"C0C0C0A4F9F880F8",
 21788 => x"C0C0C0A4F9F88080",
 21789 => x"C0C0C0A4F9F88090",
 21790 => x"C0C0C0A4F9F890C0",
 21791 => x"C0C0C0A4F9F890F9",
 21792 => x"C0C0C0A4F9F890A4",
 21793 => x"C0C0C0A4F9F890B0",
 21794 => x"C0C0C0A4F9F89099",
 21795 => x"C0C0C0A4F9F89092",
 21796 => x"C0C0C0A4F9F89082",
 21797 => x"C0C0C0A4F9F890F8",
 21798 => x"C0C0C0A4F9F89080",
 21799 => x"C0C0C0A4F9F89090",
 21800 => x"C0C0C0A4F980C0C0",
 21801 => x"C0C0C0A4F980C0F9",
 21802 => x"C0C0C0A4F980C0A4",
 21803 => x"C0C0C0A4F980C0B0",
 21804 => x"C0C0C0A4F980C099",
 21805 => x"C0C0C0A4F980C092",
 21806 => x"C0C0C0A4F980C082",
 21807 => x"C0C0C0A4F980C0F8",
 21808 => x"C0C0C0A4F980C080",
 21809 => x"C0C0C0A4F980C090",
 21810 => x"C0C0C0A4F980F9C0",
 21811 => x"C0C0C0A4F980F9F9",
 21812 => x"C0C0C0A4F980F9A4",
 21813 => x"C0C0C0A4F980F9B0",
 21814 => x"C0C0C0A4F980F999",
 21815 => x"C0C0C0A4F980F992",
 21816 => x"C0C0C0A4F980F982",
 21817 => x"C0C0C0A4F980F9F8",
 21818 => x"C0C0C0A4F980F980",
 21819 => x"C0C0C0A4F980F990",
 21820 => x"C0C0C0A4F980A4C0",
 21821 => x"C0C0C0A4F980A4F9",
 21822 => x"C0C0C0A4F980A4A4",
 21823 => x"C0C0C0A4F980A4B0",
 21824 => x"C0C0C0A4F980A499",
 21825 => x"C0C0C0A4F980A492",
 21826 => x"C0C0C0A4F980A482",
 21827 => x"C0C0C0A4F980A4F8",
 21828 => x"C0C0C0A4F980A480",
 21829 => x"C0C0C0A4F980A490",
 21830 => x"C0C0C0A4F980B0C0",
 21831 => x"C0C0C0A4F980B0F9",
 21832 => x"C0C0C0A4F980B0A4",
 21833 => x"C0C0C0A4F980B0B0",
 21834 => x"C0C0C0A4F980B099",
 21835 => x"C0C0C0A4F980B092",
 21836 => x"C0C0C0A4F980B082",
 21837 => x"C0C0C0A4F980B0F8",
 21838 => x"C0C0C0A4F980B080",
 21839 => x"C0C0C0A4F980B090",
 21840 => x"C0C0C0A4F98099C0",
 21841 => x"C0C0C0A4F98099F9",
 21842 => x"C0C0C0A4F98099A4",
 21843 => x"C0C0C0A4F98099B0",
 21844 => x"C0C0C0A4F9809999",
 21845 => x"C0C0C0A4F9809992",
 21846 => x"C0C0C0A4F9809982",
 21847 => x"C0C0C0A4F98099F8",
 21848 => x"C0C0C0A4F9809980",
 21849 => x"C0C0C0A4F9809990",
 21850 => x"C0C0C0A4F98092C0",
 21851 => x"C0C0C0A4F98092F9",
 21852 => x"C0C0C0A4F98092A4",
 21853 => x"C0C0C0A4F98092B0",
 21854 => x"C0C0C0A4F9809299",
 21855 => x"C0C0C0A4F9809292",
 21856 => x"C0C0C0A4F9809282",
 21857 => x"C0C0C0A4F98092F8",
 21858 => x"C0C0C0A4F9809280",
 21859 => x"C0C0C0A4F9809290",
 21860 => x"C0C0C0A4F98082C0",
 21861 => x"C0C0C0A4F98082F9",
 21862 => x"C0C0C0A4F98082A4",
 21863 => x"C0C0C0A4F98082B0",
 21864 => x"C0C0C0A4F9808299",
 21865 => x"C0C0C0A4F9808292",
 21866 => x"C0C0C0A4F9808282",
 21867 => x"C0C0C0A4F98082F8",
 21868 => x"C0C0C0A4F9808280",
 21869 => x"C0C0C0A4F9808290",
 21870 => x"C0C0C0A4F980F8C0",
 21871 => x"C0C0C0A4F980F8F9",
 21872 => x"C0C0C0A4F980F8A4",
 21873 => x"C0C0C0A4F980F8B0",
 21874 => x"C0C0C0A4F980F899",
 21875 => x"C0C0C0A4F980F892",
 21876 => x"C0C0C0A4F980F882",
 21877 => x"C0C0C0A4F980F8F8",
 21878 => x"C0C0C0A4F980F880",
 21879 => x"C0C0C0A4F980F890",
 21880 => x"C0C0C0A4F98080C0",
 21881 => x"C0C0C0A4F98080F9",
 21882 => x"C0C0C0A4F98080A4",
 21883 => x"C0C0C0A4F98080B0",
 21884 => x"C0C0C0A4F9808099",
 21885 => x"C0C0C0A4F9808092",
 21886 => x"C0C0C0A4F9808082",
 21887 => x"C0C0C0A4F98080F8",
 21888 => x"C0C0C0A4F9808080",
 21889 => x"C0C0C0A4F9808090",
 21890 => x"C0C0C0A4F98090C0",
 21891 => x"C0C0C0A4F98090F9",
 21892 => x"C0C0C0A4F98090A4",
 21893 => x"C0C0C0A4F98090B0",
 21894 => x"C0C0C0A4F9809099",
 21895 => x"C0C0C0A4F9809092",
 21896 => x"C0C0C0A4F9809082",
 21897 => x"C0C0C0A4F98090F8",
 21898 => x"C0C0C0A4F9809080",
 21899 => x"C0C0C0A4F9809090",
 21900 => x"C0C0C0A4F990C0C0",
 21901 => x"C0C0C0A4F990C0F9",
 21902 => x"C0C0C0A4F990C0A4",
 21903 => x"C0C0C0A4F990C0B0",
 21904 => x"C0C0C0A4F990C099",
 21905 => x"C0C0C0A4F990C092",
 21906 => x"C0C0C0A4F990C082",
 21907 => x"C0C0C0A4F990C0F8",
 21908 => x"C0C0C0A4F990C080",
 21909 => x"C0C0C0A4F990C090",
 21910 => x"C0C0C0A4F990F9C0",
 21911 => x"C0C0C0A4F990F9F9",
 21912 => x"C0C0C0A4F990F9A4",
 21913 => x"C0C0C0A4F990F9B0",
 21914 => x"C0C0C0A4F990F999",
 21915 => x"C0C0C0A4F990F992",
 21916 => x"C0C0C0A4F990F982",
 21917 => x"C0C0C0A4F990F9F8",
 21918 => x"C0C0C0A4F990F980",
 21919 => x"C0C0C0A4F990F990",
 21920 => x"C0C0C0A4F990A4C0",
 21921 => x"C0C0C0A4F990A4F9",
 21922 => x"C0C0C0A4F990A4A4",
 21923 => x"C0C0C0A4F990A4B0",
 21924 => x"C0C0C0A4F990A499",
 21925 => x"C0C0C0A4F990A492",
 21926 => x"C0C0C0A4F990A482",
 21927 => x"C0C0C0A4F990A4F8",
 21928 => x"C0C0C0A4F990A480",
 21929 => x"C0C0C0A4F990A490",
 21930 => x"C0C0C0A4F990B0C0",
 21931 => x"C0C0C0A4F990B0F9",
 21932 => x"C0C0C0A4F990B0A4",
 21933 => x"C0C0C0A4F990B0B0",
 21934 => x"C0C0C0A4F990B099",
 21935 => x"C0C0C0A4F990B092",
 21936 => x"C0C0C0A4F990B082",
 21937 => x"C0C0C0A4F990B0F8",
 21938 => x"C0C0C0A4F990B080",
 21939 => x"C0C0C0A4F990B090",
 21940 => x"C0C0C0A4F99099C0",
 21941 => x"C0C0C0A4F99099F9",
 21942 => x"C0C0C0A4F99099A4",
 21943 => x"C0C0C0A4F99099B0",
 21944 => x"C0C0C0A4F9909999",
 21945 => x"C0C0C0A4F9909992",
 21946 => x"C0C0C0A4F9909982",
 21947 => x"C0C0C0A4F99099F8",
 21948 => x"C0C0C0A4F9909980",
 21949 => x"C0C0C0A4F9909990",
 21950 => x"C0C0C0A4F99092C0",
 21951 => x"C0C0C0A4F99092F9",
 21952 => x"C0C0C0A4F99092A4",
 21953 => x"C0C0C0A4F99092B0",
 21954 => x"C0C0C0A4F9909299",
 21955 => x"C0C0C0A4F9909292",
 21956 => x"C0C0C0A4F9909282",
 21957 => x"C0C0C0A4F99092F8",
 21958 => x"C0C0C0A4F9909280",
 21959 => x"C0C0C0A4F9909290",
 21960 => x"C0C0C0A4F99082C0",
 21961 => x"C0C0C0A4F99082F9",
 21962 => x"C0C0C0A4F99082A4",
 21963 => x"C0C0C0A4F99082B0",
 21964 => x"C0C0C0A4F9908299",
 21965 => x"C0C0C0A4F9908292",
 21966 => x"C0C0C0A4F9908282",
 21967 => x"C0C0C0A4F99082F8",
 21968 => x"C0C0C0A4F9908280",
 21969 => x"C0C0C0A4F9908290",
 21970 => x"C0C0C0A4F990F8C0",
 21971 => x"C0C0C0A4F990F8F9",
 21972 => x"C0C0C0A4F990F8A4",
 21973 => x"C0C0C0A4F990F8B0",
 21974 => x"C0C0C0A4F990F899",
 21975 => x"C0C0C0A4F990F892",
 21976 => x"C0C0C0A4F990F882",
 21977 => x"C0C0C0A4F990F8F8",
 21978 => x"C0C0C0A4F990F880",
 21979 => x"C0C0C0A4F990F890",
 21980 => x"C0C0C0A4F99080C0",
 21981 => x"C0C0C0A4F99080F9",
 21982 => x"C0C0C0A4F99080A4",
 21983 => x"C0C0C0A4F99080B0",
 21984 => x"C0C0C0A4F9908099",
 21985 => x"C0C0C0A4F9908092",
 21986 => x"C0C0C0A4F9908082",
 21987 => x"C0C0C0A4F99080F8",
 21988 => x"C0C0C0A4F9908080",
 21989 => x"C0C0C0A4F9908090",
 21990 => x"C0C0C0A4F99090C0",
 21991 => x"C0C0C0A4F99090F9",
 21992 => x"C0C0C0A4F99090A4",
 21993 => x"C0C0C0A4F99090B0",
 21994 => x"C0C0C0A4F9909099",
 21995 => x"C0C0C0A4F9909092",
 21996 => x"C0C0C0A4F9909082",
 21997 => x"C0C0C0A4F99090F8",
 21998 => x"C0C0C0A4F9909080",
 21999 => x"C0C0C0A4F9909090",
 22000 => x"C0C0C0A4A4C0C0C0",
 22001 => x"C0C0C0A4A4C0C0F9",
 22002 => x"C0C0C0A4A4C0C0A4",
 22003 => x"C0C0C0A4A4C0C0B0",
 22004 => x"C0C0C0A4A4C0C099",
 22005 => x"C0C0C0A4A4C0C092",
 22006 => x"C0C0C0A4A4C0C082",
 22007 => x"C0C0C0A4A4C0C0F8",
 22008 => x"C0C0C0A4A4C0C080",
 22009 => x"C0C0C0A4A4C0C090",
 22010 => x"C0C0C0A4A4C0F9C0",
 22011 => x"C0C0C0A4A4C0F9F9",
 22012 => x"C0C0C0A4A4C0F9A4",
 22013 => x"C0C0C0A4A4C0F9B0",
 22014 => x"C0C0C0A4A4C0F999",
 22015 => x"C0C0C0A4A4C0F992",
 22016 => x"C0C0C0A4A4C0F982",
 22017 => x"C0C0C0A4A4C0F9F8",
 22018 => x"C0C0C0A4A4C0F980",
 22019 => x"C0C0C0A4A4C0F990",
 22020 => x"C0C0C0A4A4C0A4C0",
 22021 => x"C0C0C0A4A4C0A4F9",
 22022 => x"C0C0C0A4A4C0A4A4",
 22023 => x"C0C0C0A4A4C0A4B0",
 22024 => x"C0C0C0A4A4C0A499",
 22025 => x"C0C0C0A4A4C0A492",
 22026 => x"C0C0C0A4A4C0A482",
 22027 => x"C0C0C0A4A4C0A4F8",
 22028 => x"C0C0C0A4A4C0A480",
 22029 => x"C0C0C0A4A4C0A490",
 22030 => x"C0C0C0A4A4C0B0C0",
 22031 => x"C0C0C0A4A4C0B0F9",
 22032 => x"C0C0C0A4A4C0B0A4",
 22033 => x"C0C0C0A4A4C0B0B0",
 22034 => x"C0C0C0A4A4C0B099",
 22035 => x"C0C0C0A4A4C0B092",
 22036 => x"C0C0C0A4A4C0B082",
 22037 => x"C0C0C0A4A4C0B0F8",
 22038 => x"C0C0C0A4A4C0B080",
 22039 => x"C0C0C0A4A4C0B090",
 22040 => x"C0C0C0A4A4C099C0",
 22041 => x"C0C0C0A4A4C099F9",
 22042 => x"C0C0C0A4A4C099A4",
 22043 => x"C0C0C0A4A4C099B0",
 22044 => x"C0C0C0A4A4C09999",
 22045 => x"C0C0C0A4A4C09992",
 22046 => x"C0C0C0A4A4C09982",
 22047 => x"C0C0C0A4A4C099F8",
 22048 => x"C0C0C0A4A4C09980",
 22049 => x"C0C0C0A4A4C09990",
 22050 => x"C0C0C0A4A4C092C0",
 22051 => x"C0C0C0A4A4C092F9",
 22052 => x"C0C0C0A4A4C092A4",
 22053 => x"C0C0C0A4A4C092B0",
 22054 => x"C0C0C0A4A4C09299",
 22055 => x"C0C0C0A4A4C09292",
 22056 => x"C0C0C0A4A4C09282",
 22057 => x"C0C0C0A4A4C092F8",
 22058 => x"C0C0C0A4A4C09280",
 22059 => x"C0C0C0A4A4C09290",
 22060 => x"C0C0C0A4A4C082C0",
 22061 => x"C0C0C0A4A4C082F9",
 22062 => x"C0C0C0A4A4C082A4",
 22063 => x"C0C0C0A4A4C082B0",
 22064 => x"C0C0C0A4A4C08299",
 22065 => x"C0C0C0A4A4C08292",
 22066 => x"C0C0C0A4A4C08282",
 22067 => x"C0C0C0A4A4C082F8",
 22068 => x"C0C0C0A4A4C08280",
 22069 => x"C0C0C0A4A4C08290",
 22070 => x"C0C0C0A4A4C0F8C0",
 22071 => x"C0C0C0A4A4C0F8F9",
 22072 => x"C0C0C0A4A4C0F8A4",
 22073 => x"C0C0C0A4A4C0F8B0",
 22074 => x"C0C0C0A4A4C0F899",
 22075 => x"C0C0C0A4A4C0F892",
 22076 => x"C0C0C0A4A4C0F882",
 22077 => x"C0C0C0A4A4C0F8F8",
 22078 => x"C0C0C0A4A4C0F880",
 22079 => x"C0C0C0A4A4C0F890",
 22080 => x"C0C0C0A4A4C080C0",
 22081 => x"C0C0C0A4A4C080F9",
 22082 => x"C0C0C0A4A4C080A4",
 22083 => x"C0C0C0A4A4C080B0",
 22084 => x"C0C0C0A4A4C08099",
 22085 => x"C0C0C0A4A4C08092",
 22086 => x"C0C0C0A4A4C08082",
 22087 => x"C0C0C0A4A4C080F8",
 22088 => x"C0C0C0A4A4C08080",
 22089 => x"C0C0C0A4A4C08090",
 22090 => x"C0C0C0A4A4C090C0",
 22091 => x"C0C0C0A4A4C090F9",
 22092 => x"C0C0C0A4A4C090A4",
 22093 => x"C0C0C0A4A4C090B0",
 22094 => x"C0C0C0A4A4C09099",
 22095 => x"C0C0C0A4A4C09092",
 22096 => x"C0C0C0A4A4C09082",
 22097 => x"C0C0C0A4A4C090F8",
 22098 => x"C0C0C0A4A4C09080",
 22099 => x"C0C0C0A4A4C09090",
 22100 => x"C0C0C0A4A4F9C0C0",
 22101 => x"C0C0C0A4A4F9C0F9",
 22102 => x"C0C0C0A4A4F9C0A4",
 22103 => x"C0C0C0A4A4F9C0B0",
 22104 => x"C0C0C0A4A4F9C099",
 22105 => x"C0C0C0A4A4F9C092",
 22106 => x"C0C0C0A4A4F9C082",
 22107 => x"C0C0C0A4A4F9C0F8",
 22108 => x"C0C0C0A4A4F9C080",
 22109 => x"C0C0C0A4A4F9C090",
 22110 => x"C0C0C0A4A4F9F9C0",
 22111 => x"C0C0C0A4A4F9F9F9",
 22112 => x"C0C0C0A4A4F9F9A4",
 22113 => x"C0C0C0A4A4F9F9B0",
 22114 => x"C0C0C0A4A4F9F999",
 22115 => x"C0C0C0A4A4F9F992",
 22116 => x"C0C0C0A4A4F9F982",
 22117 => x"C0C0C0A4A4F9F9F8",
 22118 => x"C0C0C0A4A4F9F980",
 22119 => x"C0C0C0A4A4F9F990",
 22120 => x"C0C0C0A4A4F9A4C0",
 22121 => x"C0C0C0A4A4F9A4F9",
 22122 => x"C0C0C0A4A4F9A4A4",
 22123 => x"C0C0C0A4A4F9A4B0",
 22124 => x"C0C0C0A4A4F9A499",
 22125 => x"C0C0C0A4A4F9A492",
 22126 => x"C0C0C0A4A4F9A482",
 22127 => x"C0C0C0A4A4F9A4F8",
 22128 => x"C0C0C0A4A4F9A480",
 22129 => x"C0C0C0A4A4F9A490",
 22130 => x"C0C0C0A4A4F9B0C0",
 22131 => x"C0C0C0A4A4F9B0F9",
 22132 => x"C0C0C0A4A4F9B0A4",
 22133 => x"C0C0C0A4A4F9B0B0",
 22134 => x"C0C0C0A4A4F9B099",
 22135 => x"C0C0C0A4A4F9B092",
 22136 => x"C0C0C0A4A4F9B082",
 22137 => x"C0C0C0A4A4F9B0F8",
 22138 => x"C0C0C0A4A4F9B080",
 22139 => x"C0C0C0A4A4F9B090",
 22140 => x"C0C0C0A4A4F999C0",
 22141 => x"C0C0C0A4A4F999F9",
 22142 => x"C0C0C0A4A4F999A4",
 22143 => x"C0C0C0A4A4F999B0",
 22144 => x"C0C0C0A4A4F99999",
 22145 => x"C0C0C0A4A4F99992",
 22146 => x"C0C0C0A4A4F99982",
 22147 => x"C0C0C0A4A4F999F8",
 22148 => x"C0C0C0A4A4F99980",
 22149 => x"C0C0C0A4A4F99990",
 22150 => x"C0C0C0A4A4F992C0",
 22151 => x"C0C0C0A4A4F992F9",
 22152 => x"C0C0C0A4A4F992A4",
 22153 => x"C0C0C0A4A4F992B0",
 22154 => x"C0C0C0A4A4F99299",
 22155 => x"C0C0C0A4A4F99292",
 22156 => x"C0C0C0A4A4F99282",
 22157 => x"C0C0C0A4A4F992F8",
 22158 => x"C0C0C0A4A4F99280",
 22159 => x"C0C0C0A4A4F99290",
 22160 => x"C0C0C0A4A4F982C0",
 22161 => x"C0C0C0A4A4F982F9",
 22162 => x"C0C0C0A4A4F982A4",
 22163 => x"C0C0C0A4A4F982B0",
 22164 => x"C0C0C0A4A4F98299",
 22165 => x"C0C0C0A4A4F98292",
 22166 => x"C0C0C0A4A4F98282",
 22167 => x"C0C0C0A4A4F982F8",
 22168 => x"C0C0C0A4A4F98280",
 22169 => x"C0C0C0A4A4F98290",
 22170 => x"C0C0C0A4A4F9F8C0",
 22171 => x"C0C0C0A4A4F9F8F9",
 22172 => x"C0C0C0A4A4F9F8A4",
 22173 => x"C0C0C0A4A4F9F8B0",
 22174 => x"C0C0C0A4A4F9F899",
 22175 => x"C0C0C0A4A4F9F892",
 22176 => x"C0C0C0A4A4F9F882",
 22177 => x"C0C0C0A4A4F9F8F8",
 22178 => x"C0C0C0A4A4F9F880",
 22179 => x"C0C0C0A4A4F9F890",
 22180 => x"C0C0C0A4A4F980C0",
 22181 => x"C0C0C0A4A4F980F9",
 22182 => x"C0C0C0A4A4F980A4",
 22183 => x"C0C0C0A4A4F980B0",
 22184 => x"C0C0C0A4A4F98099",
 22185 => x"C0C0C0A4A4F98092",
 22186 => x"C0C0C0A4A4F98082",
 22187 => x"C0C0C0A4A4F980F8",
 22188 => x"C0C0C0A4A4F98080",
 22189 => x"C0C0C0A4A4F98090",
 22190 => x"C0C0C0A4A4F990C0",
 22191 => x"C0C0C0A4A4F990F9",
 22192 => x"C0C0C0A4A4F990A4",
 22193 => x"C0C0C0A4A4F990B0",
 22194 => x"C0C0C0A4A4F99099",
 22195 => x"C0C0C0A4A4F99092",
 22196 => x"C0C0C0A4A4F99082",
 22197 => x"C0C0C0A4A4F990F8",
 22198 => x"C0C0C0A4A4F99080",
 22199 => x"C0C0C0A4A4F99090",
 22200 => x"C0C0C0A4A4A4C0C0",
 22201 => x"C0C0C0A4A4A4C0F9",
 22202 => x"C0C0C0A4A4A4C0A4",
 22203 => x"C0C0C0A4A4A4C0B0",
 22204 => x"C0C0C0A4A4A4C099",
 22205 => x"C0C0C0A4A4A4C092",
 22206 => x"C0C0C0A4A4A4C082",
 22207 => x"C0C0C0A4A4A4C0F8",
 22208 => x"C0C0C0A4A4A4C080",
 22209 => x"C0C0C0A4A4A4C090",
 22210 => x"C0C0C0A4A4A4F9C0",
 22211 => x"C0C0C0A4A4A4F9F9",
 22212 => x"C0C0C0A4A4A4F9A4",
 22213 => x"C0C0C0A4A4A4F9B0",
 22214 => x"C0C0C0A4A4A4F999",
 22215 => x"C0C0C0A4A4A4F992",
 22216 => x"C0C0C0A4A4A4F982",
 22217 => x"C0C0C0A4A4A4F9F8",
 22218 => x"C0C0C0A4A4A4F980",
 22219 => x"C0C0C0A4A4A4F990",
 22220 => x"C0C0C0A4A4A4A4C0",
 22221 => x"C0C0C0A4A4A4A4F9",
 22222 => x"C0C0C0A4A4A4A4A4",
 22223 => x"C0C0C0A4A4A4A4B0",
 22224 => x"C0C0C0A4A4A4A499",
 22225 => x"C0C0C0A4A4A4A492",
 22226 => x"C0C0C0A4A4A4A482",
 22227 => x"C0C0C0A4A4A4A4F8",
 22228 => x"C0C0C0A4A4A4A480",
 22229 => x"C0C0C0A4A4A4A490",
 22230 => x"C0C0C0A4A4A4B0C0",
 22231 => x"C0C0C0A4A4A4B0F9",
 22232 => x"C0C0C0A4A4A4B0A4",
 22233 => x"C0C0C0A4A4A4B0B0",
 22234 => x"C0C0C0A4A4A4B099",
 22235 => x"C0C0C0A4A4A4B092",
 22236 => x"C0C0C0A4A4A4B082",
 22237 => x"C0C0C0A4A4A4B0F8",
 22238 => x"C0C0C0A4A4A4B080",
 22239 => x"C0C0C0A4A4A4B090",
 22240 => x"C0C0C0A4A4A499C0",
 22241 => x"C0C0C0A4A4A499F9",
 22242 => x"C0C0C0A4A4A499A4",
 22243 => x"C0C0C0A4A4A499B0",
 22244 => x"C0C0C0A4A4A49999",
 22245 => x"C0C0C0A4A4A49992",
 22246 => x"C0C0C0A4A4A49982",
 22247 => x"C0C0C0A4A4A499F8",
 22248 => x"C0C0C0A4A4A49980",
 22249 => x"C0C0C0A4A4A49990",
 22250 => x"C0C0C0A4A4A492C0",
 22251 => x"C0C0C0A4A4A492F9",
 22252 => x"C0C0C0A4A4A492A4",
 22253 => x"C0C0C0A4A4A492B0",
 22254 => x"C0C0C0A4A4A49299",
 22255 => x"C0C0C0A4A4A49292",
 22256 => x"C0C0C0A4A4A49282",
 22257 => x"C0C0C0A4A4A492F8",
 22258 => x"C0C0C0A4A4A49280",
 22259 => x"C0C0C0A4A4A49290",
 22260 => x"C0C0C0A4A4A482C0",
 22261 => x"C0C0C0A4A4A482F9",
 22262 => x"C0C0C0A4A4A482A4",
 22263 => x"C0C0C0A4A4A482B0",
 22264 => x"C0C0C0A4A4A48299",
 22265 => x"C0C0C0A4A4A48292",
 22266 => x"C0C0C0A4A4A48282",
 22267 => x"C0C0C0A4A4A482F8",
 22268 => x"C0C0C0A4A4A48280",
 22269 => x"C0C0C0A4A4A48290",
 22270 => x"C0C0C0A4A4A4F8C0",
 22271 => x"C0C0C0A4A4A4F8F9",
 22272 => x"C0C0C0A4A4A4F8A4",
 22273 => x"C0C0C0A4A4A4F8B0",
 22274 => x"C0C0C0A4A4A4F899",
 22275 => x"C0C0C0A4A4A4F892",
 22276 => x"C0C0C0A4A4A4F882",
 22277 => x"C0C0C0A4A4A4F8F8",
 22278 => x"C0C0C0A4A4A4F880",
 22279 => x"C0C0C0A4A4A4F890",
 22280 => x"C0C0C0A4A4A480C0",
 22281 => x"C0C0C0A4A4A480F9",
 22282 => x"C0C0C0A4A4A480A4",
 22283 => x"C0C0C0A4A4A480B0",
 22284 => x"C0C0C0A4A4A48099",
 22285 => x"C0C0C0A4A4A48092",
 22286 => x"C0C0C0A4A4A48082",
 22287 => x"C0C0C0A4A4A480F8",
 22288 => x"C0C0C0A4A4A48080",
 22289 => x"C0C0C0A4A4A48090",
 22290 => x"C0C0C0A4A4A490C0",
 22291 => x"C0C0C0A4A4A490F9",
 22292 => x"C0C0C0A4A4A490A4",
 22293 => x"C0C0C0A4A4A490B0",
 22294 => x"C0C0C0A4A4A49099",
 22295 => x"C0C0C0A4A4A49092",
 22296 => x"C0C0C0A4A4A49082",
 22297 => x"C0C0C0A4A4A490F8",
 22298 => x"C0C0C0A4A4A49080",
 22299 => x"C0C0C0A4A4A49090",
 22300 => x"C0C0C0A4A4B0C0C0",
 22301 => x"C0C0C0A4A4B0C0F9",
 22302 => x"C0C0C0A4A4B0C0A4",
 22303 => x"C0C0C0A4A4B0C0B0",
 22304 => x"C0C0C0A4A4B0C099",
 22305 => x"C0C0C0A4A4B0C092",
 22306 => x"C0C0C0A4A4B0C082",
 22307 => x"C0C0C0A4A4B0C0F8",
 22308 => x"C0C0C0A4A4B0C080",
 22309 => x"C0C0C0A4A4B0C090",
 22310 => x"C0C0C0A4A4B0F9C0",
 22311 => x"C0C0C0A4A4B0F9F9",
 22312 => x"C0C0C0A4A4B0F9A4",
 22313 => x"C0C0C0A4A4B0F9B0",
 22314 => x"C0C0C0A4A4B0F999",
 22315 => x"C0C0C0A4A4B0F992",
 22316 => x"C0C0C0A4A4B0F982",
 22317 => x"C0C0C0A4A4B0F9F8",
 22318 => x"C0C0C0A4A4B0F980",
 22319 => x"C0C0C0A4A4B0F990",
 22320 => x"C0C0C0A4A4B0A4C0",
 22321 => x"C0C0C0A4A4B0A4F9",
 22322 => x"C0C0C0A4A4B0A4A4",
 22323 => x"C0C0C0A4A4B0A4B0",
 22324 => x"C0C0C0A4A4B0A499",
 22325 => x"C0C0C0A4A4B0A492",
 22326 => x"C0C0C0A4A4B0A482",
 22327 => x"C0C0C0A4A4B0A4F8",
 22328 => x"C0C0C0A4A4B0A480",
 22329 => x"C0C0C0A4A4B0A490",
 22330 => x"C0C0C0A4A4B0B0C0",
 22331 => x"C0C0C0A4A4B0B0F9",
 22332 => x"C0C0C0A4A4B0B0A4",
 22333 => x"C0C0C0A4A4B0B0B0",
 22334 => x"C0C0C0A4A4B0B099",
 22335 => x"C0C0C0A4A4B0B092",
 22336 => x"C0C0C0A4A4B0B082",
 22337 => x"C0C0C0A4A4B0B0F8",
 22338 => x"C0C0C0A4A4B0B080",
 22339 => x"C0C0C0A4A4B0B090",
 22340 => x"C0C0C0A4A4B099C0",
 22341 => x"C0C0C0A4A4B099F9",
 22342 => x"C0C0C0A4A4B099A4",
 22343 => x"C0C0C0A4A4B099B0",
 22344 => x"C0C0C0A4A4B09999",
 22345 => x"C0C0C0A4A4B09992",
 22346 => x"C0C0C0A4A4B09982",
 22347 => x"C0C0C0A4A4B099F8",
 22348 => x"C0C0C0A4A4B09980",
 22349 => x"C0C0C0A4A4B09990",
 22350 => x"C0C0C0A4A4B092C0",
 22351 => x"C0C0C0A4A4B092F9",
 22352 => x"C0C0C0A4A4B092A4",
 22353 => x"C0C0C0A4A4B092B0",
 22354 => x"C0C0C0A4A4B09299",
 22355 => x"C0C0C0A4A4B09292",
 22356 => x"C0C0C0A4A4B09282",
 22357 => x"C0C0C0A4A4B092F8",
 22358 => x"C0C0C0A4A4B09280",
 22359 => x"C0C0C0A4A4B09290",
 22360 => x"C0C0C0A4A4B082C0",
 22361 => x"C0C0C0A4A4B082F9",
 22362 => x"C0C0C0A4A4B082A4",
 22363 => x"C0C0C0A4A4B082B0",
 22364 => x"C0C0C0A4A4B08299",
 22365 => x"C0C0C0A4A4B08292",
 22366 => x"C0C0C0A4A4B08282",
 22367 => x"C0C0C0A4A4B082F8",
 22368 => x"C0C0C0A4A4B08280",
 22369 => x"C0C0C0A4A4B08290",
 22370 => x"C0C0C0A4A4B0F8C0",
 22371 => x"C0C0C0A4A4B0F8F9",
 22372 => x"C0C0C0A4A4B0F8A4",
 22373 => x"C0C0C0A4A4B0F8B0",
 22374 => x"C0C0C0A4A4B0F899",
 22375 => x"C0C0C0A4A4B0F892",
 22376 => x"C0C0C0A4A4B0F882",
 22377 => x"C0C0C0A4A4B0F8F8",
 22378 => x"C0C0C0A4A4B0F880",
 22379 => x"C0C0C0A4A4B0F890",
 22380 => x"C0C0C0A4A4B080C0",
 22381 => x"C0C0C0A4A4B080F9",
 22382 => x"C0C0C0A4A4B080A4",
 22383 => x"C0C0C0A4A4B080B0",
 22384 => x"C0C0C0A4A4B08099",
 22385 => x"C0C0C0A4A4B08092",
 22386 => x"C0C0C0A4A4B08082",
 22387 => x"C0C0C0A4A4B080F8",
 22388 => x"C0C0C0A4A4B08080",
 22389 => x"C0C0C0A4A4B08090",
 22390 => x"C0C0C0A4A4B090C0",
 22391 => x"C0C0C0A4A4B090F9",
 22392 => x"C0C0C0A4A4B090A4",
 22393 => x"C0C0C0A4A4B090B0",
 22394 => x"C0C0C0A4A4B09099",
 22395 => x"C0C0C0A4A4B09092",
 22396 => x"C0C0C0A4A4B09082",
 22397 => x"C0C0C0A4A4B090F8",
 22398 => x"C0C0C0A4A4B09080",
 22399 => x"C0C0C0A4A4B09090",
 22400 => x"C0C0C0A4A499C0C0",
 22401 => x"C0C0C0A4A499C0F9",
 22402 => x"C0C0C0A4A499C0A4",
 22403 => x"C0C0C0A4A499C0B0",
 22404 => x"C0C0C0A4A499C099",
 22405 => x"C0C0C0A4A499C092",
 22406 => x"C0C0C0A4A499C082",
 22407 => x"C0C0C0A4A499C0F8",
 22408 => x"C0C0C0A4A499C080",
 22409 => x"C0C0C0A4A499C090",
 22410 => x"C0C0C0A4A499F9C0",
 22411 => x"C0C0C0A4A499F9F9",
 22412 => x"C0C0C0A4A499F9A4",
 22413 => x"C0C0C0A4A499F9B0",
 22414 => x"C0C0C0A4A499F999",
 22415 => x"C0C0C0A4A499F992",
 22416 => x"C0C0C0A4A499F982",
 22417 => x"C0C0C0A4A499F9F8",
 22418 => x"C0C0C0A4A499F980",
 22419 => x"C0C0C0A4A499F990",
 22420 => x"C0C0C0A4A499A4C0",
 22421 => x"C0C0C0A4A499A4F9",
 22422 => x"C0C0C0A4A499A4A4",
 22423 => x"C0C0C0A4A499A4B0",
 22424 => x"C0C0C0A4A499A499",
 22425 => x"C0C0C0A4A499A492",
 22426 => x"C0C0C0A4A499A482",
 22427 => x"C0C0C0A4A499A4F8",
 22428 => x"C0C0C0A4A499A480",
 22429 => x"C0C0C0A4A499A490",
 22430 => x"C0C0C0A4A499B0C0",
 22431 => x"C0C0C0A4A499B0F9",
 22432 => x"C0C0C0A4A499B0A4",
 22433 => x"C0C0C0A4A499B0B0",
 22434 => x"C0C0C0A4A499B099",
 22435 => x"C0C0C0A4A499B092",
 22436 => x"C0C0C0A4A499B082",
 22437 => x"C0C0C0A4A499B0F8",
 22438 => x"C0C0C0A4A499B080",
 22439 => x"C0C0C0A4A499B090",
 22440 => x"C0C0C0A4A49999C0",
 22441 => x"C0C0C0A4A49999F9",
 22442 => x"C0C0C0A4A49999A4",
 22443 => x"C0C0C0A4A49999B0",
 22444 => x"C0C0C0A4A4999999",
 22445 => x"C0C0C0A4A4999992",
 22446 => x"C0C0C0A4A4999982",
 22447 => x"C0C0C0A4A49999F8",
 22448 => x"C0C0C0A4A4999980",
 22449 => x"C0C0C0A4A4999990",
 22450 => x"C0C0C0A4A49992C0",
 22451 => x"C0C0C0A4A49992F9",
 22452 => x"C0C0C0A4A49992A4",
 22453 => x"C0C0C0A4A49992B0",
 22454 => x"C0C0C0A4A4999299",
 22455 => x"C0C0C0A4A4999292",
 22456 => x"C0C0C0A4A4999282",
 22457 => x"C0C0C0A4A49992F8",
 22458 => x"C0C0C0A4A4999280",
 22459 => x"C0C0C0A4A4999290",
 22460 => x"C0C0C0A4A49982C0",
 22461 => x"C0C0C0A4A49982F9",
 22462 => x"C0C0C0A4A49982A4",
 22463 => x"C0C0C0A4A49982B0",
 22464 => x"C0C0C0A4A4998299",
 22465 => x"C0C0C0A4A4998292",
 22466 => x"C0C0C0A4A4998282",
 22467 => x"C0C0C0A4A49982F8",
 22468 => x"C0C0C0A4A4998280",
 22469 => x"C0C0C0A4A4998290",
 22470 => x"C0C0C0A4A499F8C0",
 22471 => x"C0C0C0A4A499F8F9",
 22472 => x"C0C0C0A4A499F8A4",
 22473 => x"C0C0C0A4A499F8B0",
 22474 => x"C0C0C0A4A499F899",
 22475 => x"C0C0C0A4A499F892",
 22476 => x"C0C0C0A4A499F882",
 22477 => x"C0C0C0A4A499F8F8",
 22478 => x"C0C0C0A4A499F880",
 22479 => x"C0C0C0A4A499F890",
 22480 => x"C0C0C0A4A49980C0",
 22481 => x"C0C0C0A4A49980F9",
 22482 => x"C0C0C0A4A49980A4",
 22483 => x"C0C0C0A4A49980B0",
 22484 => x"C0C0C0A4A4998099",
 22485 => x"C0C0C0A4A4998092",
 22486 => x"C0C0C0A4A4998082",
 22487 => x"C0C0C0A4A49980F8",
 22488 => x"C0C0C0A4A4998080",
 22489 => x"C0C0C0A4A4998090",
 22490 => x"C0C0C0A4A49990C0",
 22491 => x"C0C0C0A4A49990F9",
 22492 => x"C0C0C0A4A49990A4",
 22493 => x"C0C0C0A4A49990B0",
 22494 => x"C0C0C0A4A4999099",
 22495 => x"C0C0C0A4A4999092",
 22496 => x"C0C0C0A4A4999082",
 22497 => x"C0C0C0A4A49990F8",
 22498 => x"C0C0C0A4A4999080",
 22499 => x"C0C0C0A4A4999090",
 22500 => x"C0C0C0A4A492C0C0",
 22501 => x"C0C0C0A4A492C0F9",
 22502 => x"C0C0C0A4A492C0A4",
 22503 => x"C0C0C0A4A492C0B0",
 22504 => x"C0C0C0A4A492C099",
 22505 => x"C0C0C0A4A492C092",
 22506 => x"C0C0C0A4A492C082",
 22507 => x"C0C0C0A4A492C0F8",
 22508 => x"C0C0C0A4A492C080",
 22509 => x"C0C0C0A4A492C090",
 22510 => x"C0C0C0A4A492F9C0",
 22511 => x"C0C0C0A4A492F9F9",
 22512 => x"C0C0C0A4A492F9A4",
 22513 => x"C0C0C0A4A492F9B0",
 22514 => x"C0C0C0A4A492F999",
 22515 => x"C0C0C0A4A492F992",
 22516 => x"C0C0C0A4A492F982",
 22517 => x"C0C0C0A4A492F9F8",
 22518 => x"C0C0C0A4A492F980",
 22519 => x"C0C0C0A4A492F990",
 22520 => x"C0C0C0A4A492A4C0",
 22521 => x"C0C0C0A4A492A4F9",
 22522 => x"C0C0C0A4A492A4A4",
 22523 => x"C0C0C0A4A492A4B0",
 22524 => x"C0C0C0A4A492A499",
 22525 => x"C0C0C0A4A492A492",
 22526 => x"C0C0C0A4A492A482",
 22527 => x"C0C0C0A4A492A4F8",
 22528 => x"C0C0C0A4A492A480",
 22529 => x"C0C0C0A4A492A490",
 22530 => x"C0C0C0A4A492B0C0",
 22531 => x"C0C0C0A4A492B0F9",
 22532 => x"C0C0C0A4A492B0A4",
 22533 => x"C0C0C0A4A492B0B0",
 22534 => x"C0C0C0A4A492B099",
 22535 => x"C0C0C0A4A492B092",
 22536 => x"C0C0C0A4A492B082",
 22537 => x"C0C0C0A4A492B0F8",
 22538 => x"C0C0C0A4A492B080",
 22539 => x"C0C0C0A4A492B090",
 22540 => x"C0C0C0A4A49299C0",
 22541 => x"C0C0C0A4A49299F9",
 22542 => x"C0C0C0A4A49299A4",
 22543 => x"C0C0C0A4A49299B0",
 22544 => x"C0C0C0A4A4929999",
 22545 => x"C0C0C0A4A4929992",
 22546 => x"C0C0C0A4A4929982",
 22547 => x"C0C0C0A4A49299F8",
 22548 => x"C0C0C0A4A4929980",
 22549 => x"C0C0C0A4A4929990",
 22550 => x"C0C0C0A4A49292C0",
 22551 => x"C0C0C0A4A49292F9",
 22552 => x"C0C0C0A4A49292A4",
 22553 => x"C0C0C0A4A49292B0",
 22554 => x"C0C0C0A4A4929299",
 22555 => x"C0C0C0A4A4929292",
 22556 => x"C0C0C0A4A4929282",
 22557 => x"C0C0C0A4A49292F8",
 22558 => x"C0C0C0A4A4929280",
 22559 => x"C0C0C0A4A4929290",
 22560 => x"C0C0C0A4A49282C0",
 22561 => x"C0C0C0A4A49282F9",
 22562 => x"C0C0C0A4A49282A4",
 22563 => x"C0C0C0A4A49282B0",
 22564 => x"C0C0C0A4A4928299",
 22565 => x"C0C0C0A4A4928292",
 22566 => x"C0C0C0A4A4928282",
 22567 => x"C0C0C0A4A49282F8",
 22568 => x"C0C0C0A4A4928280",
 22569 => x"C0C0C0A4A4928290",
 22570 => x"C0C0C0A4A492F8C0",
 22571 => x"C0C0C0A4A492F8F9",
 22572 => x"C0C0C0A4A492F8A4",
 22573 => x"C0C0C0A4A492F8B0",
 22574 => x"C0C0C0A4A492F899",
 22575 => x"C0C0C0A4A492F892",
 22576 => x"C0C0C0A4A492F882",
 22577 => x"C0C0C0A4A492F8F8",
 22578 => x"C0C0C0A4A492F880",
 22579 => x"C0C0C0A4A492F890",
 22580 => x"C0C0C0A4A49280C0",
 22581 => x"C0C0C0A4A49280F9",
 22582 => x"C0C0C0A4A49280A4",
 22583 => x"C0C0C0A4A49280B0",
 22584 => x"C0C0C0A4A4928099",
 22585 => x"C0C0C0A4A4928092",
 22586 => x"C0C0C0A4A4928082",
 22587 => x"C0C0C0A4A49280F8",
 22588 => x"C0C0C0A4A4928080",
 22589 => x"C0C0C0A4A4928090",
 22590 => x"C0C0C0A4A49290C0",
 22591 => x"C0C0C0A4A49290F9",
 22592 => x"C0C0C0A4A49290A4",
 22593 => x"C0C0C0A4A49290B0",
 22594 => x"C0C0C0A4A4929099",
 22595 => x"C0C0C0A4A4929092",
 22596 => x"C0C0C0A4A4929082",
 22597 => x"C0C0C0A4A49290F8",
 22598 => x"C0C0C0A4A4929080",
 22599 => x"C0C0C0A4A4929090",
 22600 => x"C0C0C0A4A482C0C0",
 22601 => x"C0C0C0A4A482C0F9",
 22602 => x"C0C0C0A4A482C0A4",
 22603 => x"C0C0C0A4A482C0B0",
 22604 => x"C0C0C0A4A482C099",
 22605 => x"C0C0C0A4A482C092",
 22606 => x"C0C0C0A4A482C082",
 22607 => x"C0C0C0A4A482C0F8",
 22608 => x"C0C0C0A4A482C080",
 22609 => x"C0C0C0A4A482C090",
 22610 => x"C0C0C0A4A482F9C0",
 22611 => x"C0C0C0A4A482F9F9",
 22612 => x"C0C0C0A4A482F9A4",
 22613 => x"C0C0C0A4A482F9B0",
 22614 => x"C0C0C0A4A482F999",
 22615 => x"C0C0C0A4A482F992",
 22616 => x"C0C0C0A4A482F982",
 22617 => x"C0C0C0A4A482F9F8",
 22618 => x"C0C0C0A4A482F980",
 22619 => x"C0C0C0A4A482F990",
 22620 => x"C0C0C0A4A482A4C0",
 22621 => x"C0C0C0A4A482A4F9",
 22622 => x"C0C0C0A4A482A4A4",
 22623 => x"C0C0C0A4A482A4B0",
 22624 => x"C0C0C0A4A482A499",
 22625 => x"C0C0C0A4A482A492",
 22626 => x"C0C0C0A4A482A482",
 22627 => x"C0C0C0A4A482A4F8",
 22628 => x"C0C0C0A4A482A480",
 22629 => x"C0C0C0A4A482A490",
 22630 => x"C0C0C0A4A482B0C0",
 22631 => x"C0C0C0A4A482B0F9",
 22632 => x"C0C0C0A4A482B0A4",
 22633 => x"C0C0C0A4A482B0B0",
 22634 => x"C0C0C0A4A482B099",
 22635 => x"C0C0C0A4A482B092",
 22636 => x"C0C0C0A4A482B082",
 22637 => x"C0C0C0A4A482B0F8",
 22638 => x"C0C0C0A4A482B080",
 22639 => x"C0C0C0A4A482B090",
 22640 => x"C0C0C0A4A48299C0",
 22641 => x"C0C0C0A4A48299F9",
 22642 => x"C0C0C0A4A48299A4",
 22643 => x"C0C0C0A4A48299B0",
 22644 => x"C0C0C0A4A4829999",
 22645 => x"C0C0C0A4A4829992",
 22646 => x"C0C0C0A4A4829982",
 22647 => x"C0C0C0A4A48299F8",
 22648 => x"C0C0C0A4A4829980",
 22649 => x"C0C0C0A4A4829990",
 22650 => x"C0C0C0A4A48292C0",
 22651 => x"C0C0C0A4A48292F9",
 22652 => x"C0C0C0A4A48292A4",
 22653 => x"C0C0C0A4A48292B0",
 22654 => x"C0C0C0A4A4829299",
 22655 => x"C0C0C0A4A4829292",
 22656 => x"C0C0C0A4A4829282",
 22657 => x"C0C0C0A4A48292F8",
 22658 => x"C0C0C0A4A4829280",
 22659 => x"C0C0C0A4A4829290",
 22660 => x"C0C0C0A4A48282C0",
 22661 => x"C0C0C0A4A48282F9",
 22662 => x"C0C0C0A4A48282A4",
 22663 => x"C0C0C0A4A48282B0",
 22664 => x"C0C0C0A4A4828299",
 22665 => x"C0C0C0A4A4828292",
 22666 => x"C0C0C0A4A4828282",
 22667 => x"C0C0C0A4A48282F8",
 22668 => x"C0C0C0A4A4828280",
 22669 => x"C0C0C0A4A4828290",
 22670 => x"C0C0C0A4A482F8C0",
 22671 => x"C0C0C0A4A482F8F9",
 22672 => x"C0C0C0A4A482F8A4",
 22673 => x"C0C0C0A4A482F8B0",
 22674 => x"C0C0C0A4A482F899",
 22675 => x"C0C0C0A4A482F892",
 22676 => x"C0C0C0A4A482F882",
 22677 => x"C0C0C0A4A482F8F8",
 22678 => x"C0C0C0A4A482F880",
 22679 => x"C0C0C0A4A482F890",
 22680 => x"C0C0C0A4A48280C0",
 22681 => x"C0C0C0A4A48280F9",
 22682 => x"C0C0C0A4A48280A4",
 22683 => x"C0C0C0A4A48280B0",
 22684 => x"C0C0C0A4A4828099",
 22685 => x"C0C0C0A4A4828092",
 22686 => x"C0C0C0A4A4828082",
 22687 => x"C0C0C0A4A48280F8",
 22688 => x"C0C0C0A4A4828080",
 22689 => x"C0C0C0A4A4828090",
 22690 => x"C0C0C0A4A48290C0",
 22691 => x"C0C0C0A4A48290F9",
 22692 => x"C0C0C0A4A48290A4",
 22693 => x"C0C0C0A4A48290B0",
 22694 => x"C0C0C0A4A4829099",
 22695 => x"C0C0C0A4A4829092",
 22696 => x"C0C0C0A4A4829082",
 22697 => x"C0C0C0A4A48290F8",
 22698 => x"C0C0C0A4A4829080",
 22699 => x"C0C0C0A4A4829090",
 22700 => x"C0C0C0A4A4F8C0C0",
 22701 => x"C0C0C0A4A4F8C0F9",
 22702 => x"C0C0C0A4A4F8C0A4",
 22703 => x"C0C0C0A4A4F8C0B0",
 22704 => x"C0C0C0A4A4F8C099",
 22705 => x"C0C0C0A4A4F8C092",
 22706 => x"C0C0C0A4A4F8C082",
 22707 => x"C0C0C0A4A4F8C0F8",
 22708 => x"C0C0C0A4A4F8C080",
 22709 => x"C0C0C0A4A4F8C090",
 22710 => x"C0C0C0A4A4F8F9C0",
 22711 => x"C0C0C0A4A4F8F9F9",
 22712 => x"C0C0C0A4A4F8F9A4",
 22713 => x"C0C0C0A4A4F8F9B0",
 22714 => x"C0C0C0A4A4F8F999",
 22715 => x"C0C0C0A4A4F8F992",
 22716 => x"C0C0C0A4A4F8F982",
 22717 => x"C0C0C0A4A4F8F9F8",
 22718 => x"C0C0C0A4A4F8F980",
 22719 => x"C0C0C0A4A4F8F990",
 22720 => x"C0C0C0A4A4F8A4C0",
 22721 => x"C0C0C0A4A4F8A4F9",
 22722 => x"C0C0C0A4A4F8A4A4",
 22723 => x"C0C0C0A4A4F8A4B0",
 22724 => x"C0C0C0A4A4F8A499",
 22725 => x"C0C0C0A4A4F8A492",
 22726 => x"C0C0C0A4A4F8A482",
 22727 => x"C0C0C0A4A4F8A4F8",
 22728 => x"C0C0C0A4A4F8A480",
 22729 => x"C0C0C0A4A4F8A490",
 22730 => x"C0C0C0A4A4F8B0C0",
 22731 => x"C0C0C0A4A4F8B0F9",
 22732 => x"C0C0C0A4A4F8B0A4",
 22733 => x"C0C0C0A4A4F8B0B0",
 22734 => x"C0C0C0A4A4F8B099",
 22735 => x"C0C0C0A4A4F8B092",
 22736 => x"C0C0C0A4A4F8B082",
 22737 => x"C0C0C0A4A4F8B0F8",
 22738 => x"C0C0C0A4A4F8B080",
 22739 => x"C0C0C0A4A4F8B090",
 22740 => x"C0C0C0A4A4F899C0",
 22741 => x"C0C0C0A4A4F899F9",
 22742 => x"C0C0C0A4A4F899A4",
 22743 => x"C0C0C0A4A4F899B0",
 22744 => x"C0C0C0A4A4F89999",
 22745 => x"C0C0C0A4A4F89992",
 22746 => x"C0C0C0A4A4F89982",
 22747 => x"C0C0C0A4A4F899F8",
 22748 => x"C0C0C0A4A4F89980",
 22749 => x"C0C0C0A4A4F89990",
 22750 => x"C0C0C0A4A4F892C0",
 22751 => x"C0C0C0A4A4F892F9",
 22752 => x"C0C0C0A4A4F892A4",
 22753 => x"C0C0C0A4A4F892B0",
 22754 => x"C0C0C0A4A4F89299",
 22755 => x"C0C0C0A4A4F89292",
 22756 => x"C0C0C0A4A4F89282",
 22757 => x"C0C0C0A4A4F892F8",
 22758 => x"C0C0C0A4A4F89280",
 22759 => x"C0C0C0A4A4F89290",
 22760 => x"C0C0C0A4A4F882C0",
 22761 => x"C0C0C0A4A4F882F9",
 22762 => x"C0C0C0A4A4F882A4",
 22763 => x"C0C0C0A4A4F882B0",
 22764 => x"C0C0C0A4A4F88299",
 22765 => x"C0C0C0A4A4F88292",
 22766 => x"C0C0C0A4A4F88282",
 22767 => x"C0C0C0A4A4F882F8",
 22768 => x"C0C0C0A4A4F88280",
 22769 => x"C0C0C0A4A4F88290",
 22770 => x"C0C0C0A4A4F8F8C0",
 22771 => x"C0C0C0A4A4F8F8F9",
 22772 => x"C0C0C0A4A4F8F8A4",
 22773 => x"C0C0C0A4A4F8F8B0",
 22774 => x"C0C0C0A4A4F8F899",
 22775 => x"C0C0C0A4A4F8F892",
 22776 => x"C0C0C0A4A4F8F882",
 22777 => x"C0C0C0A4A4F8F8F8",
 22778 => x"C0C0C0A4A4F8F880",
 22779 => x"C0C0C0A4A4F8F890",
 22780 => x"C0C0C0A4A4F880C0",
 22781 => x"C0C0C0A4A4F880F9",
 22782 => x"C0C0C0A4A4F880A4",
 22783 => x"C0C0C0A4A4F880B0",
 22784 => x"C0C0C0A4A4F88099",
 22785 => x"C0C0C0A4A4F88092",
 22786 => x"C0C0C0A4A4F88082",
 22787 => x"C0C0C0A4A4F880F8",
 22788 => x"C0C0C0A4A4F88080",
 22789 => x"C0C0C0A4A4F88090",
 22790 => x"C0C0C0A4A4F890C0",
 22791 => x"C0C0C0A4A4F890F9",
 22792 => x"C0C0C0A4A4F890A4",
 22793 => x"C0C0C0A4A4F890B0",
 22794 => x"C0C0C0A4A4F89099",
 22795 => x"C0C0C0A4A4F89092",
 22796 => x"C0C0C0A4A4F89082",
 22797 => x"C0C0C0A4A4F890F8",
 22798 => x"C0C0C0A4A4F89080",
 22799 => x"C0C0C0A4A4F89090",
 22800 => x"C0C0C0A4A480C0C0",
 22801 => x"C0C0C0A4A480C0F9",
 22802 => x"C0C0C0A4A480C0A4",
 22803 => x"C0C0C0A4A480C0B0",
 22804 => x"C0C0C0A4A480C099",
 22805 => x"C0C0C0A4A480C092",
 22806 => x"C0C0C0A4A480C082",
 22807 => x"C0C0C0A4A480C0F8",
 22808 => x"C0C0C0A4A480C080",
 22809 => x"C0C0C0A4A480C090",
 22810 => x"C0C0C0A4A480F9C0",
 22811 => x"C0C0C0A4A480F9F9",
 22812 => x"C0C0C0A4A480F9A4",
 22813 => x"C0C0C0A4A480F9B0",
 22814 => x"C0C0C0A4A480F999",
 22815 => x"C0C0C0A4A480F992",
 22816 => x"C0C0C0A4A480F982",
 22817 => x"C0C0C0A4A480F9F8",
 22818 => x"C0C0C0A4A480F980",
 22819 => x"C0C0C0A4A480F990",
 22820 => x"C0C0C0A4A480A4C0",
 22821 => x"C0C0C0A4A480A4F9",
 22822 => x"C0C0C0A4A480A4A4",
 22823 => x"C0C0C0A4A480A4B0",
 22824 => x"C0C0C0A4A480A499",
 22825 => x"C0C0C0A4A480A492",
 22826 => x"C0C0C0A4A480A482",
 22827 => x"C0C0C0A4A480A4F8",
 22828 => x"C0C0C0A4A480A480",
 22829 => x"C0C0C0A4A480A490",
 22830 => x"C0C0C0A4A480B0C0",
 22831 => x"C0C0C0A4A480B0F9",
 22832 => x"C0C0C0A4A480B0A4",
 22833 => x"C0C0C0A4A480B0B0",
 22834 => x"C0C0C0A4A480B099",
 22835 => x"C0C0C0A4A480B092",
 22836 => x"C0C0C0A4A480B082",
 22837 => x"C0C0C0A4A480B0F8",
 22838 => x"C0C0C0A4A480B080",
 22839 => x"C0C0C0A4A480B090",
 22840 => x"C0C0C0A4A48099C0",
 22841 => x"C0C0C0A4A48099F9",
 22842 => x"C0C0C0A4A48099A4",
 22843 => x"C0C0C0A4A48099B0",
 22844 => x"C0C0C0A4A4809999",
 22845 => x"C0C0C0A4A4809992",
 22846 => x"C0C0C0A4A4809982",
 22847 => x"C0C0C0A4A48099F8",
 22848 => x"C0C0C0A4A4809980",
 22849 => x"C0C0C0A4A4809990",
 22850 => x"C0C0C0A4A48092C0",
 22851 => x"C0C0C0A4A48092F9",
 22852 => x"C0C0C0A4A48092A4",
 22853 => x"C0C0C0A4A48092B0",
 22854 => x"C0C0C0A4A4809299",
 22855 => x"C0C0C0A4A4809292",
 22856 => x"C0C0C0A4A4809282",
 22857 => x"C0C0C0A4A48092F8",
 22858 => x"C0C0C0A4A4809280",
 22859 => x"C0C0C0A4A4809290",
 22860 => x"C0C0C0A4A48082C0",
 22861 => x"C0C0C0A4A48082F9",
 22862 => x"C0C0C0A4A48082A4",
 22863 => x"C0C0C0A4A48082B0",
 22864 => x"C0C0C0A4A4808299",
 22865 => x"C0C0C0A4A4808292",
 22866 => x"C0C0C0A4A4808282",
 22867 => x"C0C0C0A4A48082F8",
 22868 => x"C0C0C0A4A4808280",
 22869 => x"C0C0C0A4A4808290",
 22870 => x"C0C0C0A4A480F8C0",
 22871 => x"C0C0C0A4A480F8F9",
 22872 => x"C0C0C0A4A480F8A4",
 22873 => x"C0C0C0A4A480F8B0",
 22874 => x"C0C0C0A4A480F899",
 22875 => x"C0C0C0A4A480F892",
 22876 => x"C0C0C0A4A480F882",
 22877 => x"C0C0C0A4A480F8F8",
 22878 => x"C0C0C0A4A480F880",
 22879 => x"C0C0C0A4A480F890",
 22880 => x"C0C0C0A4A48080C0",
 22881 => x"C0C0C0A4A48080F9",
 22882 => x"C0C0C0A4A48080A4",
 22883 => x"C0C0C0A4A48080B0",
 22884 => x"C0C0C0A4A4808099",
 22885 => x"C0C0C0A4A4808092",
 22886 => x"C0C0C0A4A4808082",
 22887 => x"C0C0C0A4A48080F8",
 22888 => x"C0C0C0A4A4808080",
 22889 => x"C0C0C0A4A4808090",
 22890 => x"C0C0C0A4A48090C0",
 22891 => x"C0C0C0A4A48090F9",
 22892 => x"C0C0C0A4A48090A4",
 22893 => x"C0C0C0A4A48090B0",
 22894 => x"C0C0C0A4A4809099",
 22895 => x"C0C0C0A4A4809092",
 22896 => x"C0C0C0A4A4809082",
 22897 => x"C0C0C0A4A48090F8",
 22898 => x"C0C0C0A4A4809080",
 22899 => x"C0C0C0A4A4809090",
 22900 => x"C0C0C0A4A490C0C0",
 22901 => x"C0C0C0A4A490C0F9",
 22902 => x"C0C0C0A4A490C0A4",
 22903 => x"C0C0C0A4A490C0B0",
 22904 => x"C0C0C0A4A490C099",
 22905 => x"C0C0C0A4A490C092",
 22906 => x"C0C0C0A4A490C082",
 22907 => x"C0C0C0A4A490C0F8",
 22908 => x"C0C0C0A4A490C080",
 22909 => x"C0C0C0A4A490C090",
 22910 => x"C0C0C0A4A490F9C0",
 22911 => x"C0C0C0A4A490F9F9",
 22912 => x"C0C0C0A4A490F9A4",
 22913 => x"C0C0C0A4A490F9B0",
 22914 => x"C0C0C0A4A490F999",
 22915 => x"C0C0C0A4A490F992",
 22916 => x"C0C0C0A4A490F982",
 22917 => x"C0C0C0A4A490F9F8",
 22918 => x"C0C0C0A4A490F980",
 22919 => x"C0C0C0A4A490F990",
 22920 => x"C0C0C0A4A490A4C0",
 22921 => x"C0C0C0A4A490A4F9",
 22922 => x"C0C0C0A4A490A4A4",
 22923 => x"C0C0C0A4A490A4B0",
 22924 => x"C0C0C0A4A490A499",
 22925 => x"C0C0C0A4A490A492",
 22926 => x"C0C0C0A4A490A482",
 22927 => x"C0C0C0A4A490A4F8",
 22928 => x"C0C0C0A4A490A480",
 22929 => x"C0C0C0A4A490A490",
 22930 => x"C0C0C0A4A490B0C0",
 22931 => x"C0C0C0A4A490B0F9",
 22932 => x"C0C0C0A4A490B0A4",
 22933 => x"C0C0C0A4A490B0B0",
 22934 => x"C0C0C0A4A490B099",
 22935 => x"C0C0C0A4A490B092",
 22936 => x"C0C0C0A4A490B082",
 22937 => x"C0C0C0A4A490B0F8",
 22938 => x"C0C0C0A4A490B080",
 22939 => x"C0C0C0A4A490B090",
 22940 => x"C0C0C0A4A49099C0",
 22941 => x"C0C0C0A4A49099F9",
 22942 => x"C0C0C0A4A49099A4",
 22943 => x"C0C0C0A4A49099B0",
 22944 => x"C0C0C0A4A4909999",
 22945 => x"C0C0C0A4A4909992",
 22946 => x"C0C0C0A4A4909982",
 22947 => x"C0C0C0A4A49099F8",
 22948 => x"C0C0C0A4A4909980",
 22949 => x"C0C0C0A4A4909990",
 22950 => x"C0C0C0A4A49092C0",
 22951 => x"C0C0C0A4A49092F9",
 22952 => x"C0C0C0A4A49092A4",
 22953 => x"C0C0C0A4A49092B0",
 22954 => x"C0C0C0A4A4909299",
 22955 => x"C0C0C0A4A4909292",
 22956 => x"C0C0C0A4A4909282",
 22957 => x"C0C0C0A4A49092F8",
 22958 => x"C0C0C0A4A4909280",
 22959 => x"C0C0C0A4A4909290",
 22960 => x"C0C0C0A4A49082C0",
 22961 => x"C0C0C0A4A49082F9",
 22962 => x"C0C0C0A4A49082A4",
 22963 => x"C0C0C0A4A49082B0",
 22964 => x"C0C0C0A4A4908299",
 22965 => x"C0C0C0A4A4908292",
 22966 => x"C0C0C0A4A4908282",
 22967 => x"C0C0C0A4A49082F8",
 22968 => x"C0C0C0A4A4908280",
 22969 => x"C0C0C0A4A4908290",
 22970 => x"C0C0C0A4A490F8C0",
 22971 => x"C0C0C0A4A490F8F9",
 22972 => x"C0C0C0A4A490F8A4",
 22973 => x"C0C0C0A4A490F8B0",
 22974 => x"C0C0C0A4A490F899",
 22975 => x"C0C0C0A4A490F892",
 22976 => x"C0C0C0A4A490F882",
 22977 => x"C0C0C0A4A490F8F8",
 22978 => x"C0C0C0A4A490F880",
 22979 => x"C0C0C0A4A490F890",
 22980 => x"C0C0C0A4A49080C0",
 22981 => x"C0C0C0A4A49080F9",
 22982 => x"C0C0C0A4A49080A4",
 22983 => x"C0C0C0A4A49080B0",
 22984 => x"C0C0C0A4A4908099",
 22985 => x"C0C0C0A4A4908092",
 22986 => x"C0C0C0A4A4908082",
 22987 => x"C0C0C0A4A49080F8",
 22988 => x"C0C0C0A4A4908080",
 22989 => x"C0C0C0A4A4908090",
 22990 => x"C0C0C0A4A49090C0",
 22991 => x"C0C0C0A4A49090F9",
 22992 => x"C0C0C0A4A49090A4",
 22993 => x"C0C0C0A4A49090B0",
 22994 => x"C0C0C0A4A4909099",
 22995 => x"C0C0C0A4A4909092",
 22996 => x"C0C0C0A4A4909082",
 22997 => x"C0C0C0A4A49090F8",
 22998 => x"C0C0C0A4A4909080",
 22999 => x"C0C0C0A4A4909090",
 23000 => x"C0C0C0A4B0C0C0C0",
 23001 => x"C0C0C0A4B0C0C0F9",
 23002 => x"C0C0C0A4B0C0C0A4",
 23003 => x"C0C0C0A4B0C0C0B0",
 23004 => x"C0C0C0A4B0C0C099",
 23005 => x"C0C0C0A4B0C0C092",
 23006 => x"C0C0C0A4B0C0C082",
 23007 => x"C0C0C0A4B0C0C0F8",
 23008 => x"C0C0C0A4B0C0C080",
 23009 => x"C0C0C0A4B0C0C090",
 23010 => x"C0C0C0A4B0C0F9C0",
 23011 => x"C0C0C0A4B0C0F9F9",
 23012 => x"C0C0C0A4B0C0F9A4",
 23013 => x"C0C0C0A4B0C0F9B0",
 23014 => x"C0C0C0A4B0C0F999",
 23015 => x"C0C0C0A4B0C0F992",
 23016 => x"C0C0C0A4B0C0F982",
 23017 => x"C0C0C0A4B0C0F9F8",
 23018 => x"C0C0C0A4B0C0F980",
 23019 => x"C0C0C0A4B0C0F990",
 23020 => x"C0C0C0A4B0C0A4C0",
 23021 => x"C0C0C0A4B0C0A4F9",
 23022 => x"C0C0C0A4B0C0A4A4",
 23023 => x"C0C0C0A4B0C0A4B0",
 23024 => x"C0C0C0A4B0C0A499",
 23025 => x"C0C0C0A4B0C0A492",
 23026 => x"C0C0C0A4B0C0A482",
 23027 => x"C0C0C0A4B0C0A4F8",
 23028 => x"C0C0C0A4B0C0A480",
 23029 => x"C0C0C0A4B0C0A490",
 23030 => x"C0C0C0A4B0C0B0C0",
 23031 => x"C0C0C0A4B0C0B0F9",
 23032 => x"C0C0C0A4B0C0B0A4",
 23033 => x"C0C0C0A4B0C0B0B0",
 23034 => x"C0C0C0A4B0C0B099",
 23035 => x"C0C0C0A4B0C0B092",
 23036 => x"C0C0C0A4B0C0B082",
 23037 => x"C0C0C0A4B0C0B0F8",
 23038 => x"C0C0C0A4B0C0B080",
 23039 => x"C0C0C0A4B0C0B090",
 23040 => x"C0C0C0A4B0C099C0",
 23041 => x"C0C0C0A4B0C099F9",
 23042 => x"C0C0C0A4B0C099A4",
 23043 => x"C0C0C0A4B0C099B0",
 23044 => x"C0C0C0A4B0C09999",
 23045 => x"C0C0C0A4B0C09992",
 23046 => x"C0C0C0A4B0C09982",
 23047 => x"C0C0C0A4B0C099F8",
 23048 => x"C0C0C0A4B0C09980",
 23049 => x"C0C0C0A4B0C09990",
 23050 => x"C0C0C0A4B0C092C0",
 23051 => x"C0C0C0A4B0C092F9",
 23052 => x"C0C0C0A4B0C092A4",
 23053 => x"C0C0C0A4B0C092B0",
 23054 => x"C0C0C0A4B0C09299",
 23055 => x"C0C0C0A4B0C09292",
 23056 => x"C0C0C0A4B0C09282",
 23057 => x"C0C0C0A4B0C092F8",
 23058 => x"C0C0C0A4B0C09280",
 23059 => x"C0C0C0A4B0C09290",
 23060 => x"C0C0C0A4B0C082C0",
 23061 => x"C0C0C0A4B0C082F9",
 23062 => x"C0C0C0A4B0C082A4",
 23063 => x"C0C0C0A4B0C082B0",
 23064 => x"C0C0C0A4B0C08299",
 23065 => x"C0C0C0A4B0C08292",
 23066 => x"C0C0C0A4B0C08282",
 23067 => x"C0C0C0A4B0C082F8",
 23068 => x"C0C0C0A4B0C08280",
 23069 => x"C0C0C0A4B0C08290",
 23070 => x"C0C0C0A4B0C0F8C0",
 23071 => x"C0C0C0A4B0C0F8F9",
 23072 => x"C0C0C0A4B0C0F8A4",
 23073 => x"C0C0C0A4B0C0F8B0",
 23074 => x"C0C0C0A4B0C0F899",
 23075 => x"C0C0C0A4B0C0F892",
 23076 => x"C0C0C0A4B0C0F882",
 23077 => x"C0C0C0A4B0C0F8F8",
 23078 => x"C0C0C0A4B0C0F880",
 23079 => x"C0C0C0A4B0C0F890",
 23080 => x"C0C0C0A4B0C080C0",
 23081 => x"C0C0C0A4B0C080F9",
 23082 => x"C0C0C0A4B0C080A4",
 23083 => x"C0C0C0A4B0C080B0",
 23084 => x"C0C0C0A4B0C08099",
 23085 => x"C0C0C0A4B0C08092",
 23086 => x"C0C0C0A4B0C08082",
 23087 => x"C0C0C0A4B0C080F8",
 23088 => x"C0C0C0A4B0C08080",
 23089 => x"C0C0C0A4B0C08090",
 23090 => x"C0C0C0A4B0C090C0",
 23091 => x"C0C0C0A4B0C090F9",
 23092 => x"C0C0C0A4B0C090A4",
 23093 => x"C0C0C0A4B0C090B0",
 23094 => x"C0C0C0A4B0C09099",
 23095 => x"C0C0C0A4B0C09092",
 23096 => x"C0C0C0A4B0C09082",
 23097 => x"C0C0C0A4B0C090F8",
 23098 => x"C0C0C0A4B0C09080",
 23099 => x"C0C0C0A4B0C09090",
 23100 => x"C0C0C0A4B0F9C0C0",
 23101 => x"C0C0C0A4B0F9C0F9",
 23102 => x"C0C0C0A4B0F9C0A4",
 23103 => x"C0C0C0A4B0F9C0B0",
 23104 => x"C0C0C0A4B0F9C099",
 23105 => x"C0C0C0A4B0F9C092",
 23106 => x"C0C0C0A4B0F9C082",
 23107 => x"C0C0C0A4B0F9C0F8",
 23108 => x"C0C0C0A4B0F9C080",
 23109 => x"C0C0C0A4B0F9C090",
 23110 => x"C0C0C0A4B0F9F9C0",
 23111 => x"C0C0C0A4B0F9F9F9",
 23112 => x"C0C0C0A4B0F9F9A4",
 23113 => x"C0C0C0A4B0F9F9B0",
 23114 => x"C0C0C0A4B0F9F999",
 23115 => x"C0C0C0A4B0F9F992",
 23116 => x"C0C0C0A4B0F9F982",
 23117 => x"C0C0C0A4B0F9F9F8",
 23118 => x"C0C0C0A4B0F9F980",
 23119 => x"C0C0C0A4B0F9F990",
 23120 => x"C0C0C0A4B0F9A4C0",
 23121 => x"C0C0C0A4B0F9A4F9",
 23122 => x"C0C0C0A4B0F9A4A4",
 23123 => x"C0C0C0A4B0F9A4B0",
 23124 => x"C0C0C0A4B0F9A499",
 23125 => x"C0C0C0A4B0F9A492",
 23126 => x"C0C0C0A4B0F9A482",
 23127 => x"C0C0C0A4B0F9A4F8",
 23128 => x"C0C0C0A4B0F9A480",
 23129 => x"C0C0C0A4B0F9A490",
 23130 => x"C0C0C0A4B0F9B0C0",
 23131 => x"C0C0C0A4B0F9B0F9",
 23132 => x"C0C0C0A4B0F9B0A4",
 23133 => x"C0C0C0A4B0F9B0B0",
 23134 => x"C0C0C0A4B0F9B099",
 23135 => x"C0C0C0A4B0F9B092",
 23136 => x"C0C0C0A4B0F9B082",
 23137 => x"C0C0C0A4B0F9B0F8",
 23138 => x"C0C0C0A4B0F9B080",
 23139 => x"C0C0C0A4B0F9B090",
 23140 => x"C0C0C0A4B0F999C0",
 23141 => x"C0C0C0A4B0F999F9",
 23142 => x"C0C0C0A4B0F999A4",
 23143 => x"C0C0C0A4B0F999B0",
 23144 => x"C0C0C0A4B0F99999",
 23145 => x"C0C0C0A4B0F99992",
 23146 => x"C0C0C0A4B0F99982",
 23147 => x"C0C0C0A4B0F999F8",
 23148 => x"C0C0C0A4B0F99980",
 23149 => x"C0C0C0A4B0F99990",
 23150 => x"C0C0C0A4B0F992C0",
 23151 => x"C0C0C0A4B0F992F9",
 23152 => x"C0C0C0A4B0F992A4",
 23153 => x"C0C0C0A4B0F992B0",
 23154 => x"C0C0C0A4B0F99299",
 23155 => x"C0C0C0A4B0F99292",
 23156 => x"C0C0C0A4B0F99282",
 23157 => x"C0C0C0A4B0F992F8",
 23158 => x"C0C0C0A4B0F99280",
 23159 => x"C0C0C0A4B0F99290",
 23160 => x"C0C0C0A4B0F982C0",
 23161 => x"C0C0C0A4B0F982F9",
 23162 => x"C0C0C0A4B0F982A4",
 23163 => x"C0C0C0A4B0F982B0",
 23164 => x"C0C0C0A4B0F98299",
 23165 => x"C0C0C0A4B0F98292",
 23166 => x"C0C0C0A4B0F98282",
 23167 => x"C0C0C0A4B0F982F8",
 23168 => x"C0C0C0A4B0F98280",
 23169 => x"C0C0C0A4B0F98290",
 23170 => x"C0C0C0A4B0F9F8C0",
 23171 => x"C0C0C0A4B0F9F8F9",
 23172 => x"C0C0C0A4B0F9F8A4",
 23173 => x"C0C0C0A4B0F9F8B0",
 23174 => x"C0C0C0A4B0F9F899",
 23175 => x"C0C0C0A4B0F9F892",
 23176 => x"C0C0C0A4B0F9F882",
 23177 => x"C0C0C0A4B0F9F8F8",
 23178 => x"C0C0C0A4B0F9F880",
 23179 => x"C0C0C0A4B0F9F890",
 23180 => x"C0C0C0A4B0F980C0",
 23181 => x"C0C0C0A4B0F980F9",
 23182 => x"C0C0C0A4B0F980A4",
 23183 => x"C0C0C0A4B0F980B0",
 23184 => x"C0C0C0A4B0F98099",
 23185 => x"C0C0C0A4B0F98092",
 23186 => x"C0C0C0A4B0F98082",
 23187 => x"C0C0C0A4B0F980F8",
 23188 => x"C0C0C0A4B0F98080",
 23189 => x"C0C0C0A4B0F98090",
 23190 => x"C0C0C0A4B0F990C0",
 23191 => x"C0C0C0A4B0F990F9",
 23192 => x"C0C0C0A4B0F990A4",
 23193 => x"C0C0C0A4B0F990B0",
 23194 => x"C0C0C0A4B0F99099",
 23195 => x"C0C0C0A4B0F99092",
 23196 => x"C0C0C0A4B0F99082",
 23197 => x"C0C0C0A4B0F990F8",
 23198 => x"C0C0C0A4B0F99080",
 23199 => x"C0C0C0A4B0F99090",
 23200 => x"C0C0C0A4B0A4C0C0",
 23201 => x"C0C0C0A4B0A4C0F9",
 23202 => x"C0C0C0A4B0A4C0A4",
 23203 => x"C0C0C0A4B0A4C0B0",
 23204 => x"C0C0C0A4B0A4C099",
 23205 => x"C0C0C0A4B0A4C092",
 23206 => x"C0C0C0A4B0A4C082",
 23207 => x"C0C0C0A4B0A4C0F8",
 23208 => x"C0C0C0A4B0A4C080",
 23209 => x"C0C0C0A4B0A4C090",
 23210 => x"C0C0C0A4B0A4F9C0",
 23211 => x"C0C0C0A4B0A4F9F9",
 23212 => x"C0C0C0A4B0A4F9A4",
 23213 => x"C0C0C0A4B0A4F9B0",
 23214 => x"C0C0C0A4B0A4F999",
 23215 => x"C0C0C0A4B0A4F992",
 23216 => x"C0C0C0A4B0A4F982",
 23217 => x"C0C0C0A4B0A4F9F8",
 23218 => x"C0C0C0A4B0A4F980",
 23219 => x"C0C0C0A4B0A4F990",
 23220 => x"C0C0C0A4B0A4A4C0",
 23221 => x"C0C0C0A4B0A4A4F9",
 23222 => x"C0C0C0A4B0A4A4A4",
 23223 => x"C0C0C0A4B0A4A4B0",
 23224 => x"C0C0C0A4B0A4A499",
 23225 => x"C0C0C0A4B0A4A492",
 23226 => x"C0C0C0A4B0A4A482",
 23227 => x"C0C0C0A4B0A4A4F8",
 23228 => x"C0C0C0A4B0A4A480",
 23229 => x"C0C0C0A4B0A4A490",
 23230 => x"C0C0C0A4B0A4B0C0",
 23231 => x"C0C0C0A4B0A4B0F9",
 23232 => x"C0C0C0A4B0A4B0A4",
 23233 => x"C0C0C0A4B0A4B0B0",
 23234 => x"C0C0C0A4B0A4B099",
 23235 => x"C0C0C0A4B0A4B092",
 23236 => x"C0C0C0A4B0A4B082",
 23237 => x"C0C0C0A4B0A4B0F8",
 23238 => x"C0C0C0A4B0A4B080",
 23239 => x"C0C0C0A4B0A4B090",
 23240 => x"C0C0C0A4B0A499C0",
 23241 => x"C0C0C0A4B0A499F9",
 23242 => x"C0C0C0A4B0A499A4",
 23243 => x"C0C0C0A4B0A499B0",
 23244 => x"C0C0C0A4B0A49999",
 23245 => x"C0C0C0A4B0A49992",
 23246 => x"C0C0C0A4B0A49982",
 23247 => x"C0C0C0A4B0A499F8",
 23248 => x"C0C0C0A4B0A49980",
 23249 => x"C0C0C0A4B0A49990",
 23250 => x"C0C0C0A4B0A492C0",
 23251 => x"C0C0C0A4B0A492F9",
 23252 => x"C0C0C0A4B0A492A4",
 23253 => x"C0C0C0A4B0A492B0",
 23254 => x"C0C0C0A4B0A49299",
 23255 => x"C0C0C0A4B0A49292",
 23256 => x"C0C0C0A4B0A49282",
 23257 => x"C0C0C0A4B0A492F8",
 23258 => x"C0C0C0A4B0A49280",
 23259 => x"C0C0C0A4B0A49290",
 23260 => x"C0C0C0A4B0A482C0",
 23261 => x"C0C0C0A4B0A482F9",
 23262 => x"C0C0C0A4B0A482A4",
 23263 => x"C0C0C0A4B0A482B0",
 23264 => x"C0C0C0A4B0A48299",
 23265 => x"C0C0C0A4B0A48292",
 23266 => x"C0C0C0A4B0A48282",
 23267 => x"C0C0C0A4B0A482F8",
 23268 => x"C0C0C0A4B0A48280",
 23269 => x"C0C0C0A4B0A48290",
 23270 => x"C0C0C0A4B0A4F8C0",
 23271 => x"C0C0C0A4B0A4F8F9",
 23272 => x"C0C0C0A4B0A4F8A4",
 23273 => x"C0C0C0A4B0A4F8B0",
 23274 => x"C0C0C0A4B0A4F899",
 23275 => x"C0C0C0A4B0A4F892",
 23276 => x"C0C0C0A4B0A4F882",
 23277 => x"C0C0C0A4B0A4F8F8",
 23278 => x"C0C0C0A4B0A4F880",
 23279 => x"C0C0C0A4B0A4F890",
 23280 => x"C0C0C0A4B0A480C0",
 23281 => x"C0C0C0A4B0A480F9",
 23282 => x"C0C0C0A4B0A480A4",
 23283 => x"C0C0C0A4B0A480B0",
 23284 => x"C0C0C0A4B0A48099",
 23285 => x"C0C0C0A4B0A48092",
 23286 => x"C0C0C0A4B0A48082",
 23287 => x"C0C0C0A4B0A480F8",
 23288 => x"C0C0C0A4B0A48080",
 23289 => x"C0C0C0A4B0A48090",
 23290 => x"C0C0C0A4B0A490C0",
 23291 => x"C0C0C0A4B0A490F9",
 23292 => x"C0C0C0A4B0A490A4",
 23293 => x"C0C0C0A4B0A490B0",
 23294 => x"C0C0C0A4B0A49099",
 23295 => x"C0C0C0A4B0A49092",
 23296 => x"C0C0C0A4B0A49082",
 23297 => x"C0C0C0A4B0A490F8",
 23298 => x"C0C0C0A4B0A49080",
 23299 => x"C0C0C0A4B0A49090",
 23300 => x"C0C0C0A4B0B0C0C0",
 23301 => x"C0C0C0A4B0B0C0F9",
 23302 => x"C0C0C0A4B0B0C0A4",
 23303 => x"C0C0C0A4B0B0C0B0",
 23304 => x"C0C0C0A4B0B0C099",
 23305 => x"C0C0C0A4B0B0C092",
 23306 => x"C0C0C0A4B0B0C082",
 23307 => x"C0C0C0A4B0B0C0F8",
 23308 => x"C0C0C0A4B0B0C080",
 23309 => x"C0C0C0A4B0B0C090",
 23310 => x"C0C0C0A4B0B0F9C0",
 23311 => x"C0C0C0A4B0B0F9F9",
 23312 => x"C0C0C0A4B0B0F9A4",
 23313 => x"C0C0C0A4B0B0F9B0",
 23314 => x"C0C0C0A4B0B0F999",
 23315 => x"C0C0C0A4B0B0F992",
 23316 => x"C0C0C0A4B0B0F982",
 23317 => x"C0C0C0A4B0B0F9F8",
 23318 => x"C0C0C0A4B0B0F980",
 23319 => x"C0C0C0A4B0B0F990",
 23320 => x"C0C0C0A4B0B0A4C0",
 23321 => x"C0C0C0A4B0B0A4F9",
 23322 => x"C0C0C0A4B0B0A4A4",
 23323 => x"C0C0C0A4B0B0A4B0",
 23324 => x"C0C0C0A4B0B0A499",
 23325 => x"C0C0C0A4B0B0A492",
 23326 => x"C0C0C0A4B0B0A482",
 23327 => x"C0C0C0A4B0B0A4F8",
 23328 => x"C0C0C0A4B0B0A480",
 23329 => x"C0C0C0A4B0B0A490",
 23330 => x"C0C0C0A4B0B0B0C0",
 23331 => x"C0C0C0A4B0B0B0F9",
 23332 => x"C0C0C0A4B0B0B0A4",
 23333 => x"C0C0C0A4B0B0B0B0",
 23334 => x"C0C0C0A4B0B0B099",
 23335 => x"C0C0C0A4B0B0B092",
 23336 => x"C0C0C0A4B0B0B082",
 23337 => x"C0C0C0A4B0B0B0F8",
 23338 => x"C0C0C0A4B0B0B080",
 23339 => x"C0C0C0A4B0B0B090",
 23340 => x"C0C0C0A4B0B099C0",
 23341 => x"C0C0C0A4B0B099F9",
 23342 => x"C0C0C0A4B0B099A4",
 23343 => x"C0C0C0A4B0B099B0",
 23344 => x"C0C0C0A4B0B09999",
 23345 => x"C0C0C0A4B0B09992",
 23346 => x"C0C0C0A4B0B09982",
 23347 => x"C0C0C0A4B0B099F8",
 23348 => x"C0C0C0A4B0B09980",
 23349 => x"C0C0C0A4B0B09990",
 23350 => x"C0C0C0A4B0B092C0",
 23351 => x"C0C0C0A4B0B092F9",
 23352 => x"C0C0C0A4B0B092A4",
 23353 => x"C0C0C0A4B0B092B0",
 23354 => x"C0C0C0A4B0B09299",
 23355 => x"C0C0C0A4B0B09292",
 23356 => x"C0C0C0A4B0B09282",
 23357 => x"C0C0C0A4B0B092F8",
 23358 => x"C0C0C0A4B0B09280",
 23359 => x"C0C0C0A4B0B09290",
 23360 => x"C0C0C0A4B0B082C0",
 23361 => x"C0C0C0A4B0B082F9",
 23362 => x"C0C0C0A4B0B082A4",
 23363 => x"C0C0C0A4B0B082B0",
 23364 => x"C0C0C0A4B0B08299",
 23365 => x"C0C0C0A4B0B08292",
 23366 => x"C0C0C0A4B0B08282",
 23367 => x"C0C0C0A4B0B082F8",
 23368 => x"C0C0C0A4B0B08280",
 23369 => x"C0C0C0A4B0B08290",
 23370 => x"C0C0C0A4B0B0F8C0",
 23371 => x"C0C0C0A4B0B0F8F9",
 23372 => x"C0C0C0A4B0B0F8A4",
 23373 => x"C0C0C0A4B0B0F8B0",
 23374 => x"C0C0C0A4B0B0F899",
 23375 => x"C0C0C0A4B0B0F892",
 23376 => x"C0C0C0A4B0B0F882",
 23377 => x"C0C0C0A4B0B0F8F8",
 23378 => x"C0C0C0A4B0B0F880",
 23379 => x"C0C0C0A4B0B0F890",
 23380 => x"C0C0C0A4B0B080C0",
 23381 => x"C0C0C0A4B0B080F9",
 23382 => x"C0C0C0A4B0B080A4",
 23383 => x"C0C0C0A4B0B080B0",
 23384 => x"C0C0C0A4B0B08099",
 23385 => x"C0C0C0A4B0B08092",
 23386 => x"C0C0C0A4B0B08082",
 23387 => x"C0C0C0A4B0B080F8",
 23388 => x"C0C0C0A4B0B08080",
 23389 => x"C0C0C0A4B0B08090",
 23390 => x"C0C0C0A4B0B090C0",
 23391 => x"C0C0C0A4B0B090F9",
 23392 => x"C0C0C0A4B0B090A4",
 23393 => x"C0C0C0A4B0B090B0",
 23394 => x"C0C0C0A4B0B09099",
 23395 => x"C0C0C0A4B0B09092",
 23396 => x"C0C0C0A4B0B09082",
 23397 => x"C0C0C0A4B0B090F8",
 23398 => x"C0C0C0A4B0B09080",
 23399 => x"C0C0C0A4B0B09090",
 23400 => x"C0C0C0A4B099C0C0",
 23401 => x"C0C0C0A4B099C0F9",
 23402 => x"C0C0C0A4B099C0A4",
 23403 => x"C0C0C0A4B099C0B0",
 23404 => x"C0C0C0A4B099C099",
 23405 => x"C0C0C0A4B099C092",
 23406 => x"C0C0C0A4B099C082",
 23407 => x"C0C0C0A4B099C0F8",
 23408 => x"C0C0C0A4B099C080",
 23409 => x"C0C0C0A4B099C090",
 23410 => x"C0C0C0A4B099F9C0",
 23411 => x"C0C0C0A4B099F9F9",
 23412 => x"C0C0C0A4B099F9A4",
 23413 => x"C0C0C0A4B099F9B0",
 23414 => x"C0C0C0A4B099F999",
 23415 => x"C0C0C0A4B099F992",
 23416 => x"C0C0C0A4B099F982",
 23417 => x"C0C0C0A4B099F9F8",
 23418 => x"C0C0C0A4B099F980",
 23419 => x"C0C0C0A4B099F990",
 23420 => x"C0C0C0A4B099A4C0",
 23421 => x"C0C0C0A4B099A4F9",
 23422 => x"C0C0C0A4B099A4A4",
 23423 => x"C0C0C0A4B099A4B0",
 23424 => x"C0C0C0A4B099A499",
 23425 => x"C0C0C0A4B099A492",
 23426 => x"C0C0C0A4B099A482",
 23427 => x"C0C0C0A4B099A4F8",
 23428 => x"C0C0C0A4B099A480",
 23429 => x"C0C0C0A4B099A490",
 23430 => x"C0C0C0A4B099B0C0",
 23431 => x"C0C0C0A4B099B0F9",
 23432 => x"C0C0C0A4B099B0A4",
 23433 => x"C0C0C0A4B099B0B0",
 23434 => x"C0C0C0A4B099B099",
 23435 => x"C0C0C0A4B099B092",
 23436 => x"C0C0C0A4B099B082",
 23437 => x"C0C0C0A4B099B0F8",
 23438 => x"C0C0C0A4B099B080",
 23439 => x"C0C0C0A4B099B090",
 23440 => x"C0C0C0A4B09999C0",
 23441 => x"C0C0C0A4B09999F9",
 23442 => x"C0C0C0A4B09999A4",
 23443 => x"C0C0C0A4B09999B0",
 23444 => x"C0C0C0A4B0999999",
 23445 => x"C0C0C0A4B0999992",
 23446 => x"C0C0C0A4B0999982",
 23447 => x"C0C0C0A4B09999F8",
 23448 => x"C0C0C0A4B0999980",
 23449 => x"C0C0C0A4B0999990",
 23450 => x"C0C0C0A4B09992C0",
 23451 => x"C0C0C0A4B09992F9",
 23452 => x"C0C0C0A4B09992A4",
 23453 => x"C0C0C0A4B09992B0",
 23454 => x"C0C0C0A4B0999299",
 23455 => x"C0C0C0A4B0999292",
 23456 => x"C0C0C0A4B0999282",
 23457 => x"C0C0C0A4B09992F8",
 23458 => x"C0C0C0A4B0999280",
 23459 => x"C0C0C0A4B0999290",
 23460 => x"C0C0C0A4B09982C0",
 23461 => x"C0C0C0A4B09982F9",
 23462 => x"C0C0C0A4B09982A4",
 23463 => x"C0C0C0A4B09982B0",
 23464 => x"C0C0C0A4B0998299",
 23465 => x"C0C0C0A4B0998292",
 23466 => x"C0C0C0A4B0998282",
 23467 => x"C0C0C0A4B09982F8",
 23468 => x"C0C0C0A4B0998280",
 23469 => x"C0C0C0A4B0998290",
 23470 => x"C0C0C0A4B099F8C0",
 23471 => x"C0C0C0A4B099F8F9",
 23472 => x"C0C0C0A4B099F8A4",
 23473 => x"C0C0C0A4B099F8B0",
 23474 => x"C0C0C0A4B099F899",
 23475 => x"C0C0C0A4B099F892",
 23476 => x"C0C0C0A4B099F882",
 23477 => x"C0C0C0A4B099F8F8",
 23478 => x"C0C0C0A4B099F880",
 23479 => x"C0C0C0A4B099F890",
 23480 => x"C0C0C0A4B09980C0",
 23481 => x"C0C0C0A4B09980F9",
 23482 => x"C0C0C0A4B09980A4",
 23483 => x"C0C0C0A4B09980B0",
 23484 => x"C0C0C0A4B0998099",
 23485 => x"C0C0C0A4B0998092",
 23486 => x"C0C0C0A4B0998082",
 23487 => x"C0C0C0A4B09980F8",
 23488 => x"C0C0C0A4B0998080",
 23489 => x"C0C0C0A4B0998090",
 23490 => x"C0C0C0A4B09990C0",
 23491 => x"C0C0C0A4B09990F9",
 23492 => x"C0C0C0A4B09990A4",
 23493 => x"C0C0C0A4B09990B0",
 23494 => x"C0C0C0A4B0999099",
 23495 => x"C0C0C0A4B0999092",
 23496 => x"C0C0C0A4B0999082",
 23497 => x"C0C0C0A4B09990F8",
 23498 => x"C0C0C0A4B0999080",
 23499 => x"C0C0C0A4B0999090",
 23500 => x"C0C0C0A4B092C0C0",
 23501 => x"C0C0C0A4B092C0F9",
 23502 => x"C0C0C0A4B092C0A4",
 23503 => x"C0C0C0A4B092C0B0",
 23504 => x"C0C0C0A4B092C099",
 23505 => x"C0C0C0A4B092C092",
 23506 => x"C0C0C0A4B092C082",
 23507 => x"C0C0C0A4B092C0F8",
 23508 => x"C0C0C0A4B092C080",
 23509 => x"C0C0C0A4B092C090",
 23510 => x"C0C0C0A4B092F9C0",
 23511 => x"C0C0C0A4B092F9F9",
 23512 => x"C0C0C0A4B092F9A4",
 23513 => x"C0C0C0A4B092F9B0",
 23514 => x"C0C0C0A4B092F999",
 23515 => x"C0C0C0A4B092F992",
 23516 => x"C0C0C0A4B092F982",
 23517 => x"C0C0C0A4B092F9F8",
 23518 => x"C0C0C0A4B092F980",
 23519 => x"C0C0C0A4B092F990",
 23520 => x"C0C0C0A4B092A4C0",
 23521 => x"C0C0C0A4B092A4F9",
 23522 => x"C0C0C0A4B092A4A4",
 23523 => x"C0C0C0A4B092A4B0",
 23524 => x"C0C0C0A4B092A499",
 23525 => x"C0C0C0A4B092A492",
 23526 => x"C0C0C0A4B092A482",
 23527 => x"C0C0C0A4B092A4F8",
 23528 => x"C0C0C0A4B092A480",
 23529 => x"C0C0C0A4B092A490",
 23530 => x"C0C0C0A4B092B0C0",
 23531 => x"C0C0C0A4B092B0F9",
 23532 => x"C0C0C0A4B092B0A4",
 23533 => x"C0C0C0A4B092B0B0",
 23534 => x"C0C0C0A4B092B099",
 23535 => x"C0C0C0A4B092B092",
 23536 => x"C0C0C0A4B092B082",
 23537 => x"C0C0C0A4B092B0F8",
 23538 => x"C0C0C0A4B092B080",
 23539 => x"C0C0C0A4B092B090",
 23540 => x"C0C0C0A4B09299C0",
 23541 => x"C0C0C0A4B09299F9",
 23542 => x"C0C0C0A4B09299A4",
 23543 => x"C0C0C0A4B09299B0",
 23544 => x"C0C0C0A4B0929999",
 23545 => x"C0C0C0A4B0929992",
 23546 => x"C0C0C0A4B0929982",
 23547 => x"C0C0C0A4B09299F8",
 23548 => x"C0C0C0A4B0929980",
 23549 => x"C0C0C0A4B0929990",
 23550 => x"C0C0C0A4B09292C0",
 23551 => x"C0C0C0A4B09292F9",
 23552 => x"C0C0C0A4B09292A4",
 23553 => x"C0C0C0A4B09292B0",
 23554 => x"C0C0C0A4B0929299",
 23555 => x"C0C0C0A4B0929292",
 23556 => x"C0C0C0A4B0929282",
 23557 => x"C0C0C0A4B09292F8",
 23558 => x"C0C0C0A4B0929280",
 23559 => x"C0C0C0A4B0929290",
 23560 => x"C0C0C0A4B09282C0",
 23561 => x"C0C0C0A4B09282F9",
 23562 => x"C0C0C0A4B09282A4",
 23563 => x"C0C0C0A4B09282B0",
 23564 => x"C0C0C0A4B0928299",
 23565 => x"C0C0C0A4B0928292",
 23566 => x"C0C0C0A4B0928282",
 23567 => x"C0C0C0A4B09282F8",
 23568 => x"C0C0C0A4B0928280",
 23569 => x"C0C0C0A4B0928290",
 23570 => x"C0C0C0A4B092F8C0",
 23571 => x"C0C0C0A4B092F8F9",
 23572 => x"C0C0C0A4B092F8A4",
 23573 => x"C0C0C0A4B092F8B0",
 23574 => x"C0C0C0A4B092F899",
 23575 => x"C0C0C0A4B092F892",
 23576 => x"C0C0C0A4B092F882",
 23577 => x"C0C0C0A4B092F8F8",
 23578 => x"C0C0C0A4B092F880",
 23579 => x"C0C0C0A4B092F890",
 23580 => x"C0C0C0A4B09280C0",
 23581 => x"C0C0C0A4B09280F9",
 23582 => x"C0C0C0A4B09280A4",
 23583 => x"C0C0C0A4B09280B0",
 23584 => x"C0C0C0A4B0928099",
 23585 => x"C0C0C0A4B0928092",
 23586 => x"C0C0C0A4B0928082",
 23587 => x"C0C0C0A4B09280F8",
 23588 => x"C0C0C0A4B0928080",
 23589 => x"C0C0C0A4B0928090",
 23590 => x"C0C0C0A4B09290C0",
 23591 => x"C0C0C0A4B09290F9",
 23592 => x"C0C0C0A4B09290A4",
 23593 => x"C0C0C0A4B09290B0",
 23594 => x"C0C0C0A4B0929099",
 23595 => x"C0C0C0A4B0929092",
 23596 => x"C0C0C0A4B0929082",
 23597 => x"C0C0C0A4B09290F8",
 23598 => x"C0C0C0A4B0929080",
 23599 => x"C0C0C0A4B0929090",
 23600 => x"C0C0C0A4B082C0C0",
 23601 => x"C0C0C0A4B082C0F9",
 23602 => x"C0C0C0A4B082C0A4",
 23603 => x"C0C0C0A4B082C0B0",
 23604 => x"C0C0C0A4B082C099",
 23605 => x"C0C0C0A4B082C092",
 23606 => x"C0C0C0A4B082C082",
 23607 => x"C0C0C0A4B082C0F8",
 23608 => x"C0C0C0A4B082C080",
 23609 => x"C0C0C0A4B082C090",
 23610 => x"C0C0C0A4B082F9C0",
 23611 => x"C0C0C0A4B082F9F9",
 23612 => x"C0C0C0A4B082F9A4",
 23613 => x"C0C0C0A4B082F9B0",
 23614 => x"C0C0C0A4B082F999",
 23615 => x"C0C0C0A4B082F992",
 23616 => x"C0C0C0A4B082F982",
 23617 => x"C0C0C0A4B082F9F8",
 23618 => x"C0C0C0A4B082F980",
 23619 => x"C0C0C0A4B082F990",
 23620 => x"C0C0C0A4B082A4C0",
 23621 => x"C0C0C0A4B082A4F9",
 23622 => x"C0C0C0A4B082A4A4",
 23623 => x"C0C0C0A4B082A4B0",
 23624 => x"C0C0C0A4B082A499",
 23625 => x"C0C0C0A4B082A492",
 23626 => x"C0C0C0A4B082A482",
 23627 => x"C0C0C0A4B082A4F8",
 23628 => x"C0C0C0A4B082A480",
 23629 => x"C0C0C0A4B082A490",
 23630 => x"C0C0C0A4B082B0C0",
 23631 => x"C0C0C0A4B082B0F9",
 23632 => x"C0C0C0A4B082B0A4",
 23633 => x"C0C0C0A4B082B0B0",
 23634 => x"C0C0C0A4B082B099",
 23635 => x"C0C0C0A4B082B092",
 23636 => x"C0C0C0A4B082B082",
 23637 => x"C0C0C0A4B082B0F8",
 23638 => x"C0C0C0A4B082B080",
 23639 => x"C0C0C0A4B082B090",
 23640 => x"C0C0C0A4B08299C0",
 23641 => x"C0C0C0A4B08299F9",
 23642 => x"C0C0C0A4B08299A4",
 23643 => x"C0C0C0A4B08299B0",
 23644 => x"C0C0C0A4B0829999",
 23645 => x"C0C0C0A4B0829992",
 23646 => x"C0C0C0A4B0829982",
 23647 => x"C0C0C0A4B08299F8",
 23648 => x"C0C0C0A4B0829980",
 23649 => x"C0C0C0A4B0829990",
 23650 => x"C0C0C0A4B08292C0",
 23651 => x"C0C0C0A4B08292F9",
 23652 => x"C0C0C0A4B08292A4",
 23653 => x"C0C0C0A4B08292B0",
 23654 => x"C0C0C0A4B0829299",
 23655 => x"C0C0C0A4B0829292",
 23656 => x"C0C0C0A4B0829282",
 23657 => x"C0C0C0A4B08292F8",
 23658 => x"C0C0C0A4B0829280",
 23659 => x"C0C0C0A4B0829290",
 23660 => x"C0C0C0A4B08282C0",
 23661 => x"C0C0C0A4B08282F9",
 23662 => x"C0C0C0A4B08282A4",
 23663 => x"C0C0C0A4B08282B0",
 23664 => x"C0C0C0A4B0828299",
 23665 => x"C0C0C0A4B0828292",
 23666 => x"C0C0C0A4B0828282",
 23667 => x"C0C0C0A4B08282F8",
 23668 => x"C0C0C0A4B0828280",
 23669 => x"C0C0C0A4B0828290",
 23670 => x"C0C0C0A4B082F8C0",
 23671 => x"C0C0C0A4B082F8F9",
 23672 => x"C0C0C0A4B082F8A4",
 23673 => x"C0C0C0A4B082F8B0",
 23674 => x"C0C0C0A4B082F899",
 23675 => x"C0C0C0A4B082F892",
 23676 => x"C0C0C0A4B082F882",
 23677 => x"C0C0C0A4B082F8F8",
 23678 => x"C0C0C0A4B082F880",
 23679 => x"C0C0C0A4B082F890",
 23680 => x"C0C0C0A4B08280C0",
 23681 => x"C0C0C0A4B08280F9",
 23682 => x"C0C0C0A4B08280A4",
 23683 => x"C0C0C0A4B08280B0",
 23684 => x"C0C0C0A4B0828099",
 23685 => x"C0C0C0A4B0828092",
 23686 => x"C0C0C0A4B0828082",
 23687 => x"C0C0C0A4B08280F8",
 23688 => x"C0C0C0A4B0828080",
 23689 => x"C0C0C0A4B0828090",
 23690 => x"C0C0C0A4B08290C0",
 23691 => x"C0C0C0A4B08290F9",
 23692 => x"C0C0C0A4B08290A4",
 23693 => x"C0C0C0A4B08290B0",
 23694 => x"C0C0C0A4B0829099",
 23695 => x"C0C0C0A4B0829092",
 23696 => x"C0C0C0A4B0829082",
 23697 => x"C0C0C0A4B08290F8",
 23698 => x"C0C0C0A4B0829080",
 23699 => x"C0C0C0A4B0829090",
 23700 => x"C0C0C0A4B0F8C0C0",
 23701 => x"C0C0C0A4B0F8C0F9",
 23702 => x"C0C0C0A4B0F8C0A4",
 23703 => x"C0C0C0A4B0F8C0B0",
 23704 => x"C0C0C0A4B0F8C099",
 23705 => x"C0C0C0A4B0F8C092",
 23706 => x"C0C0C0A4B0F8C082",
 23707 => x"C0C0C0A4B0F8C0F8",
 23708 => x"C0C0C0A4B0F8C080",
 23709 => x"C0C0C0A4B0F8C090",
 23710 => x"C0C0C0A4B0F8F9C0",
 23711 => x"C0C0C0A4B0F8F9F9",
 23712 => x"C0C0C0A4B0F8F9A4",
 23713 => x"C0C0C0A4B0F8F9B0",
 23714 => x"C0C0C0A4B0F8F999",
 23715 => x"C0C0C0A4B0F8F992",
 23716 => x"C0C0C0A4B0F8F982",
 23717 => x"C0C0C0A4B0F8F9F8",
 23718 => x"C0C0C0A4B0F8F980",
 23719 => x"C0C0C0A4B0F8F990",
 23720 => x"C0C0C0A4B0F8A4C0",
 23721 => x"C0C0C0A4B0F8A4F9",
 23722 => x"C0C0C0A4B0F8A4A4",
 23723 => x"C0C0C0A4B0F8A4B0",
 23724 => x"C0C0C0A4B0F8A499",
 23725 => x"C0C0C0A4B0F8A492",
 23726 => x"C0C0C0A4B0F8A482",
 23727 => x"C0C0C0A4B0F8A4F8",
 23728 => x"C0C0C0A4B0F8A480",
 23729 => x"C0C0C0A4B0F8A490",
 23730 => x"C0C0C0A4B0F8B0C0",
 23731 => x"C0C0C0A4B0F8B0F9",
 23732 => x"C0C0C0A4B0F8B0A4",
 23733 => x"C0C0C0A4B0F8B0B0",
 23734 => x"C0C0C0A4B0F8B099",
 23735 => x"C0C0C0A4B0F8B092",
 23736 => x"C0C0C0A4B0F8B082",
 23737 => x"C0C0C0A4B0F8B0F8",
 23738 => x"C0C0C0A4B0F8B080",
 23739 => x"C0C0C0A4B0F8B090",
 23740 => x"C0C0C0A4B0F899C0",
 23741 => x"C0C0C0A4B0F899F9",
 23742 => x"C0C0C0A4B0F899A4",
 23743 => x"C0C0C0A4B0F899B0",
 23744 => x"C0C0C0A4B0F89999",
 23745 => x"C0C0C0A4B0F89992",
 23746 => x"C0C0C0A4B0F89982",
 23747 => x"C0C0C0A4B0F899F8",
 23748 => x"C0C0C0A4B0F89980",
 23749 => x"C0C0C0A4B0F89990",
 23750 => x"C0C0C0A4B0F892C0",
 23751 => x"C0C0C0A4B0F892F9",
 23752 => x"C0C0C0A4B0F892A4",
 23753 => x"C0C0C0A4B0F892B0",
 23754 => x"C0C0C0A4B0F89299",
 23755 => x"C0C0C0A4B0F89292",
 23756 => x"C0C0C0A4B0F89282",
 23757 => x"C0C0C0A4B0F892F8",
 23758 => x"C0C0C0A4B0F89280",
 23759 => x"C0C0C0A4B0F89290",
 23760 => x"C0C0C0A4B0F882C0",
 23761 => x"C0C0C0A4B0F882F9",
 23762 => x"C0C0C0A4B0F882A4",
 23763 => x"C0C0C0A4B0F882B0",
 23764 => x"C0C0C0A4B0F88299",
 23765 => x"C0C0C0A4B0F88292",
 23766 => x"C0C0C0A4B0F88282",
 23767 => x"C0C0C0A4B0F882F8",
 23768 => x"C0C0C0A4B0F88280",
 23769 => x"C0C0C0A4B0F88290",
 23770 => x"C0C0C0A4B0F8F8C0",
 23771 => x"C0C0C0A4B0F8F8F9",
 23772 => x"C0C0C0A4B0F8F8A4",
 23773 => x"C0C0C0A4B0F8F8B0",
 23774 => x"C0C0C0A4B0F8F899",
 23775 => x"C0C0C0A4B0F8F892",
 23776 => x"C0C0C0A4B0F8F882",
 23777 => x"C0C0C0A4B0F8F8F8",
 23778 => x"C0C0C0A4B0F8F880",
 23779 => x"C0C0C0A4B0F8F890",
 23780 => x"C0C0C0A4B0F880C0",
 23781 => x"C0C0C0A4B0F880F9",
 23782 => x"C0C0C0A4B0F880A4",
 23783 => x"C0C0C0A4B0F880B0",
 23784 => x"C0C0C0A4B0F88099",
 23785 => x"C0C0C0A4B0F88092",
 23786 => x"C0C0C0A4B0F88082",
 23787 => x"C0C0C0A4B0F880F8",
 23788 => x"C0C0C0A4B0F88080",
 23789 => x"C0C0C0A4B0F88090",
 23790 => x"C0C0C0A4B0F890C0",
 23791 => x"C0C0C0A4B0F890F9",
 23792 => x"C0C0C0A4B0F890A4",
 23793 => x"C0C0C0A4B0F890B0",
 23794 => x"C0C0C0A4B0F89099",
 23795 => x"C0C0C0A4B0F89092",
 23796 => x"C0C0C0A4B0F89082",
 23797 => x"C0C0C0A4B0F890F8",
 23798 => x"C0C0C0A4B0F89080",
 23799 => x"C0C0C0A4B0F89090",
 23800 => x"C0C0C0A4B080C0C0",
 23801 => x"C0C0C0A4B080C0F9",
 23802 => x"C0C0C0A4B080C0A4",
 23803 => x"C0C0C0A4B080C0B0",
 23804 => x"C0C0C0A4B080C099",
 23805 => x"C0C0C0A4B080C092",
 23806 => x"C0C0C0A4B080C082",
 23807 => x"C0C0C0A4B080C0F8",
 23808 => x"C0C0C0A4B080C080",
 23809 => x"C0C0C0A4B080C090",
 23810 => x"C0C0C0A4B080F9C0",
 23811 => x"C0C0C0A4B080F9F9",
 23812 => x"C0C0C0A4B080F9A4",
 23813 => x"C0C0C0A4B080F9B0",
 23814 => x"C0C0C0A4B080F999",
 23815 => x"C0C0C0A4B080F992",
 23816 => x"C0C0C0A4B080F982",
 23817 => x"C0C0C0A4B080F9F8",
 23818 => x"C0C0C0A4B080F980",
 23819 => x"C0C0C0A4B080F990",
 23820 => x"C0C0C0A4B080A4C0",
 23821 => x"C0C0C0A4B080A4F9",
 23822 => x"C0C0C0A4B080A4A4",
 23823 => x"C0C0C0A4B080A4B0",
 23824 => x"C0C0C0A4B080A499",
 23825 => x"C0C0C0A4B080A492",
 23826 => x"C0C0C0A4B080A482",
 23827 => x"C0C0C0A4B080A4F8",
 23828 => x"C0C0C0A4B080A480",
 23829 => x"C0C0C0A4B080A490",
 23830 => x"C0C0C0A4B080B0C0",
 23831 => x"C0C0C0A4B080B0F9",
 23832 => x"C0C0C0A4B080B0A4",
 23833 => x"C0C0C0A4B080B0B0",
 23834 => x"C0C0C0A4B080B099",
 23835 => x"C0C0C0A4B080B092",
 23836 => x"C0C0C0A4B080B082",
 23837 => x"C0C0C0A4B080B0F8",
 23838 => x"C0C0C0A4B080B080",
 23839 => x"C0C0C0A4B080B090",
 23840 => x"C0C0C0A4B08099C0",
 23841 => x"C0C0C0A4B08099F9",
 23842 => x"C0C0C0A4B08099A4",
 23843 => x"C0C0C0A4B08099B0",
 23844 => x"C0C0C0A4B0809999",
 23845 => x"C0C0C0A4B0809992",
 23846 => x"C0C0C0A4B0809982",
 23847 => x"C0C0C0A4B08099F8",
 23848 => x"C0C0C0A4B0809980",
 23849 => x"C0C0C0A4B0809990",
 23850 => x"C0C0C0A4B08092C0",
 23851 => x"C0C0C0A4B08092F9",
 23852 => x"C0C0C0A4B08092A4",
 23853 => x"C0C0C0A4B08092B0",
 23854 => x"C0C0C0A4B0809299",
 23855 => x"C0C0C0A4B0809292",
 23856 => x"C0C0C0A4B0809282",
 23857 => x"C0C0C0A4B08092F8",
 23858 => x"C0C0C0A4B0809280",
 23859 => x"C0C0C0A4B0809290",
 23860 => x"C0C0C0A4B08082C0",
 23861 => x"C0C0C0A4B08082F9",
 23862 => x"C0C0C0A4B08082A4",
 23863 => x"C0C0C0A4B08082B0",
 23864 => x"C0C0C0A4B0808299",
 23865 => x"C0C0C0A4B0808292",
 23866 => x"C0C0C0A4B0808282",
 23867 => x"C0C0C0A4B08082F8",
 23868 => x"C0C0C0A4B0808280",
 23869 => x"C0C0C0A4B0808290",
 23870 => x"C0C0C0A4B080F8C0",
 23871 => x"C0C0C0A4B080F8F9",
 23872 => x"C0C0C0A4B080F8A4",
 23873 => x"C0C0C0A4B080F8B0",
 23874 => x"C0C0C0A4B080F899",
 23875 => x"C0C0C0A4B080F892",
 23876 => x"C0C0C0A4B080F882",
 23877 => x"C0C0C0A4B080F8F8",
 23878 => x"C0C0C0A4B080F880",
 23879 => x"C0C0C0A4B080F890",
 23880 => x"C0C0C0A4B08080C0",
 23881 => x"C0C0C0A4B08080F9",
 23882 => x"C0C0C0A4B08080A4",
 23883 => x"C0C0C0A4B08080B0",
 23884 => x"C0C0C0A4B0808099",
 23885 => x"C0C0C0A4B0808092",
 23886 => x"C0C0C0A4B0808082",
 23887 => x"C0C0C0A4B08080F8",
 23888 => x"C0C0C0A4B0808080",
 23889 => x"C0C0C0A4B0808090",
 23890 => x"C0C0C0A4B08090C0",
 23891 => x"C0C0C0A4B08090F9",
 23892 => x"C0C0C0A4B08090A4",
 23893 => x"C0C0C0A4B08090B0",
 23894 => x"C0C0C0A4B0809099",
 23895 => x"C0C0C0A4B0809092",
 23896 => x"C0C0C0A4B0809082",
 23897 => x"C0C0C0A4B08090F8",
 23898 => x"C0C0C0A4B0809080",
 23899 => x"C0C0C0A4B0809090",
 23900 => x"C0C0C0A4B090C0C0",
 23901 => x"C0C0C0A4B090C0F9",
 23902 => x"C0C0C0A4B090C0A4",
 23903 => x"C0C0C0A4B090C0B0",
 23904 => x"C0C0C0A4B090C099",
 23905 => x"C0C0C0A4B090C092",
 23906 => x"C0C0C0A4B090C082",
 23907 => x"C0C0C0A4B090C0F8",
 23908 => x"C0C0C0A4B090C080",
 23909 => x"C0C0C0A4B090C090",
 23910 => x"C0C0C0A4B090F9C0",
 23911 => x"C0C0C0A4B090F9F9",
 23912 => x"C0C0C0A4B090F9A4",
 23913 => x"C0C0C0A4B090F9B0",
 23914 => x"C0C0C0A4B090F999",
 23915 => x"C0C0C0A4B090F992",
 23916 => x"C0C0C0A4B090F982",
 23917 => x"C0C0C0A4B090F9F8",
 23918 => x"C0C0C0A4B090F980",
 23919 => x"C0C0C0A4B090F990",
 23920 => x"C0C0C0A4B090A4C0",
 23921 => x"C0C0C0A4B090A4F9",
 23922 => x"C0C0C0A4B090A4A4",
 23923 => x"C0C0C0A4B090A4B0",
 23924 => x"C0C0C0A4B090A499",
 23925 => x"C0C0C0A4B090A492",
 23926 => x"C0C0C0A4B090A482",
 23927 => x"C0C0C0A4B090A4F8",
 23928 => x"C0C0C0A4B090A480",
 23929 => x"C0C0C0A4B090A490",
 23930 => x"C0C0C0A4B090B0C0",
 23931 => x"C0C0C0A4B090B0F9",
 23932 => x"C0C0C0A4B090B0A4",
 23933 => x"C0C0C0A4B090B0B0",
 23934 => x"C0C0C0A4B090B099",
 23935 => x"C0C0C0A4B090B092",
 23936 => x"C0C0C0A4B090B082",
 23937 => x"C0C0C0A4B090B0F8",
 23938 => x"C0C0C0A4B090B080",
 23939 => x"C0C0C0A4B090B090",
 23940 => x"C0C0C0A4B09099C0",
 23941 => x"C0C0C0A4B09099F9",
 23942 => x"C0C0C0A4B09099A4",
 23943 => x"C0C0C0A4B09099B0",
 23944 => x"C0C0C0A4B0909999",
 23945 => x"C0C0C0A4B0909992",
 23946 => x"C0C0C0A4B0909982",
 23947 => x"C0C0C0A4B09099F8",
 23948 => x"C0C0C0A4B0909980",
 23949 => x"C0C0C0A4B0909990",
 23950 => x"C0C0C0A4B09092C0",
 23951 => x"C0C0C0A4B09092F9",
 23952 => x"C0C0C0A4B09092A4",
 23953 => x"C0C0C0A4B09092B0",
 23954 => x"C0C0C0A4B0909299",
 23955 => x"C0C0C0A4B0909292",
 23956 => x"C0C0C0A4B0909282",
 23957 => x"C0C0C0A4B09092F8",
 23958 => x"C0C0C0A4B0909280",
 23959 => x"C0C0C0A4B0909290",
 23960 => x"C0C0C0A4B09082C0",
 23961 => x"C0C0C0A4B09082F9",
 23962 => x"C0C0C0A4B09082A4",
 23963 => x"C0C0C0A4B09082B0",
 23964 => x"C0C0C0A4B0908299",
 23965 => x"C0C0C0A4B0908292",
 23966 => x"C0C0C0A4B0908282",
 23967 => x"C0C0C0A4B09082F8",
 23968 => x"C0C0C0A4B0908280",
 23969 => x"C0C0C0A4B0908290",
 23970 => x"C0C0C0A4B090F8C0",
 23971 => x"C0C0C0A4B090F8F9",
 23972 => x"C0C0C0A4B090F8A4",
 23973 => x"C0C0C0A4B090F8B0",
 23974 => x"C0C0C0A4B090F899",
 23975 => x"C0C0C0A4B090F892",
 23976 => x"C0C0C0A4B090F882",
 23977 => x"C0C0C0A4B090F8F8",
 23978 => x"C0C0C0A4B090F880",
 23979 => x"C0C0C0A4B090F890",
 23980 => x"C0C0C0A4B09080C0",
 23981 => x"C0C0C0A4B09080F9",
 23982 => x"C0C0C0A4B09080A4",
 23983 => x"C0C0C0A4B09080B0",
 23984 => x"C0C0C0A4B0908099",
 23985 => x"C0C0C0A4B0908092",
 23986 => x"C0C0C0A4B0908082",
 23987 => x"C0C0C0A4B09080F8",
 23988 => x"C0C0C0A4B0908080",
 23989 => x"C0C0C0A4B0908090",
 23990 => x"C0C0C0A4B09090C0",
 23991 => x"C0C0C0A4B09090F9",
 23992 => x"C0C0C0A4B09090A4",
 23993 => x"C0C0C0A4B09090B0",
 23994 => x"C0C0C0A4B0909099",
 23995 => x"C0C0C0A4B0909092",
 23996 => x"C0C0C0A4B0909082",
 23997 => x"C0C0C0A4B09090F8",
 23998 => x"C0C0C0A4B0909080",
 23999 => x"C0C0C0A4B0909090",
 24000 => x"C0C0C0A499C0C0C0",
 24001 => x"C0C0C0A499C0C0F9",
 24002 => x"C0C0C0A499C0C0A4",
 24003 => x"C0C0C0A499C0C0B0",
 24004 => x"C0C0C0A499C0C099",
 24005 => x"C0C0C0A499C0C092",
 24006 => x"C0C0C0A499C0C082",
 24007 => x"C0C0C0A499C0C0F8",
 24008 => x"C0C0C0A499C0C080",
 24009 => x"C0C0C0A499C0C090",
 24010 => x"C0C0C0A499C0F9C0",
 24011 => x"C0C0C0A499C0F9F9",
 24012 => x"C0C0C0A499C0F9A4",
 24013 => x"C0C0C0A499C0F9B0",
 24014 => x"C0C0C0A499C0F999",
 24015 => x"C0C0C0A499C0F992",
 24016 => x"C0C0C0A499C0F982",
 24017 => x"C0C0C0A499C0F9F8",
 24018 => x"C0C0C0A499C0F980",
 24019 => x"C0C0C0A499C0F990",
 24020 => x"C0C0C0A499C0A4C0",
 24021 => x"C0C0C0A499C0A4F9",
 24022 => x"C0C0C0A499C0A4A4",
 24023 => x"C0C0C0A499C0A4B0",
 24024 => x"C0C0C0A499C0A499",
 24025 => x"C0C0C0A499C0A492",
 24026 => x"C0C0C0A499C0A482",
 24027 => x"C0C0C0A499C0A4F8",
 24028 => x"C0C0C0A499C0A480",
 24029 => x"C0C0C0A499C0A490",
 24030 => x"C0C0C0A499C0B0C0",
 24031 => x"C0C0C0A499C0B0F9",
 24032 => x"C0C0C0A499C0B0A4",
 24033 => x"C0C0C0A499C0B0B0",
 24034 => x"C0C0C0A499C0B099",
 24035 => x"C0C0C0A499C0B092",
 24036 => x"C0C0C0A499C0B082",
 24037 => x"C0C0C0A499C0B0F8",
 24038 => x"C0C0C0A499C0B080",
 24039 => x"C0C0C0A499C0B090",
 24040 => x"C0C0C0A499C099C0",
 24041 => x"C0C0C0A499C099F9",
 24042 => x"C0C0C0A499C099A4",
 24043 => x"C0C0C0A499C099B0",
 24044 => x"C0C0C0A499C09999",
 24045 => x"C0C0C0A499C09992",
 24046 => x"C0C0C0A499C09982",
 24047 => x"C0C0C0A499C099F8",
 24048 => x"C0C0C0A499C09980",
 24049 => x"C0C0C0A499C09990",
 24050 => x"C0C0C0A499C092C0",
 24051 => x"C0C0C0A499C092F9",
 24052 => x"C0C0C0A499C092A4",
 24053 => x"C0C0C0A499C092B0",
 24054 => x"C0C0C0A499C09299",
 24055 => x"C0C0C0A499C09292",
 24056 => x"C0C0C0A499C09282",
 24057 => x"C0C0C0A499C092F8",
 24058 => x"C0C0C0A499C09280",
 24059 => x"C0C0C0A499C09290",
 24060 => x"C0C0C0A499C082C0",
 24061 => x"C0C0C0A499C082F9",
 24062 => x"C0C0C0A499C082A4",
 24063 => x"C0C0C0A499C082B0",
 24064 => x"C0C0C0A499C08299",
 24065 => x"C0C0C0A499C08292",
 24066 => x"C0C0C0A499C08282",
 24067 => x"C0C0C0A499C082F8",
 24068 => x"C0C0C0A499C08280",
 24069 => x"C0C0C0A499C08290",
 24070 => x"C0C0C0A499C0F8C0",
 24071 => x"C0C0C0A499C0F8F9",
 24072 => x"C0C0C0A499C0F8A4",
 24073 => x"C0C0C0A499C0F8B0",
 24074 => x"C0C0C0A499C0F899",
 24075 => x"C0C0C0A499C0F892",
 24076 => x"C0C0C0A499C0F882",
 24077 => x"C0C0C0A499C0F8F8",
 24078 => x"C0C0C0A499C0F880",
 24079 => x"C0C0C0A499C0F890",
 24080 => x"C0C0C0A499C080C0",
 24081 => x"C0C0C0A499C080F9",
 24082 => x"C0C0C0A499C080A4",
 24083 => x"C0C0C0A499C080B0",
 24084 => x"C0C0C0A499C08099",
 24085 => x"C0C0C0A499C08092",
 24086 => x"C0C0C0A499C08082",
 24087 => x"C0C0C0A499C080F8",
 24088 => x"C0C0C0A499C08080",
 24089 => x"C0C0C0A499C08090",
 24090 => x"C0C0C0A499C090C0",
 24091 => x"C0C0C0A499C090F9",
 24092 => x"C0C0C0A499C090A4",
 24093 => x"C0C0C0A499C090B0",
 24094 => x"C0C0C0A499C09099",
 24095 => x"C0C0C0A499C09092",
 24096 => x"C0C0C0A499C09082",
 24097 => x"C0C0C0A499C090F8",
 24098 => x"C0C0C0A499C09080",
 24099 => x"C0C0C0A499C09090",
 24100 => x"C0C0C0A499F9C0C0",
 24101 => x"C0C0C0A499F9C0F9",
 24102 => x"C0C0C0A499F9C0A4",
 24103 => x"C0C0C0A499F9C0B0",
 24104 => x"C0C0C0A499F9C099",
 24105 => x"C0C0C0A499F9C092",
 24106 => x"C0C0C0A499F9C082",
 24107 => x"C0C0C0A499F9C0F8",
 24108 => x"C0C0C0A499F9C080",
 24109 => x"C0C0C0A499F9C090",
 24110 => x"C0C0C0A499F9F9C0",
 24111 => x"C0C0C0A499F9F9F9",
 24112 => x"C0C0C0A499F9F9A4",
 24113 => x"C0C0C0A499F9F9B0",
 24114 => x"C0C0C0A499F9F999",
 24115 => x"C0C0C0A499F9F992",
 24116 => x"C0C0C0A499F9F982",
 24117 => x"C0C0C0A499F9F9F8",
 24118 => x"C0C0C0A499F9F980",
 24119 => x"C0C0C0A499F9F990",
 24120 => x"C0C0C0A499F9A4C0",
 24121 => x"C0C0C0A499F9A4F9",
 24122 => x"C0C0C0A499F9A4A4",
 24123 => x"C0C0C0A499F9A4B0",
 24124 => x"C0C0C0A499F9A499",
 24125 => x"C0C0C0A499F9A492",
 24126 => x"C0C0C0A499F9A482",
 24127 => x"C0C0C0A499F9A4F8",
 24128 => x"C0C0C0A499F9A480",
 24129 => x"C0C0C0A499F9A490",
 24130 => x"C0C0C0A499F9B0C0",
 24131 => x"C0C0C0A499F9B0F9",
 24132 => x"C0C0C0A499F9B0A4",
 24133 => x"C0C0C0A499F9B0B0",
 24134 => x"C0C0C0A499F9B099",
 24135 => x"C0C0C0A499F9B092",
 24136 => x"C0C0C0A499F9B082",
 24137 => x"C0C0C0A499F9B0F8",
 24138 => x"C0C0C0A499F9B080",
 24139 => x"C0C0C0A499F9B090",
 24140 => x"C0C0C0A499F999C0",
 24141 => x"C0C0C0A499F999F9",
 24142 => x"C0C0C0A499F999A4",
 24143 => x"C0C0C0A499F999B0",
 24144 => x"C0C0C0A499F99999",
 24145 => x"C0C0C0A499F99992",
 24146 => x"C0C0C0A499F99982",
 24147 => x"C0C0C0A499F999F8",
 24148 => x"C0C0C0A499F99980",
 24149 => x"C0C0C0A499F99990",
 24150 => x"C0C0C0A499F992C0",
 24151 => x"C0C0C0A499F992F9",
 24152 => x"C0C0C0A499F992A4",
 24153 => x"C0C0C0A499F992B0",
 24154 => x"C0C0C0A499F99299",
 24155 => x"C0C0C0A499F99292",
 24156 => x"C0C0C0A499F99282",
 24157 => x"C0C0C0A499F992F8",
 24158 => x"C0C0C0A499F99280",
 24159 => x"C0C0C0A499F99290",
 24160 => x"C0C0C0A499F982C0",
 24161 => x"C0C0C0A499F982F9",
 24162 => x"C0C0C0A499F982A4",
 24163 => x"C0C0C0A499F982B0",
 24164 => x"C0C0C0A499F98299",
 24165 => x"C0C0C0A499F98292",
 24166 => x"C0C0C0A499F98282",
 24167 => x"C0C0C0A499F982F8",
 24168 => x"C0C0C0A499F98280",
 24169 => x"C0C0C0A499F98290",
 24170 => x"C0C0C0A499F9F8C0",
 24171 => x"C0C0C0A499F9F8F9",
 24172 => x"C0C0C0A499F9F8A4",
 24173 => x"C0C0C0A499F9F8B0",
 24174 => x"C0C0C0A499F9F899",
 24175 => x"C0C0C0A499F9F892",
 24176 => x"C0C0C0A499F9F882",
 24177 => x"C0C0C0A499F9F8F8",
 24178 => x"C0C0C0A499F9F880",
 24179 => x"C0C0C0A499F9F890",
 24180 => x"C0C0C0A499F980C0",
 24181 => x"C0C0C0A499F980F9",
 24182 => x"C0C0C0A499F980A4",
 24183 => x"C0C0C0A499F980B0",
 24184 => x"C0C0C0A499F98099",
 24185 => x"C0C0C0A499F98092",
 24186 => x"C0C0C0A499F98082",
 24187 => x"C0C0C0A499F980F8",
 24188 => x"C0C0C0A499F98080",
 24189 => x"C0C0C0A499F98090",
 24190 => x"C0C0C0A499F990C0",
 24191 => x"C0C0C0A499F990F9",
 24192 => x"C0C0C0A499F990A4",
 24193 => x"C0C0C0A499F990B0",
 24194 => x"C0C0C0A499F99099",
 24195 => x"C0C0C0A499F99092",
 24196 => x"C0C0C0A499F99082",
 24197 => x"C0C0C0A499F990F8",
 24198 => x"C0C0C0A499F99080",
 24199 => x"C0C0C0A499F99090",
 24200 => x"C0C0C0A499A4C0C0",
 24201 => x"C0C0C0A499A4C0F9",
 24202 => x"C0C0C0A499A4C0A4",
 24203 => x"C0C0C0A499A4C0B0",
 24204 => x"C0C0C0A499A4C099",
 24205 => x"C0C0C0A499A4C092",
 24206 => x"C0C0C0A499A4C082",
 24207 => x"C0C0C0A499A4C0F8",
 24208 => x"C0C0C0A499A4C080",
 24209 => x"C0C0C0A499A4C090",
 24210 => x"C0C0C0A499A4F9C0",
 24211 => x"C0C0C0A499A4F9F9",
 24212 => x"C0C0C0A499A4F9A4",
 24213 => x"C0C0C0A499A4F9B0",
 24214 => x"C0C0C0A499A4F999",
 24215 => x"C0C0C0A499A4F992",
 24216 => x"C0C0C0A499A4F982",
 24217 => x"C0C0C0A499A4F9F8",
 24218 => x"C0C0C0A499A4F980",
 24219 => x"C0C0C0A499A4F990",
 24220 => x"C0C0C0A499A4A4C0",
 24221 => x"C0C0C0A499A4A4F9",
 24222 => x"C0C0C0A499A4A4A4",
 24223 => x"C0C0C0A499A4A4B0",
 24224 => x"C0C0C0A499A4A499",
 24225 => x"C0C0C0A499A4A492",
 24226 => x"C0C0C0A499A4A482",
 24227 => x"C0C0C0A499A4A4F8",
 24228 => x"C0C0C0A499A4A480",
 24229 => x"C0C0C0A499A4A490",
 24230 => x"C0C0C0A499A4B0C0",
 24231 => x"C0C0C0A499A4B0F9",
 24232 => x"C0C0C0A499A4B0A4",
 24233 => x"C0C0C0A499A4B0B0",
 24234 => x"C0C0C0A499A4B099",
 24235 => x"C0C0C0A499A4B092",
 24236 => x"C0C0C0A499A4B082",
 24237 => x"C0C0C0A499A4B0F8",
 24238 => x"C0C0C0A499A4B080",
 24239 => x"C0C0C0A499A4B090",
 24240 => x"C0C0C0A499A499C0",
 24241 => x"C0C0C0A499A499F9",
 24242 => x"C0C0C0A499A499A4",
 24243 => x"C0C0C0A499A499B0",
 24244 => x"C0C0C0A499A49999",
 24245 => x"C0C0C0A499A49992",
 24246 => x"C0C0C0A499A49982",
 24247 => x"C0C0C0A499A499F8",
 24248 => x"C0C0C0A499A49980",
 24249 => x"C0C0C0A499A49990",
 24250 => x"C0C0C0A499A492C0",
 24251 => x"C0C0C0A499A492F9",
 24252 => x"C0C0C0A499A492A4",
 24253 => x"C0C0C0A499A492B0",
 24254 => x"C0C0C0A499A49299",
 24255 => x"C0C0C0A499A49292",
 24256 => x"C0C0C0A499A49282",
 24257 => x"C0C0C0A499A492F8",
 24258 => x"C0C0C0A499A49280",
 24259 => x"C0C0C0A499A49290",
 24260 => x"C0C0C0A499A482C0",
 24261 => x"C0C0C0A499A482F9",
 24262 => x"C0C0C0A499A482A4",
 24263 => x"C0C0C0A499A482B0",
 24264 => x"C0C0C0A499A48299",
 24265 => x"C0C0C0A499A48292",
 24266 => x"C0C0C0A499A48282",
 24267 => x"C0C0C0A499A482F8",
 24268 => x"C0C0C0A499A48280",
 24269 => x"C0C0C0A499A48290",
 24270 => x"C0C0C0A499A4F8C0",
 24271 => x"C0C0C0A499A4F8F9",
 24272 => x"C0C0C0A499A4F8A4",
 24273 => x"C0C0C0A499A4F8B0",
 24274 => x"C0C0C0A499A4F899",
 24275 => x"C0C0C0A499A4F892",
 24276 => x"C0C0C0A499A4F882",
 24277 => x"C0C0C0A499A4F8F8",
 24278 => x"C0C0C0A499A4F880",
 24279 => x"C0C0C0A499A4F890",
 24280 => x"C0C0C0A499A480C0",
 24281 => x"C0C0C0A499A480F9",
 24282 => x"C0C0C0A499A480A4",
 24283 => x"C0C0C0A499A480B0",
 24284 => x"C0C0C0A499A48099",
 24285 => x"C0C0C0A499A48092",
 24286 => x"C0C0C0A499A48082",
 24287 => x"C0C0C0A499A480F8",
 24288 => x"C0C0C0A499A48080",
 24289 => x"C0C0C0A499A48090",
 24290 => x"C0C0C0A499A490C0",
 24291 => x"C0C0C0A499A490F9",
 24292 => x"C0C0C0A499A490A4",
 24293 => x"C0C0C0A499A490B0",
 24294 => x"C0C0C0A499A49099",
 24295 => x"C0C0C0A499A49092",
 24296 => x"C0C0C0A499A49082",
 24297 => x"C0C0C0A499A490F8",
 24298 => x"C0C0C0A499A49080",
 24299 => x"C0C0C0A499A49090",
 24300 => x"C0C0C0A499B0C0C0",
 24301 => x"C0C0C0A499B0C0F9",
 24302 => x"C0C0C0A499B0C0A4",
 24303 => x"C0C0C0A499B0C0B0",
 24304 => x"C0C0C0A499B0C099",
 24305 => x"C0C0C0A499B0C092",
 24306 => x"C0C0C0A499B0C082",
 24307 => x"C0C0C0A499B0C0F8",
 24308 => x"C0C0C0A499B0C080",
 24309 => x"C0C0C0A499B0C090",
 24310 => x"C0C0C0A499B0F9C0",
 24311 => x"C0C0C0A499B0F9F9",
 24312 => x"C0C0C0A499B0F9A4",
 24313 => x"C0C0C0A499B0F9B0",
 24314 => x"C0C0C0A499B0F999",
 24315 => x"C0C0C0A499B0F992",
 24316 => x"C0C0C0A499B0F982",
 24317 => x"C0C0C0A499B0F9F8",
 24318 => x"C0C0C0A499B0F980",
 24319 => x"C0C0C0A499B0F990",
 24320 => x"C0C0C0A499B0A4C0",
 24321 => x"C0C0C0A499B0A4F9",
 24322 => x"C0C0C0A499B0A4A4",
 24323 => x"C0C0C0A499B0A4B0",
 24324 => x"C0C0C0A499B0A499",
 24325 => x"C0C0C0A499B0A492",
 24326 => x"C0C0C0A499B0A482",
 24327 => x"C0C0C0A499B0A4F8",
 24328 => x"C0C0C0A499B0A480",
 24329 => x"C0C0C0A499B0A490",
 24330 => x"C0C0C0A499B0B0C0",
 24331 => x"C0C0C0A499B0B0F9",
 24332 => x"C0C0C0A499B0B0A4",
 24333 => x"C0C0C0A499B0B0B0",
 24334 => x"C0C0C0A499B0B099",
 24335 => x"C0C0C0A499B0B092",
 24336 => x"C0C0C0A499B0B082",
 24337 => x"C0C0C0A499B0B0F8",
 24338 => x"C0C0C0A499B0B080",
 24339 => x"C0C0C0A499B0B090",
 24340 => x"C0C0C0A499B099C0",
 24341 => x"C0C0C0A499B099F9",
 24342 => x"C0C0C0A499B099A4",
 24343 => x"C0C0C0A499B099B0",
 24344 => x"C0C0C0A499B09999",
 24345 => x"C0C0C0A499B09992",
 24346 => x"C0C0C0A499B09982",
 24347 => x"C0C0C0A499B099F8",
 24348 => x"C0C0C0A499B09980",
 24349 => x"C0C0C0A499B09990",
 24350 => x"C0C0C0A499B092C0",
 24351 => x"C0C0C0A499B092F9",
 24352 => x"C0C0C0A499B092A4",
 24353 => x"C0C0C0A499B092B0",
 24354 => x"C0C0C0A499B09299",
 24355 => x"C0C0C0A499B09292",
 24356 => x"C0C0C0A499B09282",
 24357 => x"C0C0C0A499B092F8",
 24358 => x"C0C0C0A499B09280",
 24359 => x"C0C0C0A499B09290",
 24360 => x"C0C0C0A499B082C0",
 24361 => x"C0C0C0A499B082F9",
 24362 => x"C0C0C0A499B082A4",
 24363 => x"C0C0C0A499B082B0",
 24364 => x"C0C0C0A499B08299",
 24365 => x"C0C0C0A499B08292",
 24366 => x"C0C0C0A499B08282",
 24367 => x"C0C0C0A499B082F8",
 24368 => x"C0C0C0A499B08280",
 24369 => x"C0C0C0A499B08290",
 24370 => x"C0C0C0A499B0F8C0",
 24371 => x"C0C0C0A499B0F8F9",
 24372 => x"C0C0C0A499B0F8A4",
 24373 => x"C0C0C0A499B0F8B0",
 24374 => x"C0C0C0A499B0F899",
 24375 => x"C0C0C0A499B0F892",
 24376 => x"C0C0C0A499B0F882",
 24377 => x"C0C0C0A499B0F8F8",
 24378 => x"C0C0C0A499B0F880",
 24379 => x"C0C0C0A499B0F890",
 24380 => x"C0C0C0A499B080C0",
 24381 => x"C0C0C0A499B080F9",
 24382 => x"C0C0C0A499B080A4",
 24383 => x"C0C0C0A499B080B0",
 24384 => x"C0C0C0A499B08099",
 24385 => x"C0C0C0A499B08092",
 24386 => x"C0C0C0A499B08082",
 24387 => x"C0C0C0A499B080F8",
 24388 => x"C0C0C0A499B08080",
 24389 => x"C0C0C0A499B08090",
 24390 => x"C0C0C0A499B090C0",
 24391 => x"C0C0C0A499B090F9",
 24392 => x"C0C0C0A499B090A4",
 24393 => x"C0C0C0A499B090B0",
 24394 => x"C0C0C0A499B09099",
 24395 => x"C0C0C0A499B09092",
 24396 => x"C0C0C0A499B09082",
 24397 => x"C0C0C0A499B090F8",
 24398 => x"C0C0C0A499B09080",
 24399 => x"C0C0C0A499B09090",
 24400 => x"C0C0C0A49999C0C0",
 24401 => x"C0C0C0A49999C0F9",
 24402 => x"C0C0C0A49999C0A4",
 24403 => x"C0C0C0A49999C0B0",
 24404 => x"C0C0C0A49999C099",
 24405 => x"C0C0C0A49999C092",
 24406 => x"C0C0C0A49999C082",
 24407 => x"C0C0C0A49999C0F8",
 24408 => x"C0C0C0A49999C080",
 24409 => x"C0C0C0A49999C090",
 24410 => x"C0C0C0A49999F9C0",
 24411 => x"C0C0C0A49999F9F9",
 24412 => x"C0C0C0A49999F9A4",
 24413 => x"C0C0C0A49999F9B0",
 24414 => x"C0C0C0A49999F999",
 24415 => x"C0C0C0A49999F992",
 24416 => x"C0C0C0A49999F982",
 24417 => x"C0C0C0A49999F9F8",
 24418 => x"C0C0C0A49999F980",
 24419 => x"C0C0C0A49999F990",
 24420 => x"C0C0C0A49999A4C0",
 24421 => x"C0C0C0A49999A4F9",
 24422 => x"C0C0C0A49999A4A4",
 24423 => x"C0C0C0A49999A4B0",
 24424 => x"C0C0C0A49999A499",
 24425 => x"C0C0C0A49999A492",
 24426 => x"C0C0C0A49999A482",
 24427 => x"C0C0C0A49999A4F8",
 24428 => x"C0C0C0A49999A480",
 24429 => x"C0C0C0A49999A490",
 24430 => x"C0C0C0A49999B0C0",
 24431 => x"C0C0C0A49999B0F9",
 24432 => x"C0C0C0A49999B0A4",
 24433 => x"C0C0C0A49999B0B0",
 24434 => x"C0C0C0A49999B099",
 24435 => x"C0C0C0A49999B092",
 24436 => x"C0C0C0A49999B082",
 24437 => x"C0C0C0A49999B0F8",
 24438 => x"C0C0C0A49999B080",
 24439 => x"C0C0C0A49999B090",
 24440 => x"C0C0C0A4999999C0",
 24441 => x"C0C0C0A4999999F9",
 24442 => x"C0C0C0A4999999A4",
 24443 => x"C0C0C0A4999999B0",
 24444 => x"C0C0C0A499999999",
 24445 => x"C0C0C0A499999992",
 24446 => x"C0C0C0A499999982",
 24447 => x"C0C0C0A4999999F8",
 24448 => x"C0C0C0A499999980",
 24449 => x"C0C0C0A499999990",
 24450 => x"C0C0C0A4999992C0",
 24451 => x"C0C0C0A4999992F9",
 24452 => x"C0C0C0A4999992A4",
 24453 => x"C0C0C0A4999992B0",
 24454 => x"C0C0C0A499999299",
 24455 => x"C0C0C0A499999292",
 24456 => x"C0C0C0A499999282",
 24457 => x"C0C0C0A4999992F8",
 24458 => x"C0C0C0A499999280",
 24459 => x"C0C0C0A499999290",
 24460 => x"C0C0C0A4999982C0",
 24461 => x"C0C0C0A4999982F9",
 24462 => x"C0C0C0A4999982A4",
 24463 => x"C0C0C0A4999982B0",
 24464 => x"C0C0C0A499998299",
 24465 => x"C0C0C0A499998292",
 24466 => x"C0C0C0A499998282",
 24467 => x"C0C0C0A4999982F8",
 24468 => x"C0C0C0A499998280",
 24469 => x"C0C0C0A499998290",
 24470 => x"C0C0C0A49999F8C0",
 24471 => x"C0C0C0A49999F8F9",
 24472 => x"C0C0C0A49999F8A4",
 24473 => x"C0C0C0A49999F8B0",
 24474 => x"C0C0C0A49999F899",
 24475 => x"C0C0C0A49999F892",
 24476 => x"C0C0C0A49999F882",
 24477 => x"C0C0C0A49999F8F8",
 24478 => x"C0C0C0A49999F880",
 24479 => x"C0C0C0A49999F890",
 24480 => x"C0C0C0A4999980C0",
 24481 => x"C0C0C0A4999980F9",
 24482 => x"C0C0C0A4999980A4",
 24483 => x"C0C0C0A4999980B0",
 24484 => x"C0C0C0A499998099",
 24485 => x"C0C0C0A499998092",
 24486 => x"C0C0C0A499998082",
 24487 => x"C0C0C0A4999980F8",
 24488 => x"C0C0C0A499998080",
 24489 => x"C0C0C0A499998090",
 24490 => x"C0C0C0A4999990C0",
 24491 => x"C0C0C0A4999990F9",
 24492 => x"C0C0C0A4999990A4",
 24493 => x"C0C0C0A4999990B0",
 24494 => x"C0C0C0A499999099",
 24495 => x"C0C0C0A499999092",
 24496 => x"C0C0C0A499999082",
 24497 => x"C0C0C0A4999990F8",
 24498 => x"C0C0C0A499999080",
 24499 => x"C0C0C0A499999090",
 24500 => x"C0C0C0A49992C0C0",
 24501 => x"C0C0C0A49992C0F9",
 24502 => x"C0C0C0A49992C0A4",
 24503 => x"C0C0C0A49992C0B0",
 24504 => x"C0C0C0A49992C099",
 24505 => x"C0C0C0A49992C092",
 24506 => x"C0C0C0A49992C082",
 24507 => x"C0C0C0A49992C0F8",
 24508 => x"C0C0C0A49992C080",
 24509 => x"C0C0C0A49992C090",
 24510 => x"C0C0C0A49992F9C0",
 24511 => x"C0C0C0A49992F9F9",
 24512 => x"C0C0C0A49992F9A4",
 24513 => x"C0C0C0A49992F9B0",
 24514 => x"C0C0C0A49992F999",
 24515 => x"C0C0C0A49992F992",
 24516 => x"C0C0C0A49992F982",
 24517 => x"C0C0C0A49992F9F8",
 24518 => x"C0C0C0A49992F980",
 24519 => x"C0C0C0A49992F990",
 24520 => x"C0C0C0A49992A4C0",
 24521 => x"C0C0C0A49992A4F9",
 24522 => x"C0C0C0A49992A4A4",
 24523 => x"C0C0C0A49992A4B0",
 24524 => x"C0C0C0A49992A499",
 24525 => x"C0C0C0A49992A492",
 24526 => x"C0C0C0A49992A482",
 24527 => x"C0C0C0A49992A4F8",
 24528 => x"C0C0C0A49992A480",
 24529 => x"C0C0C0A49992A490",
 24530 => x"C0C0C0A49992B0C0",
 24531 => x"C0C0C0A49992B0F9",
 24532 => x"C0C0C0A49992B0A4",
 24533 => x"C0C0C0A49992B0B0",
 24534 => x"C0C0C0A49992B099",
 24535 => x"C0C0C0A49992B092",
 24536 => x"C0C0C0A49992B082",
 24537 => x"C0C0C0A49992B0F8",
 24538 => x"C0C0C0A49992B080",
 24539 => x"C0C0C0A49992B090",
 24540 => x"C0C0C0A4999299C0",
 24541 => x"C0C0C0A4999299F9",
 24542 => x"C0C0C0A4999299A4",
 24543 => x"C0C0C0A4999299B0",
 24544 => x"C0C0C0A499929999",
 24545 => x"C0C0C0A499929992",
 24546 => x"C0C0C0A499929982",
 24547 => x"C0C0C0A4999299F8",
 24548 => x"C0C0C0A499929980",
 24549 => x"C0C0C0A499929990",
 24550 => x"C0C0C0A4999292C0",
 24551 => x"C0C0C0A4999292F9",
 24552 => x"C0C0C0A4999292A4",
 24553 => x"C0C0C0A4999292B0",
 24554 => x"C0C0C0A499929299",
 24555 => x"C0C0C0A499929292",
 24556 => x"C0C0C0A499929282",
 24557 => x"C0C0C0A4999292F8",
 24558 => x"C0C0C0A499929280",
 24559 => x"C0C0C0A499929290",
 24560 => x"C0C0C0A4999282C0",
 24561 => x"C0C0C0A4999282F9",
 24562 => x"C0C0C0A4999282A4",
 24563 => x"C0C0C0A4999282B0",
 24564 => x"C0C0C0A499928299",
 24565 => x"C0C0C0A499928292",
 24566 => x"C0C0C0A499928282",
 24567 => x"C0C0C0A4999282F8",
 24568 => x"C0C0C0A499928280",
 24569 => x"C0C0C0A499928290",
 24570 => x"C0C0C0A49992F8C0",
 24571 => x"C0C0C0A49992F8F9",
 24572 => x"C0C0C0A49992F8A4",
 24573 => x"C0C0C0A49992F8B0",
 24574 => x"C0C0C0A49992F899",
 24575 => x"C0C0C0A49992F892",
 24576 => x"C0C0C0A49992F882",
 24577 => x"C0C0C0A49992F8F8",
 24578 => x"C0C0C0A49992F880",
 24579 => x"C0C0C0A49992F890",
 24580 => x"C0C0C0A4999280C0",
 24581 => x"C0C0C0A4999280F9",
 24582 => x"C0C0C0A4999280A4",
 24583 => x"C0C0C0A4999280B0",
 24584 => x"C0C0C0A499928099",
 24585 => x"C0C0C0A499928092",
 24586 => x"C0C0C0A499928082",
 24587 => x"C0C0C0A4999280F8",
 24588 => x"C0C0C0A499928080",
 24589 => x"C0C0C0A499928090",
 24590 => x"C0C0C0A4999290C0",
 24591 => x"C0C0C0A4999290F9",
 24592 => x"C0C0C0A4999290A4",
 24593 => x"C0C0C0A4999290B0",
 24594 => x"C0C0C0A499929099",
 24595 => x"C0C0C0A499929092",
 24596 => x"C0C0C0A499929082",
 24597 => x"C0C0C0A4999290F8",
 24598 => x"C0C0C0A499929080",
 24599 => x"C0C0C0A499929090",
 24600 => x"C0C0C0A49982C0C0",
 24601 => x"C0C0C0A49982C0F9",
 24602 => x"C0C0C0A49982C0A4",
 24603 => x"C0C0C0A49982C0B0",
 24604 => x"C0C0C0A49982C099",
 24605 => x"C0C0C0A49982C092",
 24606 => x"C0C0C0A49982C082",
 24607 => x"C0C0C0A49982C0F8",
 24608 => x"C0C0C0A49982C080",
 24609 => x"C0C0C0A49982C090",
 24610 => x"C0C0C0A49982F9C0",
 24611 => x"C0C0C0A49982F9F9",
 24612 => x"C0C0C0A49982F9A4",
 24613 => x"C0C0C0A49982F9B0",
 24614 => x"C0C0C0A49982F999",
 24615 => x"C0C0C0A49982F992",
 24616 => x"C0C0C0A49982F982",
 24617 => x"C0C0C0A49982F9F8",
 24618 => x"C0C0C0A49982F980",
 24619 => x"C0C0C0A49982F990",
 24620 => x"C0C0C0A49982A4C0",
 24621 => x"C0C0C0A49982A4F9",
 24622 => x"C0C0C0A49982A4A4",
 24623 => x"C0C0C0A49982A4B0",
 24624 => x"C0C0C0A49982A499",
 24625 => x"C0C0C0A49982A492",
 24626 => x"C0C0C0A49982A482",
 24627 => x"C0C0C0A49982A4F8",
 24628 => x"C0C0C0A49982A480",
 24629 => x"C0C0C0A49982A490",
 24630 => x"C0C0C0A49982B0C0",
 24631 => x"C0C0C0A49982B0F9",
 24632 => x"C0C0C0A49982B0A4",
 24633 => x"C0C0C0A49982B0B0",
 24634 => x"C0C0C0A49982B099",
 24635 => x"C0C0C0A49982B092",
 24636 => x"C0C0C0A49982B082",
 24637 => x"C0C0C0A49982B0F8",
 24638 => x"C0C0C0A49982B080",
 24639 => x"C0C0C0A49982B090",
 24640 => x"C0C0C0A4998299C0",
 24641 => x"C0C0C0A4998299F9",
 24642 => x"C0C0C0A4998299A4",
 24643 => x"C0C0C0A4998299B0",
 24644 => x"C0C0C0A499829999",
 24645 => x"C0C0C0A499829992",
 24646 => x"C0C0C0A499829982",
 24647 => x"C0C0C0A4998299F8",
 24648 => x"C0C0C0A499829980",
 24649 => x"C0C0C0A499829990",
 24650 => x"C0C0C0A4998292C0",
 24651 => x"C0C0C0A4998292F9",
 24652 => x"C0C0C0A4998292A4",
 24653 => x"C0C0C0A4998292B0",
 24654 => x"C0C0C0A499829299",
 24655 => x"C0C0C0A499829292",
 24656 => x"C0C0C0A499829282",
 24657 => x"C0C0C0A4998292F8",
 24658 => x"C0C0C0A499829280",
 24659 => x"C0C0C0A499829290",
 24660 => x"C0C0C0A4998282C0",
 24661 => x"C0C0C0A4998282F9",
 24662 => x"C0C0C0A4998282A4",
 24663 => x"C0C0C0A4998282B0",
 24664 => x"C0C0C0A499828299",
 24665 => x"C0C0C0A499828292",
 24666 => x"C0C0C0A499828282",
 24667 => x"C0C0C0A4998282F8",
 24668 => x"C0C0C0A499828280",
 24669 => x"C0C0C0A499828290",
 24670 => x"C0C0C0A49982F8C0",
 24671 => x"C0C0C0A49982F8F9",
 24672 => x"C0C0C0A49982F8A4",
 24673 => x"C0C0C0A49982F8B0",
 24674 => x"C0C0C0A49982F899",
 24675 => x"C0C0C0A49982F892",
 24676 => x"C0C0C0A49982F882",
 24677 => x"C0C0C0A49982F8F8",
 24678 => x"C0C0C0A49982F880",
 24679 => x"C0C0C0A49982F890",
 24680 => x"C0C0C0A4998280C0",
 24681 => x"C0C0C0A4998280F9",
 24682 => x"C0C0C0A4998280A4",
 24683 => x"C0C0C0A4998280B0",
 24684 => x"C0C0C0A499828099",
 24685 => x"C0C0C0A499828092",
 24686 => x"C0C0C0A499828082",
 24687 => x"C0C0C0A4998280F8",
 24688 => x"C0C0C0A499828080",
 24689 => x"C0C0C0A499828090",
 24690 => x"C0C0C0A4998290C0",
 24691 => x"C0C0C0A4998290F9",
 24692 => x"C0C0C0A4998290A4",
 24693 => x"C0C0C0A4998290B0",
 24694 => x"C0C0C0A499829099",
 24695 => x"C0C0C0A499829092",
 24696 => x"C0C0C0A499829082",
 24697 => x"C0C0C0A4998290F8",
 24698 => x"C0C0C0A499829080",
 24699 => x"C0C0C0A499829090",
 24700 => x"C0C0C0A499F8C0C0",
 24701 => x"C0C0C0A499F8C0F9",
 24702 => x"C0C0C0A499F8C0A4",
 24703 => x"C0C0C0A499F8C0B0",
 24704 => x"C0C0C0A499F8C099",
 24705 => x"C0C0C0A499F8C092",
 24706 => x"C0C0C0A499F8C082",
 24707 => x"C0C0C0A499F8C0F8",
 24708 => x"C0C0C0A499F8C080",
 24709 => x"C0C0C0A499F8C090",
 24710 => x"C0C0C0A499F8F9C0",
 24711 => x"C0C0C0A499F8F9F9",
 24712 => x"C0C0C0A499F8F9A4",
 24713 => x"C0C0C0A499F8F9B0",
 24714 => x"C0C0C0A499F8F999",
 24715 => x"C0C0C0A499F8F992",
 24716 => x"C0C0C0A499F8F982",
 24717 => x"C0C0C0A499F8F9F8",
 24718 => x"C0C0C0A499F8F980",
 24719 => x"C0C0C0A499F8F990",
 24720 => x"C0C0C0A499F8A4C0",
 24721 => x"C0C0C0A499F8A4F9",
 24722 => x"C0C0C0A499F8A4A4",
 24723 => x"C0C0C0A499F8A4B0",
 24724 => x"C0C0C0A499F8A499",
 24725 => x"C0C0C0A499F8A492",
 24726 => x"C0C0C0A499F8A482",
 24727 => x"C0C0C0A499F8A4F8",
 24728 => x"C0C0C0A499F8A480",
 24729 => x"C0C0C0A499F8A490",
 24730 => x"C0C0C0A499F8B0C0",
 24731 => x"C0C0C0A499F8B0F9",
 24732 => x"C0C0C0A499F8B0A4",
 24733 => x"C0C0C0A499F8B0B0",
 24734 => x"C0C0C0A499F8B099",
 24735 => x"C0C0C0A499F8B092",
 24736 => x"C0C0C0A499F8B082",
 24737 => x"C0C0C0A499F8B0F8",
 24738 => x"C0C0C0A499F8B080",
 24739 => x"C0C0C0A499F8B090",
 24740 => x"C0C0C0A499F899C0",
 24741 => x"C0C0C0A499F899F9",
 24742 => x"C0C0C0A499F899A4",
 24743 => x"C0C0C0A499F899B0",
 24744 => x"C0C0C0A499F89999",
 24745 => x"C0C0C0A499F89992",
 24746 => x"C0C0C0A499F89982",
 24747 => x"C0C0C0A499F899F8",
 24748 => x"C0C0C0A499F89980",
 24749 => x"C0C0C0A499F89990",
 24750 => x"C0C0C0A499F892C0",
 24751 => x"C0C0C0A499F892F9",
 24752 => x"C0C0C0A499F892A4",
 24753 => x"C0C0C0A499F892B0",
 24754 => x"C0C0C0A499F89299",
 24755 => x"C0C0C0A499F89292",
 24756 => x"C0C0C0A499F89282",
 24757 => x"C0C0C0A499F892F8",
 24758 => x"C0C0C0A499F89280",
 24759 => x"C0C0C0A499F89290",
 24760 => x"C0C0C0A499F882C0",
 24761 => x"C0C0C0A499F882F9",
 24762 => x"C0C0C0A499F882A4",
 24763 => x"C0C0C0A499F882B0",
 24764 => x"C0C0C0A499F88299",
 24765 => x"C0C0C0A499F88292",
 24766 => x"C0C0C0A499F88282",
 24767 => x"C0C0C0A499F882F8",
 24768 => x"C0C0C0A499F88280",
 24769 => x"C0C0C0A499F88290",
 24770 => x"C0C0C0A499F8F8C0",
 24771 => x"C0C0C0A499F8F8F9",
 24772 => x"C0C0C0A499F8F8A4",
 24773 => x"C0C0C0A499F8F8B0",
 24774 => x"C0C0C0A499F8F899",
 24775 => x"C0C0C0A499F8F892",
 24776 => x"C0C0C0A499F8F882",
 24777 => x"C0C0C0A499F8F8F8",
 24778 => x"C0C0C0A499F8F880",
 24779 => x"C0C0C0A499F8F890",
 24780 => x"C0C0C0A499F880C0",
 24781 => x"C0C0C0A499F880F9",
 24782 => x"C0C0C0A499F880A4",
 24783 => x"C0C0C0A499F880B0",
 24784 => x"C0C0C0A499F88099",
 24785 => x"C0C0C0A499F88092",
 24786 => x"C0C0C0A499F88082",
 24787 => x"C0C0C0A499F880F8",
 24788 => x"C0C0C0A499F88080",
 24789 => x"C0C0C0A499F88090",
 24790 => x"C0C0C0A499F890C0",
 24791 => x"C0C0C0A499F890F9",
 24792 => x"C0C0C0A499F890A4",
 24793 => x"C0C0C0A499F890B0",
 24794 => x"C0C0C0A499F89099",
 24795 => x"C0C0C0A499F89092",
 24796 => x"C0C0C0A499F89082",
 24797 => x"C0C0C0A499F890F8",
 24798 => x"C0C0C0A499F89080",
 24799 => x"C0C0C0A499F89090",
 24800 => x"C0C0C0A49980C0C0",
 24801 => x"C0C0C0A49980C0F9",
 24802 => x"C0C0C0A49980C0A4",
 24803 => x"C0C0C0A49980C0B0",
 24804 => x"C0C0C0A49980C099",
 24805 => x"C0C0C0A49980C092",
 24806 => x"C0C0C0A49980C082",
 24807 => x"C0C0C0A49980C0F8",
 24808 => x"C0C0C0A49980C080",
 24809 => x"C0C0C0A49980C090",
 24810 => x"C0C0C0A49980F9C0",
 24811 => x"C0C0C0A49980F9F9",
 24812 => x"C0C0C0A49980F9A4",
 24813 => x"C0C0C0A49980F9B0",
 24814 => x"C0C0C0A49980F999",
 24815 => x"C0C0C0A49980F992",
 24816 => x"C0C0C0A49980F982",
 24817 => x"C0C0C0A49980F9F8",
 24818 => x"C0C0C0A49980F980",
 24819 => x"C0C0C0A49980F990",
 24820 => x"C0C0C0A49980A4C0",
 24821 => x"C0C0C0A49980A4F9",
 24822 => x"C0C0C0A49980A4A4",
 24823 => x"C0C0C0A49980A4B0",
 24824 => x"C0C0C0A49980A499",
 24825 => x"C0C0C0A49980A492",
 24826 => x"C0C0C0A49980A482",
 24827 => x"C0C0C0A49980A4F8",
 24828 => x"C0C0C0A49980A480",
 24829 => x"C0C0C0A49980A490",
 24830 => x"C0C0C0A49980B0C0",
 24831 => x"C0C0C0A49980B0F9",
 24832 => x"C0C0C0A49980B0A4",
 24833 => x"C0C0C0A49980B0B0",
 24834 => x"C0C0C0A49980B099",
 24835 => x"C0C0C0A49980B092",
 24836 => x"C0C0C0A49980B082",
 24837 => x"C0C0C0A49980B0F8",
 24838 => x"C0C0C0A49980B080",
 24839 => x"C0C0C0A49980B090",
 24840 => x"C0C0C0A4998099C0",
 24841 => x"C0C0C0A4998099F9",
 24842 => x"C0C0C0A4998099A4",
 24843 => x"C0C0C0A4998099B0",
 24844 => x"C0C0C0A499809999",
 24845 => x"C0C0C0A499809992",
 24846 => x"C0C0C0A499809982",
 24847 => x"C0C0C0A4998099F8",
 24848 => x"C0C0C0A499809980",
 24849 => x"C0C0C0A499809990",
 24850 => x"C0C0C0A4998092C0",
 24851 => x"C0C0C0A4998092F9",
 24852 => x"C0C0C0A4998092A4",
 24853 => x"C0C0C0A4998092B0",
 24854 => x"C0C0C0A499809299",
 24855 => x"C0C0C0A499809292",
 24856 => x"C0C0C0A499809282",
 24857 => x"C0C0C0A4998092F8",
 24858 => x"C0C0C0A499809280",
 24859 => x"C0C0C0A499809290",
 24860 => x"C0C0C0A4998082C0",
 24861 => x"C0C0C0A4998082F9",
 24862 => x"C0C0C0A4998082A4",
 24863 => x"C0C0C0A4998082B0",
 24864 => x"C0C0C0A499808299",
 24865 => x"C0C0C0A499808292",
 24866 => x"C0C0C0A499808282",
 24867 => x"C0C0C0A4998082F8",
 24868 => x"C0C0C0A499808280",
 24869 => x"C0C0C0A499808290",
 24870 => x"C0C0C0A49980F8C0",
 24871 => x"C0C0C0A49980F8F9",
 24872 => x"C0C0C0A49980F8A4",
 24873 => x"C0C0C0A49980F8B0",
 24874 => x"C0C0C0A49980F899",
 24875 => x"C0C0C0A49980F892",
 24876 => x"C0C0C0A49980F882",
 24877 => x"C0C0C0A49980F8F8",
 24878 => x"C0C0C0A49980F880",
 24879 => x"C0C0C0A49980F890",
 24880 => x"C0C0C0A4998080C0",
 24881 => x"C0C0C0A4998080F9",
 24882 => x"C0C0C0A4998080A4",
 24883 => x"C0C0C0A4998080B0",
 24884 => x"C0C0C0A499808099",
 24885 => x"C0C0C0A499808092",
 24886 => x"C0C0C0A499808082",
 24887 => x"C0C0C0A4998080F8",
 24888 => x"C0C0C0A499808080",
 24889 => x"C0C0C0A499808090",
 24890 => x"C0C0C0A4998090C0",
 24891 => x"C0C0C0A4998090F9",
 24892 => x"C0C0C0A4998090A4",
 24893 => x"C0C0C0A4998090B0",
 24894 => x"C0C0C0A499809099",
 24895 => x"C0C0C0A499809092",
 24896 => x"C0C0C0A499809082",
 24897 => x"C0C0C0A4998090F8",
 24898 => x"C0C0C0A499809080",
 24899 => x"C0C0C0A499809090",
 24900 => x"C0C0C0A49990C0C0",
 24901 => x"C0C0C0A49990C0F9",
 24902 => x"C0C0C0A49990C0A4",
 24903 => x"C0C0C0A49990C0B0",
 24904 => x"C0C0C0A49990C099",
 24905 => x"C0C0C0A49990C092",
 24906 => x"C0C0C0A49990C082",
 24907 => x"C0C0C0A49990C0F8",
 24908 => x"C0C0C0A49990C080",
 24909 => x"C0C0C0A49990C090",
 24910 => x"C0C0C0A49990F9C0",
 24911 => x"C0C0C0A49990F9F9",
 24912 => x"C0C0C0A49990F9A4",
 24913 => x"C0C0C0A49990F9B0",
 24914 => x"C0C0C0A49990F999",
 24915 => x"C0C0C0A49990F992",
 24916 => x"C0C0C0A49990F982",
 24917 => x"C0C0C0A49990F9F8",
 24918 => x"C0C0C0A49990F980",
 24919 => x"C0C0C0A49990F990",
 24920 => x"C0C0C0A49990A4C0",
 24921 => x"C0C0C0A49990A4F9",
 24922 => x"C0C0C0A49990A4A4",
 24923 => x"C0C0C0A49990A4B0",
 24924 => x"C0C0C0A49990A499",
 24925 => x"C0C0C0A49990A492",
 24926 => x"C0C0C0A49990A482",
 24927 => x"C0C0C0A49990A4F8",
 24928 => x"C0C0C0A49990A480",
 24929 => x"C0C0C0A49990A490",
 24930 => x"C0C0C0A49990B0C0",
 24931 => x"C0C0C0A49990B0F9",
 24932 => x"C0C0C0A49990B0A4",
 24933 => x"C0C0C0A49990B0B0",
 24934 => x"C0C0C0A49990B099",
 24935 => x"C0C0C0A49990B092",
 24936 => x"C0C0C0A49990B082",
 24937 => x"C0C0C0A49990B0F8",
 24938 => x"C0C0C0A49990B080",
 24939 => x"C0C0C0A49990B090",
 24940 => x"C0C0C0A4999099C0",
 24941 => x"C0C0C0A4999099F9",
 24942 => x"C0C0C0A4999099A4",
 24943 => x"C0C0C0A4999099B0",
 24944 => x"C0C0C0A499909999",
 24945 => x"C0C0C0A499909992",
 24946 => x"C0C0C0A499909982",
 24947 => x"C0C0C0A4999099F8",
 24948 => x"C0C0C0A499909980",
 24949 => x"C0C0C0A499909990",
 24950 => x"C0C0C0A4999092C0",
 24951 => x"C0C0C0A4999092F9",
 24952 => x"C0C0C0A4999092A4",
 24953 => x"C0C0C0A4999092B0",
 24954 => x"C0C0C0A499909299",
 24955 => x"C0C0C0A499909292",
 24956 => x"C0C0C0A499909282",
 24957 => x"C0C0C0A4999092F8",
 24958 => x"C0C0C0A499909280",
 24959 => x"C0C0C0A499909290",
 24960 => x"C0C0C0A4999082C0",
 24961 => x"C0C0C0A4999082F9",
 24962 => x"C0C0C0A4999082A4",
 24963 => x"C0C0C0A4999082B0",
 24964 => x"C0C0C0A499908299",
 24965 => x"C0C0C0A499908292",
 24966 => x"C0C0C0A499908282",
 24967 => x"C0C0C0A4999082F8",
 24968 => x"C0C0C0A499908280",
 24969 => x"C0C0C0A499908290",
 24970 => x"C0C0C0A49990F8C0",
 24971 => x"C0C0C0A49990F8F9",
 24972 => x"C0C0C0A49990F8A4",
 24973 => x"C0C0C0A49990F8B0",
 24974 => x"C0C0C0A49990F899",
 24975 => x"C0C0C0A49990F892",
 24976 => x"C0C0C0A49990F882",
 24977 => x"C0C0C0A49990F8F8",
 24978 => x"C0C0C0A49990F880",
 24979 => x"C0C0C0A49990F890",
 24980 => x"C0C0C0A4999080C0",
 24981 => x"C0C0C0A4999080F9",
 24982 => x"C0C0C0A4999080A4",
 24983 => x"C0C0C0A4999080B0",
 24984 => x"C0C0C0A499908099",
 24985 => x"C0C0C0A499908092",
 24986 => x"C0C0C0A499908082",
 24987 => x"C0C0C0A4999080F8",
 24988 => x"C0C0C0A499908080",
 24989 => x"C0C0C0A499908090",
 24990 => x"C0C0C0A4999090C0",
 24991 => x"C0C0C0A4999090F9",
 24992 => x"C0C0C0A4999090A4",
 24993 => x"C0C0C0A4999090B0",
 24994 => x"C0C0C0A499909099",
 24995 => x"C0C0C0A499909092",
 24996 => x"C0C0C0A499909082",
 24997 => x"C0C0C0A4999090F8",
 24998 => x"C0C0C0A499909080",
 24999 => x"C0C0C0A499909090",
 25000 => x"C0C0C0A492C0C0C0",
 25001 => x"C0C0C0A492C0C0F9",
 25002 => x"C0C0C0A492C0C0A4",
 25003 => x"C0C0C0A492C0C0B0",
 25004 => x"C0C0C0A492C0C099",
 25005 => x"C0C0C0A492C0C092",
 25006 => x"C0C0C0A492C0C082",
 25007 => x"C0C0C0A492C0C0F8",
 25008 => x"C0C0C0A492C0C080",
 25009 => x"C0C0C0A492C0C090",
 25010 => x"C0C0C0A492C0F9C0",
 25011 => x"C0C0C0A492C0F9F9",
 25012 => x"C0C0C0A492C0F9A4",
 25013 => x"C0C0C0A492C0F9B0",
 25014 => x"C0C0C0A492C0F999",
 25015 => x"C0C0C0A492C0F992",
 25016 => x"C0C0C0A492C0F982",
 25017 => x"C0C0C0A492C0F9F8",
 25018 => x"C0C0C0A492C0F980",
 25019 => x"C0C0C0A492C0F990",
 25020 => x"C0C0C0A492C0A4C0",
 25021 => x"C0C0C0A492C0A4F9",
 25022 => x"C0C0C0A492C0A4A4",
 25023 => x"C0C0C0A492C0A4B0",
 25024 => x"C0C0C0A492C0A499",
 25025 => x"C0C0C0A492C0A492",
 25026 => x"C0C0C0A492C0A482",
 25027 => x"C0C0C0A492C0A4F8",
 25028 => x"C0C0C0A492C0A480",
 25029 => x"C0C0C0A492C0A490",
 25030 => x"C0C0C0A492C0B0C0",
 25031 => x"C0C0C0A492C0B0F9",
 25032 => x"C0C0C0A492C0B0A4",
 25033 => x"C0C0C0A492C0B0B0",
 25034 => x"C0C0C0A492C0B099",
 25035 => x"C0C0C0A492C0B092",
 25036 => x"C0C0C0A492C0B082",
 25037 => x"C0C0C0A492C0B0F8",
 25038 => x"C0C0C0A492C0B080",
 25039 => x"C0C0C0A492C0B090",
 25040 => x"C0C0C0A492C099C0",
 25041 => x"C0C0C0A492C099F9",
 25042 => x"C0C0C0A492C099A4",
 25043 => x"C0C0C0A492C099B0",
 25044 => x"C0C0C0A492C09999",
 25045 => x"C0C0C0A492C09992",
 25046 => x"C0C0C0A492C09982",
 25047 => x"C0C0C0A492C099F8",
 25048 => x"C0C0C0A492C09980",
 25049 => x"C0C0C0A492C09990",
 25050 => x"C0C0C0A492C092C0",
 25051 => x"C0C0C0A492C092F9",
 25052 => x"C0C0C0A492C092A4",
 25053 => x"C0C0C0A492C092B0",
 25054 => x"C0C0C0A492C09299",
 25055 => x"C0C0C0A492C09292",
 25056 => x"C0C0C0A492C09282",
 25057 => x"C0C0C0A492C092F8",
 25058 => x"C0C0C0A492C09280",
 25059 => x"C0C0C0A492C09290",
 25060 => x"C0C0C0A492C082C0",
 25061 => x"C0C0C0A492C082F9",
 25062 => x"C0C0C0A492C082A4",
 25063 => x"C0C0C0A492C082B0",
 25064 => x"C0C0C0A492C08299",
 25065 => x"C0C0C0A492C08292",
 25066 => x"C0C0C0A492C08282",
 25067 => x"C0C0C0A492C082F8",
 25068 => x"C0C0C0A492C08280",
 25069 => x"C0C0C0A492C08290",
 25070 => x"C0C0C0A492C0F8C0",
 25071 => x"C0C0C0A492C0F8F9",
 25072 => x"C0C0C0A492C0F8A4",
 25073 => x"C0C0C0A492C0F8B0",
 25074 => x"C0C0C0A492C0F899",
 25075 => x"C0C0C0A492C0F892",
 25076 => x"C0C0C0A492C0F882",
 25077 => x"C0C0C0A492C0F8F8",
 25078 => x"C0C0C0A492C0F880",
 25079 => x"C0C0C0A492C0F890",
 25080 => x"C0C0C0A492C080C0",
 25081 => x"C0C0C0A492C080F9",
 25082 => x"C0C0C0A492C080A4",
 25083 => x"C0C0C0A492C080B0",
 25084 => x"C0C0C0A492C08099",
 25085 => x"C0C0C0A492C08092",
 25086 => x"C0C0C0A492C08082",
 25087 => x"C0C0C0A492C080F8",
 25088 => x"C0C0C0A492C08080",
 25089 => x"C0C0C0A492C08090",
 25090 => x"C0C0C0A492C090C0",
 25091 => x"C0C0C0A492C090F9",
 25092 => x"C0C0C0A492C090A4",
 25093 => x"C0C0C0A492C090B0",
 25094 => x"C0C0C0A492C09099",
 25095 => x"C0C0C0A492C09092",
 25096 => x"C0C0C0A492C09082",
 25097 => x"C0C0C0A492C090F8",
 25098 => x"C0C0C0A492C09080",
 25099 => x"C0C0C0A492C09090",
 25100 => x"C0C0C0A492F9C0C0",
 25101 => x"C0C0C0A492F9C0F9",
 25102 => x"C0C0C0A492F9C0A4",
 25103 => x"C0C0C0A492F9C0B0",
 25104 => x"C0C0C0A492F9C099",
 25105 => x"C0C0C0A492F9C092",
 25106 => x"C0C0C0A492F9C082",
 25107 => x"C0C0C0A492F9C0F8",
 25108 => x"C0C0C0A492F9C080",
 25109 => x"C0C0C0A492F9C090",
 25110 => x"C0C0C0A492F9F9C0",
 25111 => x"C0C0C0A492F9F9F9",
 25112 => x"C0C0C0A492F9F9A4",
 25113 => x"C0C0C0A492F9F9B0",
 25114 => x"C0C0C0A492F9F999",
 25115 => x"C0C0C0A492F9F992",
 25116 => x"C0C0C0A492F9F982",
 25117 => x"C0C0C0A492F9F9F8",
 25118 => x"C0C0C0A492F9F980",
 25119 => x"C0C0C0A492F9F990",
 25120 => x"C0C0C0A492F9A4C0",
 25121 => x"C0C0C0A492F9A4F9",
 25122 => x"C0C0C0A492F9A4A4",
 25123 => x"C0C0C0A492F9A4B0",
 25124 => x"C0C0C0A492F9A499",
 25125 => x"C0C0C0A492F9A492",
 25126 => x"C0C0C0A492F9A482",
 25127 => x"C0C0C0A492F9A4F8",
 25128 => x"C0C0C0A492F9A480",
 25129 => x"C0C0C0A492F9A490",
 25130 => x"C0C0C0A492F9B0C0",
 25131 => x"C0C0C0A492F9B0F9",
 25132 => x"C0C0C0A492F9B0A4",
 25133 => x"C0C0C0A492F9B0B0",
 25134 => x"C0C0C0A492F9B099",
 25135 => x"C0C0C0A492F9B092",
 25136 => x"C0C0C0A492F9B082",
 25137 => x"C0C0C0A492F9B0F8",
 25138 => x"C0C0C0A492F9B080",
 25139 => x"C0C0C0A492F9B090",
 25140 => x"C0C0C0A492F999C0",
 25141 => x"C0C0C0A492F999F9",
 25142 => x"C0C0C0A492F999A4",
 25143 => x"C0C0C0A492F999B0",
 25144 => x"C0C0C0A492F99999",
 25145 => x"C0C0C0A492F99992",
 25146 => x"C0C0C0A492F99982",
 25147 => x"C0C0C0A492F999F8",
 25148 => x"C0C0C0A492F99980",
 25149 => x"C0C0C0A492F99990",
 25150 => x"C0C0C0A492F992C0",
 25151 => x"C0C0C0A492F992F9",
 25152 => x"C0C0C0A492F992A4",
 25153 => x"C0C0C0A492F992B0",
 25154 => x"C0C0C0A492F99299",
 25155 => x"C0C0C0A492F99292",
 25156 => x"C0C0C0A492F99282",
 25157 => x"C0C0C0A492F992F8",
 25158 => x"C0C0C0A492F99280",
 25159 => x"C0C0C0A492F99290",
 25160 => x"C0C0C0A492F982C0",
 25161 => x"C0C0C0A492F982F9",
 25162 => x"C0C0C0A492F982A4",
 25163 => x"C0C0C0A492F982B0",
 25164 => x"C0C0C0A492F98299",
 25165 => x"C0C0C0A492F98292",
 25166 => x"C0C0C0A492F98282",
 25167 => x"C0C0C0A492F982F8",
 25168 => x"C0C0C0A492F98280",
 25169 => x"C0C0C0A492F98290",
 25170 => x"C0C0C0A492F9F8C0",
 25171 => x"C0C0C0A492F9F8F9",
 25172 => x"C0C0C0A492F9F8A4",
 25173 => x"C0C0C0A492F9F8B0",
 25174 => x"C0C0C0A492F9F899",
 25175 => x"C0C0C0A492F9F892",
 25176 => x"C0C0C0A492F9F882",
 25177 => x"C0C0C0A492F9F8F8",
 25178 => x"C0C0C0A492F9F880",
 25179 => x"C0C0C0A492F9F890",
 25180 => x"C0C0C0A492F980C0",
 25181 => x"C0C0C0A492F980F9",
 25182 => x"C0C0C0A492F980A4",
 25183 => x"C0C0C0A492F980B0",
 25184 => x"C0C0C0A492F98099",
 25185 => x"C0C0C0A492F98092",
 25186 => x"C0C0C0A492F98082",
 25187 => x"C0C0C0A492F980F8",
 25188 => x"C0C0C0A492F98080",
 25189 => x"C0C0C0A492F98090",
 25190 => x"C0C0C0A492F990C0",
 25191 => x"C0C0C0A492F990F9",
 25192 => x"C0C0C0A492F990A4",
 25193 => x"C0C0C0A492F990B0",
 25194 => x"C0C0C0A492F99099",
 25195 => x"C0C0C0A492F99092",
 25196 => x"C0C0C0A492F99082",
 25197 => x"C0C0C0A492F990F8",
 25198 => x"C0C0C0A492F99080",
 25199 => x"C0C0C0A492F99090",
 25200 => x"C0C0C0A492A4C0C0",
 25201 => x"C0C0C0A492A4C0F9",
 25202 => x"C0C0C0A492A4C0A4",
 25203 => x"C0C0C0A492A4C0B0",
 25204 => x"C0C0C0A492A4C099",
 25205 => x"C0C0C0A492A4C092",
 25206 => x"C0C0C0A492A4C082",
 25207 => x"C0C0C0A492A4C0F8",
 25208 => x"C0C0C0A492A4C080",
 25209 => x"C0C0C0A492A4C090",
 25210 => x"C0C0C0A492A4F9C0",
 25211 => x"C0C0C0A492A4F9F9",
 25212 => x"C0C0C0A492A4F9A4",
 25213 => x"C0C0C0A492A4F9B0",
 25214 => x"C0C0C0A492A4F999",
 25215 => x"C0C0C0A492A4F992",
 25216 => x"C0C0C0A492A4F982",
 25217 => x"C0C0C0A492A4F9F8",
 25218 => x"C0C0C0A492A4F980",
 25219 => x"C0C0C0A492A4F990",
 25220 => x"C0C0C0A492A4A4C0",
 25221 => x"C0C0C0A492A4A4F9",
 25222 => x"C0C0C0A492A4A4A4",
 25223 => x"C0C0C0A492A4A4B0",
 25224 => x"C0C0C0A492A4A499",
 25225 => x"C0C0C0A492A4A492",
 25226 => x"C0C0C0A492A4A482",
 25227 => x"C0C0C0A492A4A4F8",
 25228 => x"C0C0C0A492A4A480",
 25229 => x"C0C0C0A492A4A490",
 25230 => x"C0C0C0A492A4B0C0",
 25231 => x"C0C0C0A492A4B0F9",
 25232 => x"C0C0C0A492A4B0A4",
 25233 => x"C0C0C0A492A4B0B0",
 25234 => x"C0C0C0A492A4B099",
 25235 => x"C0C0C0A492A4B092",
 25236 => x"C0C0C0A492A4B082",
 25237 => x"C0C0C0A492A4B0F8",
 25238 => x"C0C0C0A492A4B080",
 25239 => x"C0C0C0A492A4B090",
 25240 => x"C0C0C0A492A499C0",
 25241 => x"C0C0C0A492A499F9",
 25242 => x"C0C0C0A492A499A4",
 25243 => x"C0C0C0A492A499B0",
 25244 => x"C0C0C0A492A49999",
 25245 => x"C0C0C0A492A49992",
 25246 => x"C0C0C0A492A49982",
 25247 => x"C0C0C0A492A499F8",
 25248 => x"C0C0C0A492A49980",
 25249 => x"C0C0C0A492A49990",
 25250 => x"C0C0C0A492A492C0",
 25251 => x"C0C0C0A492A492F9",
 25252 => x"C0C0C0A492A492A4",
 25253 => x"C0C0C0A492A492B0",
 25254 => x"C0C0C0A492A49299",
 25255 => x"C0C0C0A492A49292",
 25256 => x"C0C0C0A492A49282",
 25257 => x"C0C0C0A492A492F8",
 25258 => x"C0C0C0A492A49280",
 25259 => x"C0C0C0A492A49290",
 25260 => x"C0C0C0A492A482C0",
 25261 => x"C0C0C0A492A482F9",
 25262 => x"C0C0C0A492A482A4",
 25263 => x"C0C0C0A492A482B0",
 25264 => x"C0C0C0A492A48299",
 25265 => x"C0C0C0A492A48292",
 25266 => x"C0C0C0A492A48282",
 25267 => x"C0C0C0A492A482F8",
 25268 => x"C0C0C0A492A48280",
 25269 => x"C0C0C0A492A48290",
 25270 => x"C0C0C0A492A4F8C0",
 25271 => x"C0C0C0A492A4F8F9",
 25272 => x"C0C0C0A492A4F8A4",
 25273 => x"C0C0C0A492A4F8B0",
 25274 => x"C0C0C0A492A4F899",
 25275 => x"C0C0C0A492A4F892",
 25276 => x"C0C0C0A492A4F882",
 25277 => x"C0C0C0A492A4F8F8",
 25278 => x"C0C0C0A492A4F880",
 25279 => x"C0C0C0A492A4F890",
 25280 => x"C0C0C0A492A480C0",
 25281 => x"C0C0C0A492A480F9",
 25282 => x"C0C0C0A492A480A4",
 25283 => x"C0C0C0A492A480B0",
 25284 => x"C0C0C0A492A48099",
 25285 => x"C0C0C0A492A48092",
 25286 => x"C0C0C0A492A48082",
 25287 => x"C0C0C0A492A480F8",
 25288 => x"C0C0C0A492A48080",
 25289 => x"C0C0C0A492A48090",
 25290 => x"C0C0C0A492A490C0",
 25291 => x"C0C0C0A492A490F9",
 25292 => x"C0C0C0A492A490A4",
 25293 => x"C0C0C0A492A490B0",
 25294 => x"C0C0C0A492A49099",
 25295 => x"C0C0C0A492A49092",
 25296 => x"C0C0C0A492A49082",
 25297 => x"C0C0C0A492A490F8",
 25298 => x"C0C0C0A492A49080",
 25299 => x"C0C0C0A492A49090",
 25300 => x"C0C0C0A492B0C0C0",
 25301 => x"C0C0C0A492B0C0F9",
 25302 => x"C0C0C0A492B0C0A4",
 25303 => x"C0C0C0A492B0C0B0",
 25304 => x"C0C0C0A492B0C099",
 25305 => x"C0C0C0A492B0C092",
 25306 => x"C0C0C0A492B0C082",
 25307 => x"C0C0C0A492B0C0F8",
 25308 => x"C0C0C0A492B0C080",
 25309 => x"C0C0C0A492B0C090",
 25310 => x"C0C0C0A492B0F9C0",
 25311 => x"C0C0C0A492B0F9F9",
 25312 => x"C0C0C0A492B0F9A4",
 25313 => x"C0C0C0A492B0F9B0",
 25314 => x"C0C0C0A492B0F999",
 25315 => x"C0C0C0A492B0F992",
 25316 => x"C0C0C0A492B0F982",
 25317 => x"C0C0C0A492B0F9F8",
 25318 => x"C0C0C0A492B0F980",
 25319 => x"C0C0C0A492B0F990",
 25320 => x"C0C0C0A492B0A4C0",
 25321 => x"C0C0C0A492B0A4F9",
 25322 => x"C0C0C0A492B0A4A4",
 25323 => x"C0C0C0A492B0A4B0",
 25324 => x"C0C0C0A492B0A499",
 25325 => x"C0C0C0A492B0A492",
 25326 => x"C0C0C0A492B0A482",
 25327 => x"C0C0C0A492B0A4F8",
 25328 => x"C0C0C0A492B0A480",
 25329 => x"C0C0C0A492B0A490",
 25330 => x"C0C0C0A492B0B0C0",
 25331 => x"C0C0C0A492B0B0F9",
 25332 => x"C0C0C0A492B0B0A4",
 25333 => x"C0C0C0A492B0B0B0",
 25334 => x"C0C0C0A492B0B099",
 25335 => x"C0C0C0A492B0B092",
 25336 => x"C0C0C0A492B0B082",
 25337 => x"C0C0C0A492B0B0F8",
 25338 => x"C0C0C0A492B0B080",
 25339 => x"C0C0C0A492B0B090",
 25340 => x"C0C0C0A492B099C0",
 25341 => x"C0C0C0A492B099F9",
 25342 => x"C0C0C0A492B099A4",
 25343 => x"C0C0C0A492B099B0",
 25344 => x"C0C0C0A492B09999",
 25345 => x"C0C0C0A492B09992",
 25346 => x"C0C0C0A492B09982",
 25347 => x"C0C0C0A492B099F8",
 25348 => x"C0C0C0A492B09980",
 25349 => x"C0C0C0A492B09990",
 25350 => x"C0C0C0A492B092C0",
 25351 => x"C0C0C0A492B092F9",
 25352 => x"C0C0C0A492B092A4",
 25353 => x"C0C0C0A492B092B0",
 25354 => x"C0C0C0A492B09299",
 25355 => x"C0C0C0A492B09292",
 25356 => x"C0C0C0A492B09282",
 25357 => x"C0C0C0A492B092F8",
 25358 => x"C0C0C0A492B09280",
 25359 => x"C0C0C0A492B09290",
 25360 => x"C0C0C0A492B082C0",
 25361 => x"C0C0C0A492B082F9",
 25362 => x"C0C0C0A492B082A4",
 25363 => x"C0C0C0A492B082B0",
 25364 => x"C0C0C0A492B08299",
 25365 => x"C0C0C0A492B08292",
 25366 => x"C0C0C0A492B08282",
 25367 => x"C0C0C0A492B082F8",
 25368 => x"C0C0C0A492B08280",
 25369 => x"C0C0C0A492B08290",
 25370 => x"C0C0C0A492B0F8C0",
 25371 => x"C0C0C0A492B0F8F9",
 25372 => x"C0C0C0A492B0F8A4",
 25373 => x"C0C0C0A492B0F8B0",
 25374 => x"C0C0C0A492B0F899",
 25375 => x"C0C0C0A492B0F892",
 25376 => x"C0C0C0A492B0F882",
 25377 => x"C0C0C0A492B0F8F8",
 25378 => x"C0C0C0A492B0F880",
 25379 => x"C0C0C0A492B0F890",
 25380 => x"C0C0C0A492B080C0",
 25381 => x"C0C0C0A492B080F9",
 25382 => x"C0C0C0A492B080A4",
 25383 => x"C0C0C0A492B080B0",
 25384 => x"C0C0C0A492B08099",
 25385 => x"C0C0C0A492B08092",
 25386 => x"C0C0C0A492B08082",
 25387 => x"C0C0C0A492B080F8",
 25388 => x"C0C0C0A492B08080",
 25389 => x"C0C0C0A492B08090",
 25390 => x"C0C0C0A492B090C0",
 25391 => x"C0C0C0A492B090F9",
 25392 => x"C0C0C0A492B090A4",
 25393 => x"C0C0C0A492B090B0",
 25394 => x"C0C0C0A492B09099",
 25395 => x"C0C0C0A492B09092",
 25396 => x"C0C0C0A492B09082",
 25397 => x"C0C0C0A492B090F8",
 25398 => x"C0C0C0A492B09080",
 25399 => x"C0C0C0A492B09090",
 25400 => x"C0C0C0A49299C0C0",
 25401 => x"C0C0C0A49299C0F9",
 25402 => x"C0C0C0A49299C0A4",
 25403 => x"C0C0C0A49299C0B0",
 25404 => x"C0C0C0A49299C099",
 25405 => x"C0C0C0A49299C092",
 25406 => x"C0C0C0A49299C082",
 25407 => x"C0C0C0A49299C0F8",
 25408 => x"C0C0C0A49299C080",
 25409 => x"C0C0C0A49299C090",
 25410 => x"C0C0C0A49299F9C0",
 25411 => x"C0C0C0A49299F9F9",
 25412 => x"C0C0C0A49299F9A4",
 25413 => x"C0C0C0A49299F9B0",
 25414 => x"C0C0C0A49299F999",
 25415 => x"C0C0C0A49299F992",
 25416 => x"C0C0C0A49299F982",
 25417 => x"C0C0C0A49299F9F8",
 25418 => x"C0C0C0A49299F980",
 25419 => x"C0C0C0A49299F990",
 25420 => x"C0C0C0A49299A4C0",
 25421 => x"C0C0C0A49299A4F9",
 25422 => x"C0C0C0A49299A4A4",
 25423 => x"C0C0C0A49299A4B0",
 25424 => x"C0C0C0A49299A499",
 25425 => x"C0C0C0A49299A492",
 25426 => x"C0C0C0A49299A482",
 25427 => x"C0C0C0A49299A4F8",
 25428 => x"C0C0C0A49299A480",
 25429 => x"C0C0C0A49299A490",
 25430 => x"C0C0C0A49299B0C0",
 25431 => x"C0C0C0A49299B0F9",
 25432 => x"C0C0C0A49299B0A4",
 25433 => x"C0C0C0A49299B0B0",
 25434 => x"C0C0C0A49299B099",
 25435 => x"C0C0C0A49299B092",
 25436 => x"C0C0C0A49299B082",
 25437 => x"C0C0C0A49299B0F8",
 25438 => x"C0C0C0A49299B080",
 25439 => x"C0C0C0A49299B090",
 25440 => x"C0C0C0A4929999C0",
 25441 => x"C0C0C0A4929999F9",
 25442 => x"C0C0C0A4929999A4",
 25443 => x"C0C0C0A4929999B0",
 25444 => x"C0C0C0A492999999",
 25445 => x"C0C0C0A492999992",
 25446 => x"C0C0C0A492999982",
 25447 => x"C0C0C0A4929999F8",
 25448 => x"C0C0C0A492999980",
 25449 => x"C0C0C0A492999990",
 25450 => x"C0C0C0A4929992C0",
 25451 => x"C0C0C0A4929992F9",
 25452 => x"C0C0C0A4929992A4",
 25453 => x"C0C0C0A4929992B0",
 25454 => x"C0C0C0A492999299",
 25455 => x"C0C0C0A492999292",
 25456 => x"C0C0C0A492999282",
 25457 => x"C0C0C0A4929992F8",
 25458 => x"C0C0C0A492999280",
 25459 => x"C0C0C0A492999290",
 25460 => x"C0C0C0A4929982C0",
 25461 => x"C0C0C0A4929982F9",
 25462 => x"C0C0C0A4929982A4",
 25463 => x"C0C0C0A4929982B0",
 25464 => x"C0C0C0A492998299",
 25465 => x"C0C0C0A492998292",
 25466 => x"C0C0C0A492998282",
 25467 => x"C0C0C0A4929982F8",
 25468 => x"C0C0C0A492998280",
 25469 => x"C0C0C0A492998290",
 25470 => x"C0C0C0A49299F8C0",
 25471 => x"C0C0C0A49299F8F9",
 25472 => x"C0C0C0A49299F8A4",
 25473 => x"C0C0C0A49299F8B0",
 25474 => x"C0C0C0A49299F899",
 25475 => x"C0C0C0A49299F892",
 25476 => x"C0C0C0A49299F882",
 25477 => x"C0C0C0A49299F8F8",
 25478 => x"C0C0C0A49299F880",
 25479 => x"C0C0C0A49299F890",
 25480 => x"C0C0C0A4929980C0",
 25481 => x"C0C0C0A4929980F9",
 25482 => x"C0C0C0A4929980A4",
 25483 => x"C0C0C0A4929980B0",
 25484 => x"C0C0C0A492998099",
 25485 => x"C0C0C0A492998092",
 25486 => x"C0C0C0A492998082",
 25487 => x"C0C0C0A4929980F8",
 25488 => x"C0C0C0A492998080",
 25489 => x"C0C0C0A492998090",
 25490 => x"C0C0C0A4929990C0",
 25491 => x"C0C0C0A4929990F9",
 25492 => x"C0C0C0A4929990A4",
 25493 => x"C0C0C0A4929990B0",
 25494 => x"C0C0C0A492999099",
 25495 => x"C0C0C0A492999092",
 25496 => x"C0C0C0A492999082",
 25497 => x"C0C0C0A4929990F8",
 25498 => x"C0C0C0A492999080",
 25499 => x"C0C0C0A492999090",
 25500 => x"C0C0C0A49292C0C0",
 25501 => x"C0C0C0A49292C0F9",
 25502 => x"C0C0C0A49292C0A4",
 25503 => x"C0C0C0A49292C0B0",
 25504 => x"C0C0C0A49292C099",
 25505 => x"C0C0C0A49292C092",
 25506 => x"C0C0C0A49292C082",
 25507 => x"C0C0C0A49292C0F8",
 25508 => x"C0C0C0A49292C080",
 25509 => x"C0C0C0A49292C090",
 25510 => x"C0C0C0A49292F9C0",
 25511 => x"C0C0C0A49292F9F9",
 25512 => x"C0C0C0A49292F9A4",
 25513 => x"C0C0C0A49292F9B0",
 25514 => x"C0C0C0A49292F999",
 25515 => x"C0C0C0A49292F992",
 25516 => x"C0C0C0A49292F982",
 25517 => x"C0C0C0A49292F9F8",
 25518 => x"C0C0C0A49292F980",
 25519 => x"C0C0C0A49292F990",
 25520 => x"C0C0C0A49292A4C0",
 25521 => x"C0C0C0A49292A4F9",
 25522 => x"C0C0C0A49292A4A4",
 25523 => x"C0C0C0A49292A4B0",
 25524 => x"C0C0C0A49292A499",
 25525 => x"C0C0C0A49292A492",
 25526 => x"C0C0C0A49292A482",
 25527 => x"C0C0C0A49292A4F8",
 25528 => x"C0C0C0A49292A480",
 25529 => x"C0C0C0A49292A490",
 25530 => x"C0C0C0A49292B0C0",
 25531 => x"C0C0C0A49292B0F9",
 25532 => x"C0C0C0A49292B0A4",
 25533 => x"C0C0C0A49292B0B0",
 25534 => x"C0C0C0A49292B099",
 25535 => x"C0C0C0A49292B092",
 25536 => x"C0C0C0A49292B082",
 25537 => x"C0C0C0A49292B0F8",
 25538 => x"C0C0C0A49292B080",
 25539 => x"C0C0C0A49292B090",
 25540 => x"C0C0C0A4929299C0",
 25541 => x"C0C0C0A4929299F9",
 25542 => x"C0C0C0A4929299A4",
 25543 => x"C0C0C0A4929299B0",
 25544 => x"C0C0C0A492929999",
 25545 => x"C0C0C0A492929992",
 25546 => x"C0C0C0A492929982",
 25547 => x"C0C0C0A4929299F8",
 25548 => x"C0C0C0A492929980",
 25549 => x"C0C0C0A492929990",
 25550 => x"C0C0C0A4929292C0",
 25551 => x"C0C0C0A4929292F9",
 25552 => x"C0C0C0A4929292A4",
 25553 => x"C0C0C0A4929292B0",
 25554 => x"C0C0C0A492929299",
 25555 => x"C0C0C0A492929292",
 25556 => x"C0C0C0A492929282",
 25557 => x"C0C0C0A4929292F8",
 25558 => x"C0C0C0A492929280",
 25559 => x"C0C0C0A492929290",
 25560 => x"C0C0C0A4929282C0",
 25561 => x"C0C0C0A4929282F9",
 25562 => x"C0C0C0A4929282A4",
 25563 => x"C0C0C0A4929282B0",
 25564 => x"C0C0C0A492928299",
 25565 => x"C0C0C0A492928292",
 25566 => x"C0C0C0A492928282",
 25567 => x"C0C0C0A4929282F8",
 25568 => x"C0C0C0A492928280",
 25569 => x"C0C0C0A492928290",
 25570 => x"C0C0C0A49292F8C0",
 25571 => x"C0C0C0A49292F8F9",
 25572 => x"C0C0C0A49292F8A4",
 25573 => x"C0C0C0A49292F8B0",
 25574 => x"C0C0C0A49292F899",
 25575 => x"C0C0C0A49292F892",
 25576 => x"C0C0C0A49292F882",
 25577 => x"C0C0C0A49292F8F8",
 25578 => x"C0C0C0A49292F880",
 25579 => x"C0C0C0A49292F890",
 25580 => x"C0C0C0A4929280C0",
 25581 => x"C0C0C0A4929280F9",
 25582 => x"C0C0C0A4929280A4",
 25583 => x"C0C0C0A4929280B0",
 25584 => x"C0C0C0A492928099",
 25585 => x"C0C0C0A492928092",
 25586 => x"C0C0C0A492928082",
 25587 => x"C0C0C0A4929280F8",
 25588 => x"C0C0C0A492928080",
 25589 => x"C0C0C0A492928090",
 25590 => x"C0C0C0A4929290C0",
 25591 => x"C0C0C0A4929290F9",
 25592 => x"C0C0C0A4929290A4",
 25593 => x"C0C0C0A4929290B0",
 25594 => x"C0C0C0A492929099",
 25595 => x"C0C0C0A492929092",
 25596 => x"C0C0C0A492929082",
 25597 => x"C0C0C0A4929290F8",
 25598 => x"C0C0C0A492929080",
 25599 => x"C0C0C0A492929090",
 25600 => x"C0C0C0A49282C0C0",
 25601 => x"C0C0C0A49282C0F9",
 25602 => x"C0C0C0A49282C0A4",
 25603 => x"C0C0C0A49282C0B0",
 25604 => x"C0C0C0A49282C099",
 25605 => x"C0C0C0A49282C092",
 25606 => x"C0C0C0A49282C082",
 25607 => x"C0C0C0A49282C0F8",
 25608 => x"C0C0C0A49282C080",
 25609 => x"C0C0C0A49282C090",
 25610 => x"C0C0C0A49282F9C0",
 25611 => x"C0C0C0A49282F9F9",
 25612 => x"C0C0C0A49282F9A4",
 25613 => x"C0C0C0A49282F9B0",
 25614 => x"C0C0C0A49282F999",
 25615 => x"C0C0C0A49282F992",
 25616 => x"C0C0C0A49282F982",
 25617 => x"C0C0C0A49282F9F8",
 25618 => x"C0C0C0A49282F980",
 25619 => x"C0C0C0A49282F990",
 25620 => x"C0C0C0A49282A4C0",
 25621 => x"C0C0C0A49282A4F9",
 25622 => x"C0C0C0A49282A4A4",
 25623 => x"C0C0C0A49282A4B0",
 25624 => x"C0C0C0A49282A499",
 25625 => x"C0C0C0A49282A492",
 25626 => x"C0C0C0A49282A482",
 25627 => x"C0C0C0A49282A4F8",
 25628 => x"C0C0C0A49282A480",
 25629 => x"C0C0C0A49282A490",
 25630 => x"C0C0C0A49282B0C0",
 25631 => x"C0C0C0A49282B0F9",
 25632 => x"C0C0C0A49282B0A4",
 25633 => x"C0C0C0A49282B0B0",
 25634 => x"C0C0C0A49282B099",
 25635 => x"C0C0C0A49282B092",
 25636 => x"C0C0C0A49282B082",
 25637 => x"C0C0C0A49282B0F8",
 25638 => x"C0C0C0A49282B080",
 25639 => x"C0C0C0A49282B090",
 25640 => x"C0C0C0A4928299C0",
 25641 => x"C0C0C0A4928299F9",
 25642 => x"C0C0C0A4928299A4",
 25643 => x"C0C0C0A4928299B0",
 25644 => x"C0C0C0A492829999",
 25645 => x"C0C0C0A492829992",
 25646 => x"C0C0C0A492829982",
 25647 => x"C0C0C0A4928299F8",
 25648 => x"C0C0C0A492829980",
 25649 => x"C0C0C0A492829990",
 25650 => x"C0C0C0A4928292C0",
 25651 => x"C0C0C0A4928292F9",
 25652 => x"C0C0C0A4928292A4",
 25653 => x"C0C0C0A4928292B0",
 25654 => x"C0C0C0A492829299",
 25655 => x"C0C0C0A492829292",
 25656 => x"C0C0C0A492829282",
 25657 => x"C0C0C0A4928292F8",
 25658 => x"C0C0C0A492829280",
 25659 => x"C0C0C0A492829290",
 25660 => x"C0C0C0A4928282C0",
 25661 => x"C0C0C0A4928282F9",
 25662 => x"C0C0C0A4928282A4",
 25663 => x"C0C0C0A4928282B0",
 25664 => x"C0C0C0A492828299",
 25665 => x"C0C0C0A492828292",
 25666 => x"C0C0C0A492828282",
 25667 => x"C0C0C0A4928282F8",
 25668 => x"C0C0C0A492828280",
 25669 => x"C0C0C0A492828290",
 25670 => x"C0C0C0A49282F8C0",
 25671 => x"C0C0C0A49282F8F9",
 25672 => x"C0C0C0A49282F8A4",
 25673 => x"C0C0C0A49282F8B0",
 25674 => x"C0C0C0A49282F899",
 25675 => x"C0C0C0A49282F892",
 25676 => x"C0C0C0A49282F882",
 25677 => x"C0C0C0A49282F8F8",
 25678 => x"C0C0C0A49282F880",
 25679 => x"C0C0C0A49282F890",
 25680 => x"C0C0C0A4928280C0",
 25681 => x"C0C0C0A4928280F9",
 25682 => x"C0C0C0A4928280A4",
 25683 => x"C0C0C0A4928280B0",
 25684 => x"C0C0C0A492828099",
 25685 => x"C0C0C0A492828092",
 25686 => x"C0C0C0A492828082",
 25687 => x"C0C0C0A4928280F8",
 25688 => x"C0C0C0A492828080",
 25689 => x"C0C0C0A492828090",
 25690 => x"C0C0C0A4928290C0",
 25691 => x"C0C0C0A4928290F9",
 25692 => x"C0C0C0A4928290A4",
 25693 => x"C0C0C0A4928290B0",
 25694 => x"C0C0C0A492829099",
 25695 => x"C0C0C0A492829092",
 25696 => x"C0C0C0A492829082",
 25697 => x"C0C0C0A4928290F8",
 25698 => x"C0C0C0A492829080",
 25699 => x"C0C0C0A492829090",
 25700 => x"C0C0C0A492F8C0C0",
 25701 => x"C0C0C0A492F8C0F9",
 25702 => x"C0C0C0A492F8C0A4",
 25703 => x"C0C0C0A492F8C0B0",
 25704 => x"C0C0C0A492F8C099",
 25705 => x"C0C0C0A492F8C092",
 25706 => x"C0C0C0A492F8C082",
 25707 => x"C0C0C0A492F8C0F8",
 25708 => x"C0C0C0A492F8C080",
 25709 => x"C0C0C0A492F8C090",
 25710 => x"C0C0C0A492F8F9C0",
 25711 => x"C0C0C0A492F8F9F9",
 25712 => x"C0C0C0A492F8F9A4",
 25713 => x"C0C0C0A492F8F9B0",
 25714 => x"C0C0C0A492F8F999",
 25715 => x"C0C0C0A492F8F992",
 25716 => x"C0C0C0A492F8F982",
 25717 => x"C0C0C0A492F8F9F8",
 25718 => x"C0C0C0A492F8F980",
 25719 => x"C0C0C0A492F8F990",
 25720 => x"C0C0C0A492F8A4C0",
 25721 => x"C0C0C0A492F8A4F9",
 25722 => x"C0C0C0A492F8A4A4",
 25723 => x"C0C0C0A492F8A4B0",
 25724 => x"C0C0C0A492F8A499",
 25725 => x"C0C0C0A492F8A492",
 25726 => x"C0C0C0A492F8A482",
 25727 => x"C0C0C0A492F8A4F8",
 25728 => x"C0C0C0A492F8A480",
 25729 => x"C0C0C0A492F8A490",
 25730 => x"C0C0C0A492F8B0C0",
 25731 => x"C0C0C0A492F8B0F9",
 25732 => x"C0C0C0A492F8B0A4",
 25733 => x"C0C0C0A492F8B0B0",
 25734 => x"C0C0C0A492F8B099",
 25735 => x"C0C0C0A492F8B092",
 25736 => x"C0C0C0A492F8B082",
 25737 => x"C0C0C0A492F8B0F8",
 25738 => x"C0C0C0A492F8B080",
 25739 => x"C0C0C0A492F8B090",
 25740 => x"C0C0C0A492F899C0",
 25741 => x"C0C0C0A492F899F9",
 25742 => x"C0C0C0A492F899A4",
 25743 => x"C0C0C0A492F899B0",
 25744 => x"C0C0C0A492F89999",
 25745 => x"C0C0C0A492F89992",
 25746 => x"C0C0C0A492F89982",
 25747 => x"C0C0C0A492F899F8",
 25748 => x"C0C0C0A492F89980",
 25749 => x"C0C0C0A492F89990",
 25750 => x"C0C0C0A492F892C0",
 25751 => x"C0C0C0A492F892F9",
 25752 => x"C0C0C0A492F892A4",
 25753 => x"C0C0C0A492F892B0",
 25754 => x"C0C0C0A492F89299",
 25755 => x"C0C0C0A492F89292",
 25756 => x"C0C0C0A492F89282",
 25757 => x"C0C0C0A492F892F8",
 25758 => x"C0C0C0A492F89280",
 25759 => x"C0C0C0A492F89290",
 25760 => x"C0C0C0A492F882C0",
 25761 => x"C0C0C0A492F882F9",
 25762 => x"C0C0C0A492F882A4",
 25763 => x"C0C0C0A492F882B0",
 25764 => x"C0C0C0A492F88299",
 25765 => x"C0C0C0A492F88292",
 25766 => x"C0C0C0A492F88282",
 25767 => x"C0C0C0A492F882F8",
 25768 => x"C0C0C0A492F88280",
 25769 => x"C0C0C0A492F88290",
 25770 => x"C0C0C0A492F8F8C0",
 25771 => x"C0C0C0A492F8F8F9",
 25772 => x"C0C0C0A492F8F8A4",
 25773 => x"C0C0C0A492F8F8B0",
 25774 => x"C0C0C0A492F8F899",
 25775 => x"C0C0C0A492F8F892",
 25776 => x"C0C0C0A492F8F882",
 25777 => x"C0C0C0A492F8F8F8",
 25778 => x"C0C0C0A492F8F880",
 25779 => x"C0C0C0A492F8F890",
 25780 => x"C0C0C0A492F880C0",
 25781 => x"C0C0C0A492F880F9",
 25782 => x"C0C0C0A492F880A4",
 25783 => x"C0C0C0A492F880B0",
 25784 => x"C0C0C0A492F88099",
 25785 => x"C0C0C0A492F88092",
 25786 => x"C0C0C0A492F88082",
 25787 => x"C0C0C0A492F880F8",
 25788 => x"C0C0C0A492F88080",
 25789 => x"C0C0C0A492F88090",
 25790 => x"C0C0C0A492F890C0",
 25791 => x"C0C0C0A492F890F9",
 25792 => x"C0C0C0A492F890A4",
 25793 => x"C0C0C0A492F890B0",
 25794 => x"C0C0C0A492F89099",
 25795 => x"C0C0C0A492F89092",
 25796 => x"C0C0C0A492F89082",
 25797 => x"C0C0C0A492F890F8",
 25798 => x"C0C0C0A492F89080",
 25799 => x"C0C0C0A492F89090",
 25800 => x"C0C0C0A49280C0C0",
 25801 => x"C0C0C0A49280C0F9",
 25802 => x"C0C0C0A49280C0A4",
 25803 => x"C0C0C0A49280C0B0",
 25804 => x"C0C0C0A49280C099",
 25805 => x"C0C0C0A49280C092",
 25806 => x"C0C0C0A49280C082",
 25807 => x"C0C0C0A49280C0F8",
 25808 => x"C0C0C0A49280C080",
 25809 => x"C0C0C0A49280C090",
 25810 => x"C0C0C0A49280F9C0",
 25811 => x"C0C0C0A49280F9F9",
 25812 => x"C0C0C0A49280F9A4",
 25813 => x"C0C0C0A49280F9B0",
 25814 => x"C0C0C0A49280F999",
 25815 => x"C0C0C0A49280F992",
 25816 => x"C0C0C0A49280F982",
 25817 => x"C0C0C0A49280F9F8",
 25818 => x"C0C0C0A49280F980",
 25819 => x"C0C0C0A49280F990",
 25820 => x"C0C0C0A49280A4C0",
 25821 => x"C0C0C0A49280A4F9",
 25822 => x"C0C0C0A49280A4A4",
 25823 => x"C0C0C0A49280A4B0",
 25824 => x"C0C0C0A49280A499",
 25825 => x"C0C0C0A49280A492",
 25826 => x"C0C0C0A49280A482",
 25827 => x"C0C0C0A49280A4F8",
 25828 => x"C0C0C0A49280A480",
 25829 => x"C0C0C0A49280A490",
 25830 => x"C0C0C0A49280B0C0",
 25831 => x"C0C0C0A49280B0F9",
 25832 => x"C0C0C0A49280B0A4",
 25833 => x"C0C0C0A49280B0B0",
 25834 => x"C0C0C0A49280B099",
 25835 => x"C0C0C0A49280B092",
 25836 => x"C0C0C0A49280B082",
 25837 => x"C0C0C0A49280B0F8",
 25838 => x"C0C0C0A49280B080",
 25839 => x"C0C0C0A49280B090",
 25840 => x"C0C0C0A4928099C0",
 25841 => x"C0C0C0A4928099F9",
 25842 => x"C0C0C0A4928099A4",
 25843 => x"C0C0C0A4928099B0",
 25844 => x"C0C0C0A492809999",
 25845 => x"C0C0C0A492809992",
 25846 => x"C0C0C0A492809982",
 25847 => x"C0C0C0A4928099F8",
 25848 => x"C0C0C0A492809980",
 25849 => x"C0C0C0A492809990",
 25850 => x"C0C0C0A4928092C0",
 25851 => x"C0C0C0A4928092F9",
 25852 => x"C0C0C0A4928092A4",
 25853 => x"C0C0C0A4928092B0",
 25854 => x"C0C0C0A492809299",
 25855 => x"C0C0C0A492809292",
 25856 => x"C0C0C0A492809282",
 25857 => x"C0C0C0A4928092F8",
 25858 => x"C0C0C0A492809280",
 25859 => x"C0C0C0A492809290",
 25860 => x"C0C0C0A4928082C0",
 25861 => x"C0C0C0A4928082F9",
 25862 => x"C0C0C0A4928082A4",
 25863 => x"C0C0C0A4928082B0",
 25864 => x"C0C0C0A492808299",
 25865 => x"C0C0C0A492808292",
 25866 => x"C0C0C0A492808282",
 25867 => x"C0C0C0A4928082F8",
 25868 => x"C0C0C0A492808280",
 25869 => x"C0C0C0A492808290",
 25870 => x"C0C0C0A49280F8C0",
 25871 => x"C0C0C0A49280F8F9",
 25872 => x"C0C0C0A49280F8A4",
 25873 => x"C0C0C0A49280F8B0",
 25874 => x"C0C0C0A49280F899",
 25875 => x"C0C0C0A49280F892",
 25876 => x"C0C0C0A49280F882",
 25877 => x"C0C0C0A49280F8F8",
 25878 => x"C0C0C0A49280F880",
 25879 => x"C0C0C0A49280F890",
 25880 => x"C0C0C0A4928080C0",
 25881 => x"C0C0C0A4928080F9",
 25882 => x"C0C0C0A4928080A4",
 25883 => x"C0C0C0A4928080B0",
 25884 => x"C0C0C0A492808099",
 25885 => x"C0C0C0A492808092",
 25886 => x"C0C0C0A492808082",
 25887 => x"C0C0C0A4928080F8",
 25888 => x"C0C0C0A492808080",
 25889 => x"C0C0C0A492808090",
 25890 => x"C0C0C0A4928090C0",
 25891 => x"C0C0C0A4928090F9",
 25892 => x"C0C0C0A4928090A4",
 25893 => x"C0C0C0A4928090B0",
 25894 => x"C0C0C0A492809099",
 25895 => x"C0C0C0A492809092",
 25896 => x"C0C0C0A492809082",
 25897 => x"C0C0C0A4928090F8",
 25898 => x"C0C0C0A492809080",
 25899 => x"C0C0C0A492809090",
 25900 => x"C0C0C0A49290C0C0",
 25901 => x"C0C0C0A49290C0F9",
 25902 => x"C0C0C0A49290C0A4",
 25903 => x"C0C0C0A49290C0B0",
 25904 => x"C0C0C0A49290C099",
 25905 => x"C0C0C0A49290C092",
 25906 => x"C0C0C0A49290C082",
 25907 => x"C0C0C0A49290C0F8",
 25908 => x"C0C0C0A49290C080",
 25909 => x"C0C0C0A49290C090",
 25910 => x"C0C0C0A49290F9C0",
 25911 => x"C0C0C0A49290F9F9",
 25912 => x"C0C0C0A49290F9A4",
 25913 => x"C0C0C0A49290F9B0",
 25914 => x"C0C0C0A49290F999",
 25915 => x"C0C0C0A49290F992",
 25916 => x"C0C0C0A49290F982",
 25917 => x"C0C0C0A49290F9F8",
 25918 => x"C0C0C0A49290F980",
 25919 => x"C0C0C0A49290F990",
 25920 => x"C0C0C0A49290A4C0",
 25921 => x"C0C0C0A49290A4F9",
 25922 => x"C0C0C0A49290A4A4",
 25923 => x"C0C0C0A49290A4B0",
 25924 => x"C0C0C0A49290A499",
 25925 => x"C0C0C0A49290A492",
 25926 => x"C0C0C0A49290A482",
 25927 => x"C0C0C0A49290A4F8",
 25928 => x"C0C0C0A49290A480",
 25929 => x"C0C0C0A49290A490",
 25930 => x"C0C0C0A49290B0C0",
 25931 => x"C0C0C0A49290B0F9",
 25932 => x"C0C0C0A49290B0A4",
 25933 => x"C0C0C0A49290B0B0",
 25934 => x"C0C0C0A49290B099",
 25935 => x"C0C0C0A49290B092",
 25936 => x"C0C0C0A49290B082",
 25937 => x"C0C0C0A49290B0F8",
 25938 => x"C0C0C0A49290B080",
 25939 => x"C0C0C0A49290B090",
 25940 => x"C0C0C0A4929099C0",
 25941 => x"C0C0C0A4929099F9",
 25942 => x"C0C0C0A4929099A4",
 25943 => x"C0C0C0A4929099B0",
 25944 => x"C0C0C0A492909999",
 25945 => x"C0C0C0A492909992",
 25946 => x"C0C0C0A492909982",
 25947 => x"C0C0C0A4929099F8",
 25948 => x"C0C0C0A492909980",
 25949 => x"C0C0C0A492909990",
 25950 => x"C0C0C0A4929092C0",
 25951 => x"C0C0C0A4929092F9",
 25952 => x"C0C0C0A4929092A4",
 25953 => x"C0C0C0A4929092B0",
 25954 => x"C0C0C0A492909299",
 25955 => x"C0C0C0A492909292",
 25956 => x"C0C0C0A492909282",
 25957 => x"C0C0C0A4929092F8",
 25958 => x"C0C0C0A492909280",
 25959 => x"C0C0C0A492909290",
 25960 => x"C0C0C0A4929082C0",
 25961 => x"C0C0C0A4929082F9",
 25962 => x"C0C0C0A4929082A4",
 25963 => x"C0C0C0A4929082B0",
 25964 => x"C0C0C0A492908299",
 25965 => x"C0C0C0A492908292",
 25966 => x"C0C0C0A492908282",
 25967 => x"C0C0C0A4929082F8",
 25968 => x"C0C0C0A492908280",
 25969 => x"C0C0C0A492908290",
 25970 => x"C0C0C0A49290F8C0",
 25971 => x"C0C0C0A49290F8F9",
 25972 => x"C0C0C0A49290F8A4",
 25973 => x"C0C0C0A49290F8B0",
 25974 => x"C0C0C0A49290F899",
 25975 => x"C0C0C0A49290F892",
 25976 => x"C0C0C0A49290F882",
 25977 => x"C0C0C0A49290F8F8",
 25978 => x"C0C0C0A49290F880",
 25979 => x"C0C0C0A49290F890",
 25980 => x"C0C0C0A4929080C0",
 25981 => x"C0C0C0A4929080F9",
 25982 => x"C0C0C0A4929080A4",
 25983 => x"C0C0C0A4929080B0",
 25984 => x"C0C0C0A492908099",
 25985 => x"C0C0C0A492908092",
 25986 => x"C0C0C0A492908082",
 25987 => x"C0C0C0A4929080F8",
 25988 => x"C0C0C0A492908080",
 25989 => x"C0C0C0A492908090",
 25990 => x"C0C0C0A4929090C0",
 25991 => x"C0C0C0A4929090F9",
 25992 => x"C0C0C0A4929090A4",
 25993 => x"C0C0C0A4929090B0",
 25994 => x"C0C0C0A492909099",
 25995 => x"C0C0C0A492909092",
 25996 => x"C0C0C0A492909082",
 25997 => x"C0C0C0A4929090F8",
 25998 => x"C0C0C0A492909080",
 25999 => x"C0C0C0A492909090",
 26000 => x"C0C0C0A482C0C0C0",
 26001 => x"C0C0C0A482C0C0F9",
 26002 => x"C0C0C0A482C0C0A4",
 26003 => x"C0C0C0A482C0C0B0",
 26004 => x"C0C0C0A482C0C099",
 26005 => x"C0C0C0A482C0C092",
 26006 => x"C0C0C0A482C0C082",
 26007 => x"C0C0C0A482C0C0F8",
 26008 => x"C0C0C0A482C0C080",
 26009 => x"C0C0C0A482C0C090",
 26010 => x"C0C0C0A482C0F9C0",
 26011 => x"C0C0C0A482C0F9F9",
 26012 => x"C0C0C0A482C0F9A4",
 26013 => x"C0C0C0A482C0F9B0",
 26014 => x"C0C0C0A482C0F999",
 26015 => x"C0C0C0A482C0F992",
 26016 => x"C0C0C0A482C0F982",
 26017 => x"C0C0C0A482C0F9F8",
 26018 => x"C0C0C0A482C0F980",
 26019 => x"C0C0C0A482C0F990",
 26020 => x"C0C0C0A482C0A4C0",
 26021 => x"C0C0C0A482C0A4F9",
 26022 => x"C0C0C0A482C0A4A4",
 26023 => x"C0C0C0A482C0A4B0",
 26024 => x"C0C0C0A482C0A499",
 26025 => x"C0C0C0A482C0A492",
 26026 => x"C0C0C0A482C0A482",
 26027 => x"C0C0C0A482C0A4F8",
 26028 => x"C0C0C0A482C0A480",
 26029 => x"C0C0C0A482C0A490",
 26030 => x"C0C0C0A482C0B0C0",
 26031 => x"C0C0C0A482C0B0F9",
 26032 => x"C0C0C0A482C0B0A4",
 26033 => x"C0C0C0A482C0B0B0",
 26034 => x"C0C0C0A482C0B099",
 26035 => x"C0C0C0A482C0B092",
 26036 => x"C0C0C0A482C0B082",
 26037 => x"C0C0C0A482C0B0F8",
 26038 => x"C0C0C0A482C0B080",
 26039 => x"C0C0C0A482C0B090",
 26040 => x"C0C0C0A482C099C0",
 26041 => x"C0C0C0A482C099F9",
 26042 => x"C0C0C0A482C099A4",
 26043 => x"C0C0C0A482C099B0",
 26044 => x"C0C0C0A482C09999",
 26045 => x"C0C0C0A482C09992",
 26046 => x"C0C0C0A482C09982",
 26047 => x"C0C0C0A482C099F8",
 26048 => x"C0C0C0A482C09980",
 26049 => x"C0C0C0A482C09990",
 26050 => x"C0C0C0A482C092C0",
 26051 => x"C0C0C0A482C092F9",
 26052 => x"C0C0C0A482C092A4",
 26053 => x"C0C0C0A482C092B0",
 26054 => x"C0C0C0A482C09299",
 26055 => x"C0C0C0A482C09292",
 26056 => x"C0C0C0A482C09282",
 26057 => x"C0C0C0A482C092F8",
 26058 => x"C0C0C0A482C09280",
 26059 => x"C0C0C0A482C09290",
 26060 => x"C0C0C0A482C082C0",
 26061 => x"C0C0C0A482C082F9",
 26062 => x"C0C0C0A482C082A4",
 26063 => x"C0C0C0A482C082B0",
 26064 => x"C0C0C0A482C08299",
 26065 => x"C0C0C0A482C08292",
 26066 => x"C0C0C0A482C08282",
 26067 => x"C0C0C0A482C082F8",
 26068 => x"C0C0C0A482C08280",
 26069 => x"C0C0C0A482C08290",
 26070 => x"C0C0C0A482C0F8C0",
 26071 => x"C0C0C0A482C0F8F9",
 26072 => x"C0C0C0A482C0F8A4",
 26073 => x"C0C0C0A482C0F8B0",
 26074 => x"C0C0C0A482C0F899",
 26075 => x"C0C0C0A482C0F892",
 26076 => x"C0C0C0A482C0F882",
 26077 => x"C0C0C0A482C0F8F8",
 26078 => x"C0C0C0A482C0F880",
 26079 => x"C0C0C0A482C0F890",
 26080 => x"C0C0C0A482C080C0",
 26081 => x"C0C0C0A482C080F9",
 26082 => x"C0C0C0A482C080A4",
 26083 => x"C0C0C0A482C080B0",
 26084 => x"C0C0C0A482C08099",
 26085 => x"C0C0C0A482C08092",
 26086 => x"C0C0C0A482C08082",
 26087 => x"C0C0C0A482C080F8",
 26088 => x"C0C0C0A482C08080",
 26089 => x"C0C0C0A482C08090",
 26090 => x"C0C0C0A482C090C0",
 26091 => x"C0C0C0A482C090F9",
 26092 => x"C0C0C0A482C090A4",
 26093 => x"C0C0C0A482C090B0",
 26094 => x"C0C0C0A482C09099",
 26095 => x"C0C0C0A482C09092",
 26096 => x"C0C0C0A482C09082",
 26097 => x"C0C0C0A482C090F8",
 26098 => x"C0C0C0A482C09080",
 26099 => x"C0C0C0A482C09090",
 26100 => x"C0C0C0A482F9C0C0",
 26101 => x"C0C0C0A482F9C0F9",
 26102 => x"C0C0C0A482F9C0A4",
 26103 => x"C0C0C0A482F9C0B0",
 26104 => x"C0C0C0A482F9C099",
 26105 => x"C0C0C0A482F9C092",
 26106 => x"C0C0C0A482F9C082",
 26107 => x"C0C0C0A482F9C0F8",
 26108 => x"C0C0C0A482F9C080",
 26109 => x"C0C0C0A482F9C090",
 26110 => x"C0C0C0A482F9F9C0",
 26111 => x"C0C0C0A482F9F9F9",
 26112 => x"C0C0C0A482F9F9A4",
 26113 => x"C0C0C0A482F9F9B0",
 26114 => x"C0C0C0A482F9F999",
 26115 => x"C0C0C0A482F9F992",
 26116 => x"C0C0C0A482F9F982",
 26117 => x"C0C0C0A482F9F9F8",
 26118 => x"C0C0C0A482F9F980",
 26119 => x"C0C0C0A482F9F990",
 26120 => x"C0C0C0A482F9A4C0",
 26121 => x"C0C0C0A482F9A4F9",
 26122 => x"C0C0C0A482F9A4A4",
 26123 => x"C0C0C0A482F9A4B0",
 26124 => x"C0C0C0A482F9A499",
 26125 => x"C0C0C0A482F9A492",
 26126 => x"C0C0C0A482F9A482",
 26127 => x"C0C0C0A482F9A4F8",
 26128 => x"C0C0C0A482F9A480",
 26129 => x"C0C0C0A482F9A490",
 26130 => x"C0C0C0A482F9B0C0",
 26131 => x"C0C0C0A482F9B0F9",
 26132 => x"C0C0C0A482F9B0A4",
 26133 => x"C0C0C0A482F9B0B0",
 26134 => x"C0C0C0A482F9B099",
 26135 => x"C0C0C0A482F9B092",
 26136 => x"C0C0C0A482F9B082",
 26137 => x"C0C0C0A482F9B0F8",
 26138 => x"C0C0C0A482F9B080",
 26139 => x"C0C0C0A482F9B090",
 26140 => x"C0C0C0A482F999C0",
 26141 => x"C0C0C0A482F999F9",
 26142 => x"C0C0C0A482F999A4",
 26143 => x"C0C0C0A482F999B0",
 26144 => x"C0C0C0A482F99999",
 26145 => x"C0C0C0A482F99992",
 26146 => x"C0C0C0A482F99982",
 26147 => x"C0C0C0A482F999F8",
 26148 => x"C0C0C0A482F99980",
 26149 => x"C0C0C0A482F99990",
 26150 => x"C0C0C0A482F992C0",
 26151 => x"C0C0C0A482F992F9",
 26152 => x"C0C0C0A482F992A4",
 26153 => x"C0C0C0A482F992B0",
 26154 => x"C0C0C0A482F99299",
 26155 => x"C0C0C0A482F99292",
 26156 => x"C0C0C0A482F99282",
 26157 => x"C0C0C0A482F992F8",
 26158 => x"C0C0C0A482F99280",
 26159 => x"C0C0C0A482F99290",
 26160 => x"C0C0C0A482F982C0",
 26161 => x"C0C0C0A482F982F9",
 26162 => x"C0C0C0A482F982A4",
 26163 => x"C0C0C0A482F982B0",
 26164 => x"C0C0C0A482F98299",
 26165 => x"C0C0C0A482F98292",
 26166 => x"C0C0C0A482F98282",
 26167 => x"C0C0C0A482F982F8",
 26168 => x"C0C0C0A482F98280",
 26169 => x"C0C0C0A482F98290",
 26170 => x"C0C0C0A482F9F8C0",
 26171 => x"C0C0C0A482F9F8F9",
 26172 => x"C0C0C0A482F9F8A4",
 26173 => x"C0C0C0A482F9F8B0",
 26174 => x"C0C0C0A482F9F899",
 26175 => x"C0C0C0A482F9F892",
 26176 => x"C0C0C0A482F9F882",
 26177 => x"C0C0C0A482F9F8F8",
 26178 => x"C0C0C0A482F9F880",
 26179 => x"C0C0C0A482F9F890",
 26180 => x"C0C0C0A482F980C0",
 26181 => x"C0C0C0A482F980F9",
 26182 => x"C0C0C0A482F980A4",
 26183 => x"C0C0C0A482F980B0",
 26184 => x"C0C0C0A482F98099",
 26185 => x"C0C0C0A482F98092",
 26186 => x"C0C0C0A482F98082",
 26187 => x"C0C0C0A482F980F8",
 26188 => x"C0C0C0A482F98080",
 26189 => x"C0C0C0A482F98090",
 26190 => x"C0C0C0A482F990C0",
 26191 => x"C0C0C0A482F990F9",
 26192 => x"C0C0C0A482F990A4",
 26193 => x"C0C0C0A482F990B0",
 26194 => x"C0C0C0A482F99099",
 26195 => x"C0C0C0A482F99092",
 26196 => x"C0C0C0A482F99082",
 26197 => x"C0C0C0A482F990F8",
 26198 => x"C0C0C0A482F99080",
 26199 => x"C0C0C0A482F99090",
 26200 => x"C0C0C0A482A4C0C0",
 26201 => x"C0C0C0A482A4C0F9",
 26202 => x"C0C0C0A482A4C0A4",
 26203 => x"C0C0C0A482A4C0B0",
 26204 => x"C0C0C0A482A4C099",
 26205 => x"C0C0C0A482A4C092",
 26206 => x"C0C0C0A482A4C082",
 26207 => x"C0C0C0A482A4C0F8",
 26208 => x"C0C0C0A482A4C080",
 26209 => x"C0C0C0A482A4C090",
 26210 => x"C0C0C0A482A4F9C0",
 26211 => x"C0C0C0A482A4F9F9",
 26212 => x"C0C0C0A482A4F9A4",
 26213 => x"C0C0C0A482A4F9B0",
 26214 => x"C0C0C0A482A4F999",
 26215 => x"C0C0C0A482A4F992",
 26216 => x"C0C0C0A482A4F982",
 26217 => x"C0C0C0A482A4F9F8",
 26218 => x"C0C0C0A482A4F980",
 26219 => x"C0C0C0A482A4F990",
 26220 => x"C0C0C0A482A4A4C0",
 26221 => x"C0C0C0A482A4A4F9",
 26222 => x"C0C0C0A482A4A4A4",
 26223 => x"C0C0C0A482A4A4B0",
 26224 => x"C0C0C0A482A4A499",
 26225 => x"C0C0C0A482A4A492",
 26226 => x"C0C0C0A482A4A482",
 26227 => x"C0C0C0A482A4A4F8",
 26228 => x"C0C0C0A482A4A480",
 26229 => x"C0C0C0A482A4A490",
 26230 => x"C0C0C0A482A4B0C0",
 26231 => x"C0C0C0A482A4B0F9",
 26232 => x"C0C0C0A482A4B0A4",
 26233 => x"C0C0C0A482A4B0B0",
 26234 => x"C0C0C0A482A4B099",
 26235 => x"C0C0C0A482A4B092",
 26236 => x"C0C0C0A482A4B082",
 26237 => x"C0C0C0A482A4B0F8",
 26238 => x"C0C0C0A482A4B080",
 26239 => x"C0C0C0A482A4B090",
 26240 => x"C0C0C0A482A499C0",
 26241 => x"C0C0C0A482A499F9",
 26242 => x"C0C0C0A482A499A4",
 26243 => x"C0C0C0A482A499B0",
 26244 => x"C0C0C0A482A49999",
 26245 => x"C0C0C0A482A49992",
 26246 => x"C0C0C0A482A49982",
 26247 => x"C0C0C0A482A499F8",
 26248 => x"C0C0C0A482A49980",
 26249 => x"C0C0C0A482A49990",
 26250 => x"C0C0C0A482A492C0",
 26251 => x"C0C0C0A482A492F9",
 26252 => x"C0C0C0A482A492A4",
 26253 => x"C0C0C0A482A492B0",
 26254 => x"C0C0C0A482A49299",
 26255 => x"C0C0C0A482A49292",
 26256 => x"C0C0C0A482A49282",
 26257 => x"C0C0C0A482A492F8",
 26258 => x"C0C0C0A482A49280",
 26259 => x"C0C0C0A482A49290",
 26260 => x"C0C0C0A482A482C0",
 26261 => x"C0C0C0A482A482F9",
 26262 => x"C0C0C0A482A482A4",
 26263 => x"C0C0C0A482A482B0",
 26264 => x"C0C0C0A482A48299",
 26265 => x"C0C0C0A482A48292",
 26266 => x"C0C0C0A482A48282",
 26267 => x"C0C0C0A482A482F8",
 26268 => x"C0C0C0A482A48280",
 26269 => x"C0C0C0A482A48290",
 26270 => x"C0C0C0A482A4F8C0",
 26271 => x"C0C0C0A482A4F8F9",
 26272 => x"C0C0C0A482A4F8A4",
 26273 => x"C0C0C0A482A4F8B0",
 26274 => x"C0C0C0A482A4F899",
 26275 => x"C0C0C0A482A4F892",
 26276 => x"C0C0C0A482A4F882",
 26277 => x"C0C0C0A482A4F8F8",
 26278 => x"C0C0C0A482A4F880",
 26279 => x"C0C0C0A482A4F890",
 26280 => x"C0C0C0A482A480C0",
 26281 => x"C0C0C0A482A480F9",
 26282 => x"C0C0C0A482A480A4",
 26283 => x"C0C0C0A482A480B0",
 26284 => x"C0C0C0A482A48099",
 26285 => x"C0C0C0A482A48092",
 26286 => x"C0C0C0A482A48082",
 26287 => x"C0C0C0A482A480F8",
 26288 => x"C0C0C0A482A48080",
 26289 => x"C0C0C0A482A48090",
 26290 => x"C0C0C0A482A490C0",
 26291 => x"C0C0C0A482A490F9",
 26292 => x"C0C0C0A482A490A4",
 26293 => x"C0C0C0A482A490B0",
 26294 => x"C0C0C0A482A49099",
 26295 => x"C0C0C0A482A49092",
 26296 => x"C0C0C0A482A49082",
 26297 => x"C0C0C0A482A490F8",
 26298 => x"C0C0C0A482A49080",
 26299 => x"C0C0C0A482A49090",
 26300 => x"C0C0C0A482B0C0C0",
 26301 => x"C0C0C0A482B0C0F9",
 26302 => x"C0C0C0A482B0C0A4",
 26303 => x"C0C0C0A482B0C0B0",
 26304 => x"C0C0C0A482B0C099",
 26305 => x"C0C0C0A482B0C092",
 26306 => x"C0C0C0A482B0C082",
 26307 => x"C0C0C0A482B0C0F8",
 26308 => x"C0C0C0A482B0C080",
 26309 => x"C0C0C0A482B0C090",
 26310 => x"C0C0C0A482B0F9C0",
 26311 => x"C0C0C0A482B0F9F9",
 26312 => x"C0C0C0A482B0F9A4",
 26313 => x"C0C0C0A482B0F9B0",
 26314 => x"C0C0C0A482B0F999",
 26315 => x"C0C0C0A482B0F992",
 26316 => x"C0C0C0A482B0F982",
 26317 => x"C0C0C0A482B0F9F8",
 26318 => x"C0C0C0A482B0F980",
 26319 => x"C0C0C0A482B0F990",
 26320 => x"C0C0C0A482B0A4C0",
 26321 => x"C0C0C0A482B0A4F9",
 26322 => x"C0C0C0A482B0A4A4",
 26323 => x"C0C0C0A482B0A4B0",
 26324 => x"C0C0C0A482B0A499",
 26325 => x"C0C0C0A482B0A492",
 26326 => x"C0C0C0A482B0A482",
 26327 => x"C0C0C0A482B0A4F8",
 26328 => x"C0C0C0A482B0A480",
 26329 => x"C0C0C0A482B0A490",
 26330 => x"C0C0C0A482B0B0C0",
 26331 => x"C0C0C0A482B0B0F9",
 26332 => x"C0C0C0A482B0B0A4",
 26333 => x"C0C0C0A482B0B0B0",
 26334 => x"C0C0C0A482B0B099",
 26335 => x"C0C0C0A482B0B092",
 26336 => x"C0C0C0A482B0B082",
 26337 => x"C0C0C0A482B0B0F8",
 26338 => x"C0C0C0A482B0B080",
 26339 => x"C0C0C0A482B0B090",
 26340 => x"C0C0C0A482B099C0",
 26341 => x"C0C0C0A482B099F9",
 26342 => x"C0C0C0A482B099A4",
 26343 => x"C0C0C0A482B099B0",
 26344 => x"C0C0C0A482B09999",
 26345 => x"C0C0C0A482B09992",
 26346 => x"C0C0C0A482B09982",
 26347 => x"C0C0C0A482B099F8",
 26348 => x"C0C0C0A482B09980",
 26349 => x"C0C0C0A482B09990",
 26350 => x"C0C0C0A482B092C0",
 26351 => x"C0C0C0A482B092F9",
 26352 => x"C0C0C0A482B092A4",
 26353 => x"C0C0C0A482B092B0",
 26354 => x"C0C0C0A482B09299",
 26355 => x"C0C0C0A482B09292",
 26356 => x"C0C0C0A482B09282",
 26357 => x"C0C0C0A482B092F8",
 26358 => x"C0C0C0A482B09280",
 26359 => x"C0C0C0A482B09290",
 26360 => x"C0C0C0A482B082C0",
 26361 => x"C0C0C0A482B082F9",
 26362 => x"C0C0C0A482B082A4",
 26363 => x"C0C0C0A482B082B0",
 26364 => x"C0C0C0A482B08299",
 26365 => x"C0C0C0A482B08292",
 26366 => x"C0C0C0A482B08282",
 26367 => x"C0C0C0A482B082F8",
 26368 => x"C0C0C0A482B08280",
 26369 => x"C0C0C0A482B08290",
 26370 => x"C0C0C0A482B0F8C0",
 26371 => x"C0C0C0A482B0F8F9",
 26372 => x"C0C0C0A482B0F8A4",
 26373 => x"C0C0C0A482B0F8B0",
 26374 => x"C0C0C0A482B0F899",
 26375 => x"C0C0C0A482B0F892",
 26376 => x"C0C0C0A482B0F882",
 26377 => x"C0C0C0A482B0F8F8",
 26378 => x"C0C0C0A482B0F880",
 26379 => x"C0C0C0A482B0F890",
 26380 => x"C0C0C0A482B080C0",
 26381 => x"C0C0C0A482B080F9",
 26382 => x"C0C0C0A482B080A4",
 26383 => x"C0C0C0A482B080B0",
 26384 => x"C0C0C0A482B08099",
 26385 => x"C0C0C0A482B08092",
 26386 => x"C0C0C0A482B08082",
 26387 => x"C0C0C0A482B080F8",
 26388 => x"C0C0C0A482B08080",
 26389 => x"C0C0C0A482B08090",
 26390 => x"C0C0C0A482B090C0",
 26391 => x"C0C0C0A482B090F9",
 26392 => x"C0C0C0A482B090A4",
 26393 => x"C0C0C0A482B090B0",
 26394 => x"C0C0C0A482B09099",
 26395 => x"C0C0C0A482B09092",
 26396 => x"C0C0C0A482B09082",
 26397 => x"C0C0C0A482B090F8",
 26398 => x"C0C0C0A482B09080",
 26399 => x"C0C0C0A482B09090",
 26400 => x"C0C0C0A48299C0C0",
 26401 => x"C0C0C0A48299C0F9",
 26402 => x"C0C0C0A48299C0A4",
 26403 => x"C0C0C0A48299C0B0",
 26404 => x"C0C0C0A48299C099",
 26405 => x"C0C0C0A48299C092",
 26406 => x"C0C0C0A48299C082",
 26407 => x"C0C0C0A48299C0F8",
 26408 => x"C0C0C0A48299C080",
 26409 => x"C0C0C0A48299C090",
 26410 => x"C0C0C0A48299F9C0",
 26411 => x"C0C0C0A48299F9F9",
 26412 => x"C0C0C0A48299F9A4",
 26413 => x"C0C0C0A48299F9B0",
 26414 => x"C0C0C0A48299F999",
 26415 => x"C0C0C0A48299F992",
 26416 => x"C0C0C0A48299F982",
 26417 => x"C0C0C0A48299F9F8",
 26418 => x"C0C0C0A48299F980",
 26419 => x"C0C0C0A48299F990",
 26420 => x"C0C0C0A48299A4C0",
 26421 => x"C0C0C0A48299A4F9",
 26422 => x"C0C0C0A48299A4A4",
 26423 => x"C0C0C0A48299A4B0",
 26424 => x"C0C0C0A48299A499",
 26425 => x"C0C0C0A48299A492",
 26426 => x"C0C0C0A48299A482",
 26427 => x"C0C0C0A48299A4F8",
 26428 => x"C0C0C0A48299A480",
 26429 => x"C0C0C0A48299A490",
 26430 => x"C0C0C0A48299B0C0",
 26431 => x"C0C0C0A48299B0F9",
 26432 => x"C0C0C0A48299B0A4",
 26433 => x"C0C0C0A48299B0B0",
 26434 => x"C0C0C0A48299B099",
 26435 => x"C0C0C0A48299B092",
 26436 => x"C0C0C0A48299B082",
 26437 => x"C0C0C0A48299B0F8",
 26438 => x"C0C0C0A48299B080",
 26439 => x"C0C0C0A48299B090",
 26440 => x"C0C0C0A4829999C0",
 26441 => x"C0C0C0A4829999F9",
 26442 => x"C0C0C0A4829999A4",
 26443 => x"C0C0C0A4829999B0",
 26444 => x"C0C0C0A482999999",
 26445 => x"C0C0C0A482999992",
 26446 => x"C0C0C0A482999982",
 26447 => x"C0C0C0A4829999F8",
 26448 => x"C0C0C0A482999980",
 26449 => x"C0C0C0A482999990",
 26450 => x"C0C0C0A4829992C0",
 26451 => x"C0C0C0A4829992F9",
 26452 => x"C0C0C0A4829992A4",
 26453 => x"C0C0C0A4829992B0",
 26454 => x"C0C0C0A482999299",
 26455 => x"C0C0C0A482999292",
 26456 => x"C0C0C0A482999282",
 26457 => x"C0C0C0A4829992F8",
 26458 => x"C0C0C0A482999280",
 26459 => x"C0C0C0A482999290",
 26460 => x"C0C0C0A4829982C0",
 26461 => x"C0C0C0A4829982F9",
 26462 => x"C0C0C0A4829982A4",
 26463 => x"C0C0C0A4829982B0",
 26464 => x"C0C0C0A482998299",
 26465 => x"C0C0C0A482998292",
 26466 => x"C0C0C0A482998282",
 26467 => x"C0C0C0A4829982F8",
 26468 => x"C0C0C0A482998280",
 26469 => x"C0C0C0A482998290",
 26470 => x"C0C0C0A48299F8C0",
 26471 => x"C0C0C0A48299F8F9",
 26472 => x"C0C0C0A48299F8A4",
 26473 => x"C0C0C0A48299F8B0",
 26474 => x"C0C0C0A48299F899",
 26475 => x"C0C0C0A48299F892",
 26476 => x"C0C0C0A48299F882",
 26477 => x"C0C0C0A48299F8F8",
 26478 => x"C0C0C0A48299F880",
 26479 => x"C0C0C0A48299F890",
 26480 => x"C0C0C0A4829980C0",
 26481 => x"C0C0C0A4829980F9",
 26482 => x"C0C0C0A4829980A4",
 26483 => x"C0C0C0A4829980B0",
 26484 => x"C0C0C0A482998099",
 26485 => x"C0C0C0A482998092",
 26486 => x"C0C0C0A482998082",
 26487 => x"C0C0C0A4829980F8",
 26488 => x"C0C0C0A482998080",
 26489 => x"C0C0C0A482998090",
 26490 => x"C0C0C0A4829990C0",
 26491 => x"C0C0C0A4829990F9",
 26492 => x"C0C0C0A4829990A4",
 26493 => x"C0C0C0A4829990B0",
 26494 => x"C0C0C0A482999099",
 26495 => x"C0C0C0A482999092",
 26496 => x"C0C0C0A482999082",
 26497 => x"C0C0C0A4829990F8",
 26498 => x"C0C0C0A482999080",
 26499 => x"C0C0C0A482999090",
 26500 => x"C0C0C0A48292C0C0",
 26501 => x"C0C0C0A48292C0F9",
 26502 => x"C0C0C0A48292C0A4",
 26503 => x"C0C0C0A48292C0B0",
 26504 => x"C0C0C0A48292C099",
 26505 => x"C0C0C0A48292C092",
 26506 => x"C0C0C0A48292C082",
 26507 => x"C0C0C0A48292C0F8",
 26508 => x"C0C0C0A48292C080",
 26509 => x"C0C0C0A48292C090",
 26510 => x"C0C0C0A48292F9C0",
 26511 => x"C0C0C0A48292F9F9",
 26512 => x"C0C0C0A48292F9A4",
 26513 => x"C0C0C0A48292F9B0",
 26514 => x"C0C0C0A48292F999",
 26515 => x"C0C0C0A48292F992",
 26516 => x"C0C0C0A48292F982",
 26517 => x"C0C0C0A48292F9F8",
 26518 => x"C0C0C0A48292F980",
 26519 => x"C0C0C0A48292F990",
 26520 => x"C0C0C0A48292A4C0",
 26521 => x"C0C0C0A48292A4F9",
 26522 => x"C0C0C0A48292A4A4",
 26523 => x"C0C0C0A48292A4B0",
 26524 => x"C0C0C0A48292A499",
 26525 => x"C0C0C0A48292A492",
 26526 => x"C0C0C0A48292A482",
 26527 => x"C0C0C0A48292A4F8",
 26528 => x"C0C0C0A48292A480",
 26529 => x"C0C0C0A48292A490",
 26530 => x"C0C0C0A48292B0C0",
 26531 => x"C0C0C0A48292B0F9",
 26532 => x"C0C0C0A48292B0A4",
 26533 => x"C0C0C0A48292B0B0",
 26534 => x"C0C0C0A48292B099",
 26535 => x"C0C0C0A48292B092",
 26536 => x"C0C0C0A48292B082",
 26537 => x"C0C0C0A48292B0F8",
 26538 => x"C0C0C0A48292B080",
 26539 => x"C0C0C0A48292B090",
 26540 => x"C0C0C0A4829299C0",
 26541 => x"C0C0C0A4829299F9",
 26542 => x"C0C0C0A4829299A4",
 26543 => x"C0C0C0A4829299B0",
 26544 => x"C0C0C0A482929999",
 26545 => x"C0C0C0A482929992",
 26546 => x"C0C0C0A482929982",
 26547 => x"C0C0C0A4829299F8",
 26548 => x"C0C0C0A482929980",
 26549 => x"C0C0C0A482929990",
 26550 => x"C0C0C0A4829292C0",
 26551 => x"C0C0C0A4829292F9",
 26552 => x"C0C0C0A4829292A4",
 26553 => x"C0C0C0A4829292B0",
 26554 => x"C0C0C0A482929299",
 26555 => x"C0C0C0A482929292",
 26556 => x"C0C0C0A482929282",
 26557 => x"C0C0C0A4829292F8",
 26558 => x"C0C0C0A482929280",
 26559 => x"C0C0C0A482929290",
 26560 => x"C0C0C0A4829282C0",
 26561 => x"C0C0C0A4829282F9",
 26562 => x"C0C0C0A4829282A4",
 26563 => x"C0C0C0A4829282B0",
 26564 => x"C0C0C0A482928299",
 26565 => x"C0C0C0A482928292",
 26566 => x"C0C0C0A482928282",
 26567 => x"C0C0C0A4829282F8",
 26568 => x"C0C0C0A482928280",
 26569 => x"C0C0C0A482928290",
 26570 => x"C0C0C0A48292F8C0",
 26571 => x"C0C0C0A48292F8F9",
 26572 => x"C0C0C0A48292F8A4",
 26573 => x"C0C0C0A48292F8B0",
 26574 => x"C0C0C0A48292F899",
 26575 => x"C0C0C0A48292F892",
 26576 => x"C0C0C0A48292F882",
 26577 => x"C0C0C0A48292F8F8",
 26578 => x"C0C0C0A48292F880",
 26579 => x"C0C0C0A48292F890",
 26580 => x"C0C0C0A4829280C0",
 26581 => x"C0C0C0A4829280F9",
 26582 => x"C0C0C0A4829280A4",
 26583 => x"C0C0C0A4829280B0",
 26584 => x"C0C0C0A482928099",
 26585 => x"C0C0C0A482928092",
 26586 => x"C0C0C0A482928082",
 26587 => x"C0C0C0A4829280F8",
 26588 => x"C0C0C0A482928080",
 26589 => x"C0C0C0A482928090",
 26590 => x"C0C0C0A4829290C0",
 26591 => x"C0C0C0A4829290F9",
 26592 => x"C0C0C0A4829290A4",
 26593 => x"C0C0C0A4829290B0",
 26594 => x"C0C0C0A482929099",
 26595 => x"C0C0C0A482929092",
 26596 => x"C0C0C0A482929082",
 26597 => x"C0C0C0A4829290F8",
 26598 => x"C0C0C0A482929080",
 26599 => x"C0C0C0A482929090",
 26600 => x"C0C0C0A48282C0C0",
 26601 => x"C0C0C0A48282C0F9",
 26602 => x"C0C0C0A48282C0A4",
 26603 => x"C0C0C0A48282C0B0",
 26604 => x"C0C0C0A48282C099",
 26605 => x"C0C0C0A48282C092",
 26606 => x"C0C0C0A48282C082",
 26607 => x"C0C0C0A48282C0F8",
 26608 => x"C0C0C0A48282C080",
 26609 => x"C0C0C0A48282C090",
 26610 => x"C0C0C0A48282F9C0",
 26611 => x"C0C0C0A48282F9F9",
 26612 => x"C0C0C0A48282F9A4",
 26613 => x"C0C0C0A48282F9B0",
 26614 => x"C0C0C0A48282F999",
 26615 => x"C0C0C0A48282F992",
 26616 => x"C0C0C0A48282F982",
 26617 => x"C0C0C0A48282F9F8",
 26618 => x"C0C0C0A48282F980",
 26619 => x"C0C0C0A48282F990",
 26620 => x"C0C0C0A48282A4C0",
 26621 => x"C0C0C0A48282A4F9",
 26622 => x"C0C0C0A48282A4A4",
 26623 => x"C0C0C0A48282A4B0",
 26624 => x"C0C0C0A48282A499",
 26625 => x"C0C0C0A48282A492",
 26626 => x"C0C0C0A48282A482",
 26627 => x"C0C0C0A48282A4F8",
 26628 => x"C0C0C0A48282A480",
 26629 => x"C0C0C0A48282A490",
 26630 => x"C0C0C0A48282B0C0",
 26631 => x"C0C0C0A48282B0F9",
 26632 => x"C0C0C0A48282B0A4",
 26633 => x"C0C0C0A48282B0B0",
 26634 => x"C0C0C0A48282B099",
 26635 => x"C0C0C0A48282B092",
 26636 => x"C0C0C0A48282B082",
 26637 => x"C0C0C0A48282B0F8",
 26638 => x"C0C0C0A48282B080",
 26639 => x"C0C0C0A48282B090",
 26640 => x"C0C0C0A4828299C0",
 26641 => x"C0C0C0A4828299F9",
 26642 => x"C0C0C0A4828299A4",
 26643 => x"C0C0C0A4828299B0",
 26644 => x"C0C0C0A482829999",
 26645 => x"C0C0C0A482829992",
 26646 => x"C0C0C0A482829982",
 26647 => x"C0C0C0A4828299F8",
 26648 => x"C0C0C0A482829980",
 26649 => x"C0C0C0A482829990",
 26650 => x"C0C0C0A4828292C0",
 26651 => x"C0C0C0A4828292F9",
 26652 => x"C0C0C0A4828292A4",
 26653 => x"C0C0C0A4828292B0",
 26654 => x"C0C0C0A482829299",
 26655 => x"C0C0C0A482829292",
 26656 => x"C0C0C0A482829282",
 26657 => x"C0C0C0A4828292F8",
 26658 => x"C0C0C0A482829280",
 26659 => x"C0C0C0A482829290",
 26660 => x"C0C0C0A4828282C0",
 26661 => x"C0C0C0A4828282F9",
 26662 => x"C0C0C0A4828282A4",
 26663 => x"C0C0C0A4828282B0",
 26664 => x"C0C0C0A482828299",
 26665 => x"C0C0C0A482828292",
 26666 => x"C0C0C0A482828282",
 26667 => x"C0C0C0A4828282F8",
 26668 => x"C0C0C0A482828280",
 26669 => x"C0C0C0A482828290",
 26670 => x"C0C0C0A48282F8C0",
 26671 => x"C0C0C0A48282F8F9",
 26672 => x"C0C0C0A48282F8A4",
 26673 => x"C0C0C0A48282F8B0",
 26674 => x"C0C0C0A48282F899",
 26675 => x"C0C0C0A48282F892",
 26676 => x"C0C0C0A48282F882",
 26677 => x"C0C0C0A48282F8F8",
 26678 => x"C0C0C0A48282F880",
 26679 => x"C0C0C0A48282F890",
 26680 => x"C0C0C0A4828280C0",
 26681 => x"C0C0C0A4828280F9",
 26682 => x"C0C0C0A4828280A4",
 26683 => x"C0C0C0A4828280B0",
 26684 => x"C0C0C0A482828099",
 26685 => x"C0C0C0A482828092",
 26686 => x"C0C0C0A482828082",
 26687 => x"C0C0C0A4828280F8",
 26688 => x"C0C0C0A482828080",
 26689 => x"C0C0C0A482828090",
 26690 => x"C0C0C0A4828290C0",
 26691 => x"C0C0C0A4828290F9",
 26692 => x"C0C0C0A4828290A4",
 26693 => x"C0C0C0A4828290B0",
 26694 => x"C0C0C0A482829099",
 26695 => x"C0C0C0A482829092",
 26696 => x"C0C0C0A482829082",
 26697 => x"C0C0C0A4828290F8",
 26698 => x"C0C0C0A482829080",
 26699 => x"C0C0C0A482829090",
 26700 => x"C0C0C0A482F8C0C0",
 26701 => x"C0C0C0A482F8C0F9",
 26702 => x"C0C0C0A482F8C0A4",
 26703 => x"C0C0C0A482F8C0B0",
 26704 => x"C0C0C0A482F8C099",
 26705 => x"C0C0C0A482F8C092",
 26706 => x"C0C0C0A482F8C082",
 26707 => x"C0C0C0A482F8C0F8",
 26708 => x"C0C0C0A482F8C080",
 26709 => x"C0C0C0A482F8C090",
 26710 => x"C0C0C0A482F8F9C0",
 26711 => x"C0C0C0A482F8F9F9",
 26712 => x"C0C0C0A482F8F9A4",
 26713 => x"C0C0C0A482F8F9B0",
 26714 => x"C0C0C0A482F8F999",
 26715 => x"C0C0C0A482F8F992",
 26716 => x"C0C0C0A482F8F982",
 26717 => x"C0C0C0A482F8F9F8",
 26718 => x"C0C0C0A482F8F980",
 26719 => x"C0C0C0A482F8F990",
 26720 => x"C0C0C0A482F8A4C0",
 26721 => x"C0C0C0A482F8A4F9",
 26722 => x"C0C0C0A482F8A4A4",
 26723 => x"C0C0C0A482F8A4B0",
 26724 => x"C0C0C0A482F8A499",
 26725 => x"C0C0C0A482F8A492",
 26726 => x"C0C0C0A482F8A482",
 26727 => x"C0C0C0A482F8A4F8",
 26728 => x"C0C0C0A482F8A480",
 26729 => x"C0C0C0A482F8A490",
 26730 => x"C0C0C0A482F8B0C0",
 26731 => x"C0C0C0A482F8B0F9",
 26732 => x"C0C0C0A482F8B0A4",
 26733 => x"C0C0C0A482F8B0B0",
 26734 => x"C0C0C0A482F8B099",
 26735 => x"C0C0C0A482F8B092",
 26736 => x"C0C0C0A482F8B082",
 26737 => x"C0C0C0A482F8B0F8",
 26738 => x"C0C0C0A482F8B080",
 26739 => x"C0C0C0A482F8B090",
 26740 => x"C0C0C0A482F899C0",
 26741 => x"C0C0C0A482F899F9",
 26742 => x"C0C0C0A482F899A4",
 26743 => x"C0C0C0A482F899B0",
 26744 => x"C0C0C0A482F89999",
 26745 => x"C0C0C0A482F89992",
 26746 => x"C0C0C0A482F89982",
 26747 => x"C0C0C0A482F899F8",
 26748 => x"C0C0C0A482F89980",
 26749 => x"C0C0C0A482F89990",
 26750 => x"C0C0C0A482F892C0",
 26751 => x"C0C0C0A482F892F9",
 26752 => x"C0C0C0A482F892A4",
 26753 => x"C0C0C0A482F892B0",
 26754 => x"C0C0C0A482F89299",
 26755 => x"C0C0C0A482F89292",
 26756 => x"C0C0C0A482F89282",
 26757 => x"C0C0C0A482F892F8",
 26758 => x"C0C0C0A482F89280",
 26759 => x"C0C0C0A482F89290",
 26760 => x"C0C0C0A482F882C0",
 26761 => x"C0C0C0A482F882F9",
 26762 => x"C0C0C0A482F882A4",
 26763 => x"C0C0C0A482F882B0",
 26764 => x"C0C0C0A482F88299",
 26765 => x"C0C0C0A482F88292",
 26766 => x"C0C0C0A482F88282",
 26767 => x"C0C0C0A482F882F8",
 26768 => x"C0C0C0A482F88280",
 26769 => x"C0C0C0A482F88290",
 26770 => x"C0C0C0A482F8F8C0",
 26771 => x"C0C0C0A482F8F8F9",
 26772 => x"C0C0C0A482F8F8A4",
 26773 => x"C0C0C0A482F8F8B0",
 26774 => x"C0C0C0A482F8F899",
 26775 => x"C0C0C0A482F8F892",
 26776 => x"C0C0C0A482F8F882",
 26777 => x"C0C0C0A482F8F8F8",
 26778 => x"C0C0C0A482F8F880",
 26779 => x"C0C0C0A482F8F890",
 26780 => x"C0C0C0A482F880C0",
 26781 => x"C0C0C0A482F880F9",
 26782 => x"C0C0C0A482F880A4",
 26783 => x"C0C0C0A482F880B0",
 26784 => x"C0C0C0A482F88099",
 26785 => x"C0C0C0A482F88092",
 26786 => x"C0C0C0A482F88082",
 26787 => x"C0C0C0A482F880F8",
 26788 => x"C0C0C0A482F88080",
 26789 => x"C0C0C0A482F88090",
 26790 => x"C0C0C0A482F890C0",
 26791 => x"C0C0C0A482F890F9",
 26792 => x"C0C0C0A482F890A4",
 26793 => x"C0C0C0A482F890B0",
 26794 => x"C0C0C0A482F89099",
 26795 => x"C0C0C0A482F89092",
 26796 => x"C0C0C0A482F89082",
 26797 => x"C0C0C0A482F890F8",
 26798 => x"C0C0C0A482F89080",
 26799 => x"C0C0C0A482F89090",
 26800 => x"C0C0C0A48280C0C0",
 26801 => x"C0C0C0A48280C0F9",
 26802 => x"C0C0C0A48280C0A4",
 26803 => x"C0C0C0A48280C0B0",
 26804 => x"C0C0C0A48280C099",
 26805 => x"C0C0C0A48280C092",
 26806 => x"C0C0C0A48280C082",
 26807 => x"C0C0C0A48280C0F8",
 26808 => x"C0C0C0A48280C080",
 26809 => x"C0C0C0A48280C090",
 26810 => x"C0C0C0A48280F9C0",
 26811 => x"C0C0C0A48280F9F9",
 26812 => x"C0C0C0A48280F9A4",
 26813 => x"C0C0C0A48280F9B0",
 26814 => x"C0C0C0A48280F999",
 26815 => x"C0C0C0A48280F992",
 26816 => x"C0C0C0A48280F982",
 26817 => x"C0C0C0A48280F9F8",
 26818 => x"C0C0C0A48280F980",
 26819 => x"C0C0C0A48280F990",
 26820 => x"C0C0C0A48280A4C0",
 26821 => x"C0C0C0A48280A4F9",
 26822 => x"C0C0C0A48280A4A4",
 26823 => x"C0C0C0A48280A4B0",
 26824 => x"C0C0C0A48280A499",
 26825 => x"C0C0C0A48280A492",
 26826 => x"C0C0C0A48280A482",
 26827 => x"C0C0C0A48280A4F8",
 26828 => x"C0C0C0A48280A480",
 26829 => x"C0C0C0A48280A490",
 26830 => x"C0C0C0A48280B0C0",
 26831 => x"C0C0C0A48280B0F9",
 26832 => x"C0C0C0A48280B0A4",
 26833 => x"C0C0C0A48280B0B0",
 26834 => x"C0C0C0A48280B099",
 26835 => x"C0C0C0A48280B092",
 26836 => x"C0C0C0A48280B082",
 26837 => x"C0C0C0A48280B0F8",
 26838 => x"C0C0C0A48280B080",
 26839 => x"C0C0C0A48280B090",
 26840 => x"C0C0C0A4828099C0",
 26841 => x"C0C0C0A4828099F9",
 26842 => x"C0C0C0A4828099A4",
 26843 => x"C0C0C0A4828099B0",
 26844 => x"C0C0C0A482809999",
 26845 => x"C0C0C0A482809992",
 26846 => x"C0C0C0A482809982",
 26847 => x"C0C0C0A4828099F8",
 26848 => x"C0C0C0A482809980",
 26849 => x"C0C0C0A482809990",
 26850 => x"C0C0C0A4828092C0",
 26851 => x"C0C0C0A4828092F9",
 26852 => x"C0C0C0A4828092A4",
 26853 => x"C0C0C0A4828092B0",
 26854 => x"C0C0C0A482809299",
 26855 => x"C0C0C0A482809292",
 26856 => x"C0C0C0A482809282",
 26857 => x"C0C0C0A4828092F8",
 26858 => x"C0C0C0A482809280",
 26859 => x"C0C0C0A482809290",
 26860 => x"C0C0C0A4828082C0",
 26861 => x"C0C0C0A4828082F9",
 26862 => x"C0C0C0A4828082A4",
 26863 => x"C0C0C0A4828082B0",
 26864 => x"C0C0C0A482808299",
 26865 => x"C0C0C0A482808292",
 26866 => x"C0C0C0A482808282",
 26867 => x"C0C0C0A4828082F8",
 26868 => x"C0C0C0A482808280",
 26869 => x"C0C0C0A482808290",
 26870 => x"C0C0C0A48280F8C0",
 26871 => x"C0C0C0A48280F8F9",
 26872 => x"C0C0C0A48280F8A4",
 26873 => x"C0C0C0A48280F8B0",
 26874 => x"C0C0C0A48280F899",
 26875 => x"C0C0C0A48280F892",
 26876 => x"C0C0C0A48280F882",
 26877 => x"C0C0C0A48280F8F8",
 26878 => x"C0C0C0A48280F880",
 26879 => x"C0C0C0A48280F890",
 26880 => x"C0C0C0A4828080C0",
 26881 => x"C0C0C0A4828080F9",
 26882 => x"C0C0C0A4828080A4",
 26883 => x"C0C0C0A4828080B0",
 26884 => x"C0C0C0A482808099",
 26885 => x"C0C0C0A482808092",
 26886 => x"C0C0C0A482808082",
 26887 => x"C0C0C0A4828080F8",
 26888 => x"C0C0C0A482808080",
 26889 => x"C0C0C0A482808090",
 26890 => x"C0C0C0A4828090C0",
 26891 => x"C0C0C0A4828090F9",
 26892 => x"C0C0C0A4828090A4",
 26893 => x"C0C0C0A4828090B0",
 26894 => x"C0C0C0A482809099",
 26895 => x"C0C0C0A482809092",
 26896 => x"C0C0C0A482809082",
 26897 => x"C0C0C0A4828090F8",
 26898 => x"C0C0C0A482809080",
 26899 => x"C0C0C0A482809090",
 26900 => x"C0C0C0A48290C0C0",
 26901 => x"C0C0C0A48290C0F9",
 26902 => x"C0C0C0A48290C0A4",
 26903 => x"C0C0C0A48290C0B0",
 26904 => x"C0C0C0A48290C099",
 26905 => x"C0C0C0A48290C092",
 26906 => x"C0C0C0A48290C082",
 26907 => x"C0C0C0A48290C0F8",
 26908 => x"C0C0C0A48290C080",
 26909 => x"C0C0C0A48290C090",
 26910 => x"C0C0C0A48290F9C0",
 26911 => x"C0C0C0A48290F9F9",
 26912 => x"C0C0C0A48290F9A4",
 26913 => x"C0C0C0A48290F9B0",
 26914 => x"C0C0C0A48290F999",
 26915 => x"C0C0C0A48290F992",
 26916 => x"C0C0C0A48290F982",
 26917 => x"C0C0C0A48290F9F8",
 26918 => x"C0C0C0A48290F980",
 26919 => x"C0C0C0A48290F990",
 26920 => x"C0C0C0A48290A4C0",
 26921 => x"C0C0C0A48290A4F9",
 26922 => x"C0C0C0A48290A4A4",
 26923 => x"C0C0C0A48290A4B0",
 26924 => x"C0C0C0A48290A499",
 26925 => x"C0C0C0A48290A492",
 26926 => x"C0C0C0A48290A482",
 26927 => x"C0C0C0A48290A4F8",
 26928 => x"C0C0C0A48290A480",
 26929 => x"C0C0C0A48290A490",
 26930 => x"C0C0C0A48290B0C0",
 26931 => x"C0C0C0A48290B0F9",
 26932 => x"C0C0C0A48290B0A4",
 26933 => x"C0C0C0A48290B0B0",
 26934 => x"C0C0C0A48290B099",
 26935 => x"C0C0C0A48290B092",
 26936 => x"C0C0C0A48290B082",
 26937 => x"C0C0C0A48290B0F8",
 26938 => x"C0C0C0A48290B080",
 26939 => x"C0C0C0A48290B090",
 26940 => x"C0C0C0A4829099C0",
 26941 => x"C0C0C0A4829099F9",
 26942 => x"C0C0C0A4829099A4",
 26943 => x"C0C0C0A4829099B0",
 26944 => x"C0C0C0A482909999",
 26945 => x"C0C0C0A482909992",
 26946 => x"C0C0C0A482909982",
 26947 => x"C0C0C0A4829099F8",
 26948 => x"C0C0C0A482909980",
 26949 => x"C0C0C0A482909990",
 26950 => x"C0C0C0A4829092C0",
 26951 => x"C0C0C0A4829092F9",
 26952 => x"C0C0C0A4829092A4",
 26953 => x"C0C0C0A4829092B0",
 26954 => x"C0C0C0A482909299",
 26955 => x"C0C0C0A482909292",
 26956 => x"C0C0C0A482909282",
 26957 => x"C0C0C0A4829092F8",
 26958 => x"C0C0C0A482909280",
 26959 => x"C0C0C0A482909290",
 26960 => x"C0C0C0A4829082C0",
 26961 => x"C0C0C0A4829082F9",
 26962 => x"C0C0C0A4829082A4",
 26963 => x"C0C0C0A4829082B0",
 26964 => x"C0C0C0A482908299",
 26965 => x"C0C0C0A482908292",
 26966 => x"C0C0C0A482908282",
 26967 => x"C0C0C0A4829082F8",
 26968 => x"C0C0C0A482908280",
 26969 => x"C0C0C0A482908290",
 26970 => x"C0C0C0A48290F8C0",
 26971 => x"C0C0C0A48290F8F9",
 26972 => x"C0C0C0A48290F8A4",
 26973 => x"C0C0C0A48290F8B0",
 26974 => x"C0C0C0A48290F899",
 26975 => x"C0C0C0A48290F892",
 26976 => x"C0C0C0A48290F882",
 26977 => x"C0C0C0A48290F8F8",
 26978 => x"C0C0C0A48290F880",
 26979 => x"C0C0C0A48290F890",
 26980 => x"C0C0C0A4829080C0",
 26981 => x"C0C0C0A4829080F9",
 26982 => x"C0C0C0A4829080A4",
 26983 => x"C0C0C0A4829080B0",
 26984 => x"C0C0C0A482908099",
 26985 => x"C0C0C0A482908092",
 26986 => x"C0C0C0A482908082",
 26987 => x"C0C0C0A4829080F8",
 26988 => x"C0C0C0A482908080",
 26989 => x"C0C0C0A482908090",
 26990 => x"C0C0C0A4829090C0",
 26991 => x"C0C0C0A4829090F9",
 26992 => x"C0C0C0A4829090A4",
 26993 => x"C0C0C0A4829090B0",
 26994 => x"C0C0C0A482909099",
 26995 => x"C0C0C0A482909092",
 26996 => x"C0C0C0A482909082",
 26997 => x"C0C0C0A4829090F8",
 26998 => x"C0C0C0A482909080",
 26999 => x"C0C0C0A482909090",
 27000 => x"C0C0C0A4F8C0C0C0",
 27001 => x"C0C0C0A4F8C0C0F9",
 27002 => x"C0C0C0A4F8C0C0A4",
 27003 => x"C0C0C0A4F8C0C0B0",
 27004 => x"C0C0C0A4F8C0C099",
 27005 => x"C0C0C0A4F8C0C092",
 27006 => x"C0C0C0A4F8C0C082",
 27007 => x"C0C0C0A4F8C0C0F8",
 27008 => x"C0C0C0A4F8C0C080",
 27009 => x"C0C0C0A4F8C0C090",
 27010 => x"C0C0C0A4F8C0F9C0",
 27011 => x"C0C0C0A4F8C0F9F9",
 27012 => x"C0C0C0A4F8C0F9A4",
 27013 => x"C0C0C0A4F8C0F9B0",
 27014 => x"C0C0C0A4F8C0F999",
 27015 => x"C0C0C0A4F8C0F992",
 27016 => x"C0C0C0A4F8C0F982",
 27017 => x"C0C0C0A4F8C0F9F8",
 27018 => x"C0C0C0A4F8C0F980",
 27019 => x"C0C0C0A4F8C0F990",
 27020 => x"C0C0C0A4F8C0A4C0",
 27021 => x"C0C0C0A4F8C0A4F9",
 27022 => x"C0C0C0A4F8C0A4A4",
 27023 => x"C0C0C0A4F8C0A4B0",
 27024 => x"C0C0C0A4F8C0A499",
 27025 => x"C0C0C0A4F8C0A492",
 27026 => x"C0C0C0A4F8C0A482",
 27027 => x"C0C0C0A4F8C0A4F8",
 27028 => x"C0C0C0A4F8C0A480",
 27029 => x"C0C0C0A4F8C0A490",
 27030 => x"C0C0C0A4F8C0B0C0",
 27031 => x"C0C0C0A4F8C0B0F9",
 27032 => x"C0C0C0A4F8C0B0A4",
 27033 => x"C0C0C0A4F8C0B0B0",
 27034 => x"C0C0C0A4F8C0B099",
 27035 => x"C0C0C0A4F8C0B092",
 27036 => x"C0C0C0A4F8C0B082",
 27037 => x"C0C0C0A4F8C0B0F8",
 27038 => x"C0C0C0A4F8C0B080",
 27039 => x"C0C0C0A4F8C0B090",
 27040 => x"C0C0C0A4F8C099C0",
 27041 => x"C0C0C0A4F8C099F9",
 27042 => x"C0C0C0A4F8C099A4",
 27043 => x"C0C0C0A4F8C099B0",
 27044 => x"C0C0C0A4F8C09999",
 27045 => x"C0C0C0A4F8C09992",
 27046 => x"C0C0C0A4F8C09982",
 27047 => x"C0C0C0A4F8C099F8",
 27048 => x"C0C0C0A4F8C09980",
 27049 => x"C0C0C0A4F8C09990",
 27050 => x"C0C0C0A4F8C092C0",
 27051 => x"C0C0C0A4F8C092F9",
 27052 => x"C0C0C0A4F8C092A4",
 27053 => x"C0C0C0A4F8C092B0",
 27054 => x"C0C0C0A4F8C09299",
 27055 => x"C0C0C0A4F8C09292",
 27056 => x"C0C0C0A4F8C09282",
 27057 => x"C0C0C0A4F8C092F8",
 27058 => x"C0C0C0A4F8C09280",
 27059 => x"C0C0C0A4F8C09290",
 27060 => x"C0C0C0A4F8C082C0",
 27061 => x"C0C0C0A4F8C082F9",
 27062 => x"C0C0C0A4F8C082A4",
 27063 => x"C0C0C0A4F8C082B0",
 27064 => x"C0C0C0A4F8C08299",
 27065 => x"C0C0C0A4F8C08292",
 27066 => x"C0C0C0A4F8C08282",
 27067 => x"C0C0C0A4F8C082F8",
 27068 => x"C0C0C0A4F8C08280",
 27069 => x"C0C0C0A4F8C08290",
 27070 => x"C0C0C0A4F8C0F8C0",
 27071 => x"C0C0C0A4F8C0F8F9",
 27072 => x"C0C0C0A4F8C0F8A4",
 27073 => x"C0C0C0A4F8C0F8B0",
 27074 => x"C0C0C0A4F8C0F899",
 27075 => x"C0C0C0A4F8C0F892",
 27076 => x"C0C0C0A4F8C0F882",
 27077 => x"C0C0C0A4F8C0F8F8",
 27078 => x"C0C0C0A4F8C0F880",
 27079 => x"C0C0C0A4F8C0F890",
 27080 => x"C0C0C0A4F8C080C0",
 27081 => x"C0C0C0A4F8C080F9",
 27082 => x"C0C0C0A4F8C080A4",
 27083 => x"C0C0C0A4F8C080B0",
 27084 => x"C0C0C0A4F8C08099",
 27085 => x"C0C0C0A4F8C08092",
 27086 => x"C0C0C0A4F8C08082",
 27087 => x"C0C0C0A4F8C080F8",
 27088 => x"C0C0C0A4F8C08080",
 27089 => x"C0C0C0A4F8C08090",
 27090 => x"C0C0C0A4F8C090C0",
 27091 => x"C0C0C0A4F8C090F9",
 27092 => x"C0C0C0A4F8C090A4",
 27093 => x"C0C0C0A4F8C090B0",
 27094 => x"C0C0C0A4F8C09099",
 27095 => x"C0C0C0A4F8C09092",
 27096 => x"C0C0C0A4F8C09082",
 27097 => x"C0C0C0A4F8C090F8",
 27098 => x"C0C0C0A4F8C09080",
 27099 => x"C0C0C0A4F8C09090",
 27100 => x"C0C0C0A4F8F9C0C0",
 27101 => x"C0C0C0A4F8F9C0F9",
 27102 => x"C0C0C0A4F8F9C0A4",
 27103 => x"C0C0C0A4F8F9C0B0",
 27104 => x"C0C0C0A4F8F9C099",
 27105 => x"C0C0C0A4F8F9C092",
 27106 => x"C0C0C0A4F8F9C082",
 27107 => x"C0C0C0A4F8F9C0F8",
 27108 => x"C0C0C0A4F8F9C080",
 27109 => x"C0C0C0A4F8F9C090",
 27110 => x"C0C0C0A4F8F9F9C0",
 27111 => x"C0C0C0A4F8F9F9F9",
 27112 => x"C0C0C0A4F8F9F9A4",
 27113 => x"C0C0C0A4F8F9F9B0",
 27114 => x"C0C0C0A4F8F9F999",
 27115 => x"C0C0C0A4F8F9F992",
 27116 => x"C0C0C0A4F8F9F982",
 27117 => x"C0C0C0A4F8F9F9F8",
 27118 => x"C0C0C0A4F8F9F980",
 27119 => x"C0C0C0A4F8F9F990",
 27120 => x"C0C0C0A4F8F9A4C0",
 27121 => x"C0C0C0A4F8F9A4F9",
 27122 => x"C0C0C0A4F8F9A4A4",
 27123 => x"C0C0C0A4F8F9A4B0",
 27124 => x"C0C0C0A4F8F9A499",
 27125 => x"C0C0C0A4F8F9A492",
 27126 => x"C0C0C0A4F8F9A482",
 27127 => x"C0C0C0A4F8F9A4F8",
 27128 => x"C0C0C0A4F8F9A480",
 27129 => x"C0C0C0A4F8F9A490",
 27130 => x"C0C0C0A4F8F9B0C0",
 27131 => x"C0C0C0A4F8F9B0F9",
 27132 => x"C0C0C0A4F8F9B0A4",
 27133 => x"C0C0C0A4F8F9B0B0",
 27134 => x"C0C0C0A4F8F9B099",
 27135 => x"C0C0C0A4F8F9B092",
 27136 => x"C0C0C0A4F8F9B082",
 27137 => x"C0C0C0A4F8F9B0F8",
 27138 => x"C0C0C0A4F8F9B080",
 27139 => x"C0C0C0A4F8F9B090",
 27140 => x"C0C0C0A4F8F999C0",
 27141 => x"C0C0C0A4F8F999F9",
 27142 => x"C0C0C0A4F8F999A4",
 27143 => x"C0C0C0A4F8F999B0",
 27144 => x"C0C0C0A4F8F99999",
 27145 => x"C0C0C0A4F8F99992",
 27146 => x"C0C0C0A4F8F99982",
 27147 => x"C0C0C0A4F8F999F8",
 27148 => x"C0C0C0A4F8F99980",
 27149 => x"C0C0C0A4F8F99990",
 27150 => x"C0C0C0A4F8F992C0",
 27151 => x"C0C0C0A4F8F992F9",
 27152 => x"C0C0C0A4F8F992A4",
 27153 => x"C0C0C0A4F8F992B0",
 27154 => x"C0C0C0A4F8F99299",
 27155 => x"C0C0C0A4F8F99292",
 27156 => x"C0C0C0A4F8F99282",
 27157 => x"C0C0C0A4F8F992F8",
 27158 => x"C0C0C0A4F8F99280",
 27159 => x"C0C0C0A4F8F99290",
 27160 => x"C0C0C0A4F8F982C0",
 27161 => x"C0C0C0A4F8F982F9",
 27162 => x"C0C0C0A4F8F982A4",
 27163 => x"C0C0C0A4F8F982B0",
 27164 => x"C0C0C0A4F8F98299",
 27165 => x"C0C0C0A4F8F98292",
 27166 => x"C0C0C0A4F8F98282",
 27167 => x"C0C0C0A4F8F982F8",
 27168 => x"C0C0C0A4F8F98280",
 27169 => x"C0C0C0A4F8F98290",
 27170 => x"C0C0C0A4F8F9F8C0",
 27171 => x"C0C0C0A4F8F9F8F9",
 27172 => x"C0C0C0A4F8F9F8A4",
 27173 => x"C0C0C0A4F8F9F8B0",
 27174 => x"C0C0C0A4F8F9F899",
 27175 => x"C0C0C0A4F8F9F892",
 27176 => x"C0C0C0A4F8F9F882",
 27177 => x"C0C0C0A4F8F9F8F8",
 27178 => x"C0C0C0A4F8F9F880",
 27179 => x"C0C0C0A4F8F9F890",
 27180 => x"C0C0C0A4F8F980C0",
 27181 => x"C0C0C0A4F8F980F9",
 27182 => x"C0C0C0A4F8F980A4",
 27183 => x"C0C0C0A4F8F980B0",
 27184 => x"C0C0C0A4F8F98099",
 27185 => x"C0C0C0A4F8F98092",
 27186 => x"C0C0C0A4F8F98082",
 27187 => x"C0C0C0A4F8F980F8",
 27188 => x"C0C0C0A4F8F98080",
 27189 => x"C0C0C0A4F8F98090",
 27190 => x"C0C0C0A4F8F990C0",
 27191 => x"C0C0C0A4F8F990F9",
 27192 => x"C0C0C0A4F8F990A4",
 27193 => x"C0C0C0A4F8F990B0",
 27194 => x"C0C0C0A4F8F99099",
 27195 => x"C0C0C0A4F8F99092",
 27196 => x"C0C0C0A4F8F99082",
 27197 => x"C0C0C0A4F8F990F8",
 27198 => x"C0C0C0A4F8F99080",
 27199 => x"C0C0C0A4F8F99090",
 27200 => x"C0C0C0A4F8A4C0C0",
 27201 => x"C0C0C0A4F8A4C0F9",
 27202 => x"C0C0C0A4F8A4C0A4",
 27203 => x"C0C0C0A4F8A4C0B0",
 27204 => x"C0C0C0A4F8A4C099",
 27205 => x"C0C0C0A4F8A4C092",
 27206 => x"C0C0C0A4F8A4C082",
 27207 => x"C0C0C0A4F8A4C0F8",
 27208 => x"C0C0C0A4F8A4C080",
 27209 => x"C0C0C0A4F8A4C090",
 27210 => x"C0C0C0A4F8A4F9C0",
 27211 => x"C0C0C0A4F8A4F9F9",
 27212 => x"C0C0C0A4F8A4F9A4",
 27213 => x"C0C0C0A4F8A4F9B0",
 27214 => x"C0C0C0A4F8A4F999",
 27215 => x"C0C0C0A4F8A4F992",
 27216 => x"C0C0C0A4F8A4F982",
 27217 => x"C0C0C0A4F8A4F9F8",
 27218 => x"C0C0C0A4F8A4F980",
 27219 => x"C0C0C0A4F8A4F990",
 27220 => x"C0C0C0A4F8A4A4C0",
 27221 => x"C0C0C0A4F8A4A4F9",
 27222 => x"C0C0C0A4F8A4A4A4",
 27223 => x"C0C0C0A4F8A4A4B0",
 27224 => x"C0C0C0A4F8A4A499",
 27225 => x"C0C0C0A4F8A4A492",
 27226 => x"C0C0C0A4F8A4A482",
 27227 => x"C0C0C0A4F8A4A4F8",
 27228 => x"C0C0C0A4F8A4A480",
 27229 => x"C0C0C0A4F8A4A490",
 27230 => x"C0C0C0A4F8A4B0C0",
 27231 => x"C0C0C0A4F8A4B0F9",
 27232 => x"C0C0C0A4F8A4B0A4",
 27233 => x"C0C0C0A4F8A4B0B0",
 27234 => x"C0C0C0A4F8A4B099",
 27235 => x"C0C0C0A4F8A4B092",
 27236 => x"C0C0C0A4F8A4B082",
 27237 => x"C0C0C0A4F8A4B0F8",
 27238 => x"C0C0C0A4F8A4B080",
 27239 => x"C0C0C0A4F8A4B090",
 27240 => x"C0C0C0A4F8A499C0",
 27241 => x"C0C0C0A4F8A499F9",
 27242 => x"C0C0C0A4F8A499A4",
 27243 => x"C0C0C0A4F8A499B0",
 27244 => x"C0C0C0A4F8A49999",
 27245 => x"C0C0C0A4F8A49992",
 27246 => x"C0C0C0A4F8A49982",
 27247 => x"C0C0C0A4F8A499F8",
 27248 => x"C0C0C0A4F8A49980",
 27249 => x"C0C0C0A4F8A49990",
 27250 => x"C0C0C0A4F8A492C0",
 27251 => x"C0C0C0A4F8A492F9",
 27252 => x"C0C0C0A4F8A492A4",
 27253 => x"C0C0C0A4F8A492B0",
 27254 => x"C0C0C0A4F8A49299",
 27255 => x"C0C0C0A4F8A49292",
 27256 => x"C0C0C0A4F8A49282",
 27257 => x"C0C0C0A4F8A492F8",
 27258 => x"C0C0C0A4F8A49280",
 27259 => x"C0C0C0A4F8A49290",
 27260 => x"C0C0C0A4F8A482C0",
 27261 => x"C0C0C0A4F8A482F9",
 27262 => x"C0C0C0A4F8A482A4",
 27263 => x"C0C0C0A4F8A482B0",
 27264 => x"C0C0C0A4F8A48299",
 27265 => x"C0C0C0A4F8A48292",
 27266 => x"C0C0C0A4F8A48282",
 27267 => x"C0C0C0A4F8A482F8",
 27268 => x"C0C0C0A4F8A48280",
 27269 => x"C0C0C0A4F8A48290",
 27270 => x"C0C0C0A4F8A4F8C0",
 27271 => x"C0C0C0A4F8A4F8F9",
 27272 => x"C0C0C0A4F8A4F8A4",
 27273 => x"C0C0C0A4F8A4F8B0",
 27274 => x"C0C0C0A4F8A4F899",
 27275 => x"C0C0C0A4F8A4F892",
 27276 => x"C0C0C0A4F8A4F882",
 27277 => x"C0C0C0A4F8A4F8F8",
 27278 => x"C0C0C0A4F8A4F880",
 27279 => x"C0C0C0A4F8A4F890",
 27280 => x"C0C0C0A4F8A480C0",
 27281 => x"C0C0C0A4F8A480F9",
 27282 => x"C0C0C0A4F8A480A4",
 27283 => x"C0C0C0A4F8A480B0",
 27284 => x"C0C0C0A4F8A48099",
 27285 => x"C0C0C0A4F8A48092",
 27286 => x"C0C0C0A4F8A48082",
 27287 => x"C0C0C0A4F8A480F8",
 27288 => x"C0C0C0A4F8A48080",
 27289 => x"C0C0C0A4F8A48090",
 27290 => x"C0C0C0A4F8A490C0",
 27291 => x"C0C0C0A4F8A490F9",
 27292 => x"C0C0C0A4F8A490A4",
 27293 => x"C0C0C0A4F8A490B0",
 27294 => x"C0C0C0A4F8A49099",
 27295 => x"C0C0C0A4F8A49092",
 27296 => x"C0C0C0A4F8A49082",
 27297 => x"C0C0C0A4F8A490F8",
 27298 => x"C0C0C0A4F8A49080",
 27299 => x"C0C0C0A4F8A49090",
 27300 => x"C0C0C0A4F8B0C0C0",
 27301 => x"C0C0C0A4F8B0C0F9",
 27302 => x"C0C0C0A4F8B0C0A4",
 27303 => x"C0C0C0A4F8B0C0B0",
 27304 => x"C0C0C0A4F8B0C099",
 27305 => x"C0C0C0A4F8B0C092",
 27306 => x"C0C0C0A4F8B0C082",
 27307 => x"C0C0C0A4F8B0C0F8",
 27308 => x"C0C0C0A4F8B0C080",
 27309 => x"C0C0C0A4F8B0C090",
 27310 => x"C0C0C0A4F8B0F9C0",
 27311 => x"C0C0C0A4F8B0F9F9",
 27312 => x"C0C0C0A4F8B0F9A4",
 27313 => x"C0C0C0A4F8B0F9B0",
 27314 => x"C0C0C0A4F8B0F999",
 27315 => x"C0C0C0A4F8B0F992",
 27316 => x"C0C0C0A4F8B0F982",
 27317 => x"C0C0C0A4F8B0F9F8",
 27318 => x"C0C0C0A4F8B0F980",
 27319 => x"C0C0C0A4F8B0F990",
 27320 => x"C0C0C0A4F8B0A4C0",
 27321 => x"C0C0C0A4F8B0A4F9",
 27322 => x"C0C0C0A4F8B0A4A4",
 27323 => x"C0C0C0A4F8B0A4B0",
 27324 => x"C0C0C0A4F8B0A499",
 27325 => x"C0C0C0A4F8B0A492",
 27326 => x"C0C0C0A4F8B0A482",
 27327 => x"C0C0C0A4F8B0A4F8",
 27328 => x"C0C0C0A4F8B0A480",
 27329 => x"C0C0C0A4F8B0A490",
 27330 => x"C0C0C0A4F8B0B0C0",
 27331 => x"C0C0C0A4F8B0B0F9",
 27332 => x"C0C0C0A4F8B0B0A4",
 27333 => x"C0C0C0A4F8B0B0B0",
 27334 => x"C0C0C0A4F8B0B099",
 27335 => x"C0C0C0A4F8B0B092",
 27336 => x"C0C0C0A4F8B0B082",
 27337 => x"C0C0C0A4F8B0B0F8",
 27338 => x"C0C0C0A4F8B0B080",
 27339 => x"C0C0C0A4F8B0B090",
 27340 => x"C0C0C0A4F8B099C0",
 27341 => x"C0C0C0A4F8B099F9",
 27342 => x"C0C0C0A4F8B099A4",
 27343 => x"C0C0C0A4F8B099B0",
 27344 => x"C0C0C0A4F8B09999",
 27345 => x"C0C0C0A4F8B09992",
 27346 => x"C0C0C0A4F8B09982",
 27347 => x"C0C0C0A4F8B099F8",
 27348 => x"C0C0C0A4F8B09980",
 27349 => x"C0C0C0A4F8B09990",
 27350 => x"C0C0C0A4F8B092C0",
 27351 => x"C0C0C0A4F8B092F9",
 27352 => x"C0C0C0A4F8B092A4",
 27353 => x"C0C0C0A4F8B092B0",
 27354 => x"C0C0C0A4F8B09299",
 27355 => x"C0C0C0A4F8B09292",
 27356 => x"C0C0C0A4F8B09282",
 27357 => x"C0C0C0A4F8B092F8",
 27358 => x"C0C0C0A4F8B09280",
 27359 => x"C0C0C0A4F8B09290",
 27360 => x"C0C0C0A4F8B082C0",
 27361 => x"C0C0C0A4F8B082F9",
 27362 => x"C0C0C0A4F8B082A4",
 27363 => x"C0C0C0A4F8B082B0",
 27364 => x"C0C0C0A4F8B08299",
 27365 => x"C0C0C0A4F8B08292",
 27366 => x"C0C0C0A4F8B08282",
 27367 => x"C0C0C0A4F8B082F8",
 27368 => x"C0C0C0A4F8B08280",
 27369 => x"C0C0C0A4F8B08290",
 27370 => x"C0C0C0A4F8B0F8C0",
 27371 => x"C0C0C0A4F8B0F8F9",
 27372 => x"C0C0C0A4F8B0F8A4",
 27373 => x"C0C0C0A4F8B0F8B0",
 27374 => x"C0C0C0A4F8B0F899",
 27375 => x"C0C0C0A4F8B0F892",
 27376 => x"C0C0C0A4F8B0F882",
 27377 => x"C0C0C0A4F8B0F8F8",
 27378 => x"C0C0C0A4F8B0F880",
 27379 => x"C0C0C0A4F8B0F890",
 27380 => x"C0C0C0A4F8B080C0",
 27381 => x"C0C0C0A4F8B080F9",
 27382 => x"C0C0C0A4F8B080A4",
 27383 => x"C0C0C0A4F8B080B0",
 27384 => x"C0C0C0A4F8B08099",
 27385 => x"C0C0C0A4F8B08092",
 27386 => x"C0C0C0A4F8B08082",
 27387 => x"C0C0C0A4F8B080F8",
 27388 => x"C0C0C0A4F8B08080",
 27389 => x"C0C0C0A4F8B08090",
 27390 => x"C0C0C0A4F8B090C0",
 27391 => x"C0C0C0A4F8B090F9",
 27392 => x"C0C0C0A4F8B090A4",
 27393 => x"C0C0C0A4F8B090B0",
 27394 => x"C0C0C0A4F8B09099",
 27395 => x"C0C0C0A4F8B09092",
 27396 => x"C0C0C0A4F8B09082",
 27397 => x"C0C0C0A4F8B090F8",
 27398 => x"C0C0C0A4F8B09080",
 27399 => x"C0C0C0A4F8B09090",
 27400 => x"C0C0C0A4F899C0C0",
 27401 => x"C0C0C0A4F899C0F9",
 27402 => x"C0C0C0A4F899C0A4",
 27403 => x"C0C0C0A4F899C0B0",
 27404 => x"C0C0C0A4F899C099",
 27405 => x"C0C0C0A4F899C092",
 27406 => x"C0C0C0A4F899C082",
 27407 => x"C0C0C0A4F899C0F8",
 27408 => x"C0C0C0A4F899C080",
 27409 => x"C0C0C0A4F899C090",
 27410 => x"C0C0C0A4F899F9C0",
 27411 => x"C0C0C0A4F899F9F9",
 27412 => x"C0C0C0A4F899F9A4",
 27413 => x"C0C0C0A4F899F9B0",
 27414 => x"C0C0C0A4F899F999",
 27415 => x"C0C0C0A4F899F992",
 27416 => x"C0C0C0A4F899F982",
 27417 => x"C0C0C0A4F899F9F8",
 27418 => x"C0C0C0A4F899F980",
 27419 => x"C0C0C0A4F899F990",
 27420 => x"C0C0C0A4F899A4C0",
 27421 => x"C0C0C0A4F899A4F9",
 27422 => x"C0C0C0A4F899A4A4",
 27423 => x"C0C0C0A4F899A4B0",
 27424 => x"C0C0C0A4F899A499",
 27425 => x"C0C0C0A4F899A492",
 27426 => x"C0C0C0A4F899A482",
 27427 => x"C0C0C0A4F899A4F8",
 27428 => x"C0C0C0A4F899A480",
 27429 => x"C0C0C0A4F899A490",
 27430 => x"C0C0C0A4F899B0C0",
 27431 => x"C0C0C0A4F899B0F9",
 27432 => x"C0C0C0A4F899B0A4",
 27433 => x"C0C0C0A4F899B0B0",
 27434 => x"C0C0C0A4F899B099",
 27435 => x"C0C0C0A4F899B092",
 27436 => x"C0C0C0A4F899B082",
 27437 => x"C0C0C0A4F899B0F8",
 27438 => x"C0C0C0A4F899B080",
 27439 => x"C0C0C0A4F899B090",
 27440 => x"C0C0C0A4F89999C0",
 27441 => x"C0C0C0A4F89999F9",
 27442 => x"C0C0C0A4F89999A4",
 27443 => x"C0C0C0A4F89999B0",
 27444 => x"C0C0C0A4F8999999",
 27445 => x"C0C0C0A4F8999992",
 27446 => x"C0C0C0A4F8999982",
 27447 => x"C0C0C0A4F89999F8",
 27448 => x"C0C0C0A4F8999980",
 27449 => x"C0C0C0A4F8999990",
 27450 => x"C0C0C0A4F89992C0",
 27451 => x"C0C0C0A4F89992F9",
 27452 => x"C0C0C0A4F89992A4",
 27453 => x"C0C0C0A4F89992B0",
 27454 => x"C0C0C0A4F8999299",
 27455 => x"C0C0C0A4F8999292",
 27456 => x"C0C0C0A4F8999282",
 27457 => x"C0C0C0A4F89992F8",
 27458 => x"C0C0C0A4F8999280",
 27459 => x"C0C0C0A4F8999290",
 27460 => x"C0C0C0A4F89982C0",
 27461 => x"C0C0C0A4F89982F9",
 27462 => x"C0C0C0A4F89982A4",
 27463 => x"C0C0C0A4F89982B0",
 27464 => x"C0C0C0A4F8998299",
 27465 => x"C0C0C0A4F8998292",
 27466 => x"C0C0C0A4F8998282",
 27467 => x"C0C0C0A4F89982F8",
 27468 => x"C0C0C0A4F8998280",
 27469 => x"C0C0C0A4F8998290",
 27470 => x"C0C0C0A4F899F8C0",
 27471 => x"C0C0C0A4F899F8F9",
 27472 => x"C0C0C0A4F899F8A4",
 27473 => x"C0C0C0A4F899F8B0",
 27474 => x"C0C0C0A4F899F899",
 27475 => x"C0C0C0A4F899F892",
 27476 => x"C0C0C0A4F899F882",
 27477 => x"C0C0C0A4F899F8F8",
 27478 => x"C0C0C0A4F899F880",
 27479 => x"C0C0C0A4F899F890",
 27480 => x"C0C0C0A4F89980C0",
 27481 => x"C0C0C0A4F89980F9",
 27482 => x"C0C0C0A4F89980A4",
 27483 => x"C0C0C0A4F89980B0",
 27484 => x"C0C0C0A4F8998099",
 27485 => x"C0C0C0A4F8998092",
 27486 => x"C0C0C0A4F8998082",
 27487 => x"C0C0C0A4F89980F8",
 27488 => x"C0C0C0A4F8998080",
 27489 => x"C0C0C0A4F8998090",
 27490 => x"C0C0C0A4F89990C0",
 27491 => x"C0C0C0A4F89990F9",
 27492 => x"C0C0C0A4F89990A4",
 27493 => x"C0C0C0A4F89990B0",
 27494 => x"C0C0C0A4F8999099",
 27495 => x"C0C0C0A4F8999092",
 27496 => x"C0C0C0A4F8999082",
 27497 => x"C0C0C0A4F89990F8",
 27498 => x"C0C0C0A4F8999080",
 27499 => x"C0C0C0A4F8999090",
 27500 => x"C0C0C0A4F892C0C0",
 27501 => x"C0C0C0A4F892C0F9",
 27502 => x"C0C0C0A4F892C0A4",
 27503 => x"C0C0C0A4F892C0B0",
 27504 => x"C0C0C0A4F892C099",
 27505 => x"C0C0C0A4F892C092",
 27506 => x"C0C0C0A4F892C082",
 27507 => x"C0C0C0A4F892C0F8",
 27508 => x"C0C0C0A4F892C080",
 27509 => x"C0C0C0A4F892C090",
 27510 => x"C0C0C0A4F892F9C0",
 27511 => x"C0C0C0A4F892F9F9",
 27512 => x"C0C0C0A4F892F9A4",
 27513 => x"C0C0C0A4F892F9B0",
 27514 => x"C0C0C0A4F892F999",
 27515 => x"C0C0C0A4F892F992",
 27516 => x"C0C0C0A4F892F982",
 27517 => x"C0C0C0A4F892F9F8",
 27518 => x"C0C0C0A4F892F980",
 27519 => x"C0C0C0A4F892F990",
 27520 => x"C0C0C0A4F892A4C0",
 27521 => x"C0C0C0A4F892A4F9",
 27522 => x"C0C0C0A4F892A4A4",
 27523 => x"C0C0C0A4F892A4B0",
 27524 => x"C0C0C0A4F892A499",
 27525 => x"C0C0C0A4F892A492",
 27526 => x"C0C0C0A4F892A482",
 27527 => x"C0C0C0A4F892A4F8",
 27528 => x"C0C0C0A4F892A480",
 27529 => x"C0C0C0A4F892A490",
 27530 => x"C0C0C0A4F892B0C0",
 27531 => x"C0C0C0A4F892B0F9",
 27532 => x"C0C0C0A4F892B0A4",
 27533 => x"C0C0C0A4F892B0B0",
 27534 => x"C0C0C0A4F892B099",
 27535 => x"C0C0C0A4F892B092",
 27536 => x"C0C0C0A4F892B082",
 27537 => x"C0C0C0A4F892B0F8",
 27538 => x"C0C0C0A4F892B080",
 27539 => x"C0C0C0A4F892B090",
 27540 => x"C0C0C0A4F89299C0",
 27541 => x"C0C0C0A4F89299F9",
 27542 => x"C0C0C0A4F89299A4",
 27543 => x"C0C0C0A4F89299B0",
 27544 => x"C0C0C0A4F8929999",
 27545 => x"C0C0C0A4F8929992",
 27546 => x"C0C0C0A4F8929982",
 27547 => x"C0C0C0A4F89299F8",
 27548 => x"C0C0C0A4F8929980",
 27549 => x"C0C0C0A4F8929990",
 27550 => x"C0C0C0A4F89292C0",
 27551 => x"C0C0C0A4F89292F9",
 27552 => x"C0C0C0A4F89292A4",
 27553 => x"C0C0C0A4F89292B0",
 27554 => x"C0C0C0A4F8929299",
 27555 => x"C0C0C0A4F8929292",
 27556 => x"C0C0C0A4F8929282",
 27557 => x"C0C0C0A4F89292F8",
 27558 => x"C0C0C0A4F8929280",
 27559 => x"C0C0C0A4F8929290",
 27560 => x"C0C0C0A4F89282C0",
 27561 => x"C0C0C0A4F89282F9",
 27562 => x"C0C0C0A4F89282A4",
 27563 => x"C0C0C0A4F89282B0",
 27564 => x"C0C0C0A4F8928299",
 27565 => x"C0C0C0A4F8928292",
 27566 => x"C0C0C0A4F8928282",
 27567 => x"C0C0C0A4F89282F8",
 27568 => x"C0C0C0A4F8928280",
 27569 => x"C0C0C0A4F8928290",
 27570 => x"C0C0C0A4F892F8C0",
 27571 => x"C0C0C0A4F892F8F9",
 27572 => x"C0C0C0A4F892F8A4",
 27573 => x"C0C0C0A4F892F8B0",
 27574 => x"C0C0C0A4F892F899",
 27575 => x"C0C0C0A4F892F892",
 27576 => x"C0C0C0A4F892F882",
 27577 => x"C0C0C0A4F892F8F8",
 27578 => x"C0C0C0A4F892F880",
 27579 => x"C0C0C0A4F892F890",
 27580 => x"C0C0C0A4F89280C0",
 27581 => x"C0C0C0A4F89280F9",
 27582 => x"C0C0C0A4F89280A4",
 27583 => x"C0C0C0A4F89280B0",
 27584 => x"C0C0C0A4F8928099",
 27585 => x"C0C0C0A4F8928092",
 27586 => x"C0C0C0A4F8928082",
 27587 => x"C0C0C0A4F89280F8",
 27588 => x"C0C0C0A4F8928080",
 27589 => x"C0C0C0A4F8928090",
 27590 => x"C0C0C0A4F89290C0",
 27591 => x"C0C0C0A4F89290F9",
 27592 => x"C0C0C0A4F89290A4",
 27593 => x"C0C0C0A4F89290B0",
 27594 => x"C0C0C0A4F8929099",
 27595 => x"C0C0C0A4F8929092",
 27596 => x"C0C0C0A4F8929082",
 27597 => x"C0C0C0A4F89290F8",
 27598 => x"C0C0C0A4F8929080",
 27599 => x"C0C0C0A4F8929090",
 27600 => x"C0C0C0A4F882C0C0",
 27601 => x"C0C0C0A4F882C0F9",
 27602 => x"C0C0C0A4F882C0A4",
 27603 => x"C0C0C0A4F882C0B0",
 27604 => x"C0C0C0A4F882C099",
 27605 => x"C0C0C0A4F882C092",
 27606 => x"C0C0C0A4F882C082",
 27607 => x"C0C0C0A4F882C0F8",
 27608 => x"C0C0C0A4F882C080",
 27609 => x"C0C0C0A4F882C090",
 27610 => x"C0C0C0A4F882F9C0",
 27611 => x"C0C0C0A4F882F9F9",
 27612 => x"C0C0C0A4F882F9A4",
 27613 => x"C0C0C0A4F882F9B0",
 27614 => x"C0C0C0A4F882F999",
 27615 => x"C0C0C0A4F882F992",
 27616 => x"C0C0C0A4F882F982",
 27617 => x"C0C0C0A4F882F9F8",
 27618 => x"C0C0C0A4F882F980",
 27619 => x"C0C0C0A4F882F990",
 27620 => x"C0C0C0A4F882A4C0",
 27621 => x"C0C0C0A4F882A4F9",
 27622 => x"C0C0C0A4F882A4A4",
 27623 => x"C0C0C0A4F882A4B0",
 27624 => x"C0C0C0A4F882A499",
 27625 => x"C0C0C0A4F882A492",
 27626 => x"C0C0C0A4F882A482",
 27627 => x"C0C0C0A4F882A4F8",
 27628 => x"C0C0C0A4F882A480",
 27629 => x"C0C0C0A4F882A490",
 27630 => x"C0C0C0A4F882B0C0",
 27631 => x"C0C0C0A4F882B0F9",
 27632 => x"C0C0C0A4F882B0A4",
 27633 => x"C0C0C0A4F882B0B0",
 27634 => x"C0C0C0A4F882B099",
 27635 => x"C0C0C0A4F882B092",
 27636 => x"C0C0C0A4F882B082",
 27637 => x"C0C0C0A4F882B0F8",
 27638 => x"C0C0C0A4F882B080",
 27639 => x"C0C0C0A4F882B090",
 27640 => x"C0C0C0A4F88299C0",
 27641 => x"C0C0C0A4F88299F9",
 27642 => x"C0C0C0A4F88299A4",
 27643 => x"C0C0C0A4F88299B0",
 27644 => x"C0C0C0A4F8829999",
 27645 => x"C0C0C0A4F8829992",
 27646 => x"C0C0C0A4F8829982",
 27647 => x"C0C0C0A4F88299F8",
 27648 => x"C0C0C0A4F8829980",
 27649 => x"C0C0C0A4F8829990",
 27650 => x"C0C0C0A4F88292C0",
 27651 => x"C0C0C0A4F88292F9",
 27652 => x"C0C0C0A4F88292A4",
 27653 => x"C0C0C0A4F88292B0",
 27654 => x"C0C0C0A4F8829299",
 27655 => x"C0C0C0A4F8829292",
 27656 => x"C0C0C0A4F8829282",
 27657 => x"C0C0C0A4F88292F8",
 27658 => x"C0C0C0A4F8829280",
 27659 => x"C0C0C0A4F8829290",
 27660 => x"C0C0C0A4F88282C0",
 27661 => x"C0C0C0A4F88282F9",
 27662 => x"C0C0C0A4F88282A4",
 27663 => x"C0C0C0A4F88282B0",
 27664 => x"C0C0C0A4F8828299",
 27665 => x"C0C0C0A4F8828292",
 27666 => x"C0C0C0A4F8828282",
 27667 => x"C0C0C0A4F88282F8",
 27668 => x"C0C0C0A4F8828280",
 27669 => x"C0C0C0A4F8828290",
 27670 => x"C0C0C0A4F882F8C0",
 27671 => x"C0C0C0A4F882F8F9",
 27672 => x"C0C0C0A4F882F8A4",
 27673 => x"C0C0C0A4F882F8B0",
 27674 => x"C0C0C0A4F882F899",
 27675 => x"C0C0C0A4F882F892",
 27676 => x"C0C0C0A4F882F882",
 27677 => x"C0C0C0A4F882F8F8",
 27678 => x"C0C0C0A4F882F880",
 27679 => x"C0C0C0A4F882F890",
 27680 => x"C0C0C0A4F88280C0",
 27681 => x"C0C0C0A4F88280F9",
 27682 => x"C0C0C0A4F88280A4",
 27683 => x"C0C0C0A4F88280B0",
 27684 => x"C0C0C0A4F8828099",
 27685 => x"C0C0C0A4F8828092",
 27686 => x"C0C0C0A4F8828082",
 27687 => x"C0C0C0A4F88280F8",
 27688 => x"C0C0C0A4F8828080",
 27689 => x"C0C0C0A4F8828090",
 27690 => x"C0C0C0A4F88290C0",
 27691 => x"C0C0C0A4F88290F9",
 27692 => x"C0C0C0A4F88290A4",
 27693 => x"C0C0C0A4F88290B0",
 27694 => x"C0C0C0A4F8829099",
 27695 => x"C0C0C0A4F8829092",
 27696 => x"C0C0C0A4F8829082",
 27697 => x"C0C0C0A4F88290F8",
 27698 => x"C0C0C0A4F8829080",
 27699 => x"C0C0C0A4F8829090",
 27700 => x"C0C0C0A4F8F8C0C0",
 27701 => x"C0C0C0A4F8F8C0F9",
 27702 => x"C0C0C0A4F8F8C0A4",
 27703 => x"C0C0C0A4F8F8C0B0",
 27704 => x"C0C0C0A4F8F8C099",
 27705 => x"C0C0C0A4F8F8C092",
 27706 => x"C0C0C0A4F8F8C082",
 27707 => x"C0C0C0A4F8F8C0F8",
 27708 => x"C0C0C0A4F8F8C080",
 27709 => x"C0C0C0A4F8F8C090",
 27710 => x"C0C0C0A4F8F8F9C0",
 27711 => x"C0C0C0A4F8F8F9F9",
 27712 => x"C0C0C0A4F8F8F9A4",
 27713 => x"C0C0C0A4F8F8F9B0",
 27714 => x"C0C0C0A4F8F8F999",
 27715 => x"C0C0C0A4F8F8F992",
 27716 => x"C0C0C0A4F8F8F982",
 27717 => x"C0C0C0A4F8F8F9F8",
 27718 => x"C0C0C0A4F8F8F980",
 27719 => x"C0C0C0A4F8F8F990",
 27720 => x"C0C0C0A4F8F8A4C0",
 27721 => x"C0C0C0A4F8F8A4F9",
 27722 => x"C0C0C0A4F8F8A4A4",
 27723 => x"C0C0C0A4F8F8A4B0",
 27724 => x"C0C0C0A4F8F8A499",
 27725 => x"C0C0C0A4F8F8A492",
 27726 => x"C0C0C0A4F8F8A482",
 27727 => x"C0C0C0A4F8F8A4F8",
 27728 => x"C0C0C0A4F8F8A480",
 27729 => x"C0C0C0A4F8F8A490",
 27730 => x"C0C0C0A4F8F8B0C0",
 27731 => x"C0C0C0A4F8F8B0F9",
 27732 => x"C0C0C0A4F8F8B0A4",
 27733 => x"C0C0C0A4F8F8B0B0",
 27734 => x"C0C0C0A4F8F8B099",
 27735 => x"C0C0C0A4F8F8B092",
 27736 => x"C0C0C0A4F8F8B082",
 27737 => x"C0C0C0A4F8F8B0F8",
 27738 => x"C0C0C0A4F8F8B080",
 27739 => x"C0C0C0A4F8F8B090",
 27740 => x"C0C0C0A4F8F899C0",
 27741 => x"C0C0C0A4F8F899F9",
 27742 => x"C0C0C0A4F8F899A4",
 27743 => x"C0C0C0A4F8F899B0",
 27744 => x"C0C0C0A4F8F89999",
 27745 => x"C0C0C0A4F8F89992",
 27746 => x"C0C0C0A4F8F89982",
 27747 => x"C0C0C0A4F8F899F8",
 27748 => x"C0C0C0A4F8F89980",
 27749 => x"C0C0C0A4F8F89990",
 27750 => x"C0C0C0A4F8F892C0",
 27751 => x"C0C0C0A4F8F892F9",
 27752 => x"C0C0C0A4F8F892A4",
 27753 => x"C0C0C0A4F8F892B0",
 27754 => x"C0C0C0A4F8F89299",
 27755 => x"C0C0C0A4F8F89292",
 27756 => x"C0C0C0A4F8F89282",
 27757 => x"C0C0C0A4F8F892F8",
 27758 => x"C0C0C0A4F8F89280",
 27759 => x"C0C0C0A4F8F89290",
 27760 => x"C0C0C0A4F8F882C0",
 27761 => x"C0C0C0A4F8F882F9",
 27762 => x"C0C0C0A4F8F882A4",
 27763 => x"C0C0C0A4F8F882B0",
 27764 => x"C0C0C0A4F8F88299",
 27765 => x"C0C0C0A4F8F88292",
 27766 => x"C0C0C0A4F8F88282",
 27767 => x"C0C0C0A4F8F882F8",
 27768 => x"C0C0C0A4F8F88280",
 27769 => x"C0C0C0A4F8F88290",
 27770 => x"C0C0C0A4F8F8F8C0",
 27771 => x"C0C0C0A4F8F8F8F9",
 27772 => x"C0C0C0A4F8F8F8A4",
 27773 => x"C0C0C0A4F8F8F8B0",
 27774 => x"C0C0C0A4F8F8F899",
 27775 => x"C0C0C0A4F8F8F892",
 27776 => x"C0C0C0A4F8F8F882",
 27777 => x"C0C0C0A4F8F8F8F8",
 27778 => x"C0C0C0A4F8F8F880",
 27779 => x"C0C0C0A4F8F8F890",
 27780 => x"C0C0C0A4F8F880C0",
 27781 => x"C0C0C0A4F8F880F9",
 27782 => x"C0C0C0A4F8F880A4",
 27783 => x"C0C0C0A4F8F880B0",
 27784 => x"C0C0C0A4F8F88099",
 27785 => x"C0C0C0A4F8F88092",
 27786 => x"C0C0C0A4F8F88082",
 27787 => x"C0C0C0A4F8F880F8",
 27788 => x"C0C0C0A4F8F88080",
 27789 => x"C0C0C0A4F8F88090",
 27790 => x"C0C0C0A4F8F890C0",
 27791 => x"C0C0C0A4F8F890F9",
 27792 => x"C0C0C0A4F8F890A4",
 27793 => x"C0C0C0A4F8F890B0",
 27794 => x"C0C0C0A4F8F89099",
 27795 => x"C0C0C0A4F8F89092",
 27796 => x"C0C0C0A4F8F89082",
 27797 => x"C0C0C0A4F8F890F8",
 27798 => x"C0C0C0A4F8F89080",
 27799 => x"C0C0C0A4F8F89090",
 27800 => x"C0C0C0A4F880C0C0",
 27801 => x"C0C0C0A4F880C0F9",
 27802 => x"C0C0C0A4F880C0A4",
 27803 => x"C0C0C0A4F880C0B0",
 27804 => x"C0C0C0A4F880C099",
 27805 => x"C0C0C0A4F880C092",
 27806 => x"C0C0C0A4F880C082",
 27807 => x"C0C0C0A4F880C0F8",
 27808 => x"C0C0C0A4F880C080",
 27809 => x"C0C0C0A4F880C090",
 27810 => x"C0C0C0A4F880F9C0",
 27811 => x"C0C0C0A4F880F9F9",
 27812 => x"C0C0C0A4F880F9A4",
 27813 => x"C0C0C0A4F880F9B0",
 27814 => x"C0C0C0A4F880F999",
 27815 => x"C0C0C0A4F880F992",
 27816 => x"C0C0C0A4F880F982",
 27817 => x"C0C0C0A4F880F9F8",
 27818 => x"C0C0C0A4F880F980",
 27819 => x"C0C0C0A4F880F990",
 27820 => x"C0C0C0A4F880A4C0",
 27821 => x"C0C0C0A4F880A4F9",
 27822 => x"C0C0C0A4F880A4A4",
 27823 => x"C0C0C0A4F880A4B0",
 27824 => x"C0C0C0A4F880A499",
 27825 => x"C0C0C0A4F880A492",
 27826 => x"C0C0C0A4F880A482",
 27827 => x"C0C0C0A4F880A4F8",
 27828 => x"C0C0C0A4F880A480",
 27829 => x"C0C0C0A4F880A490",
 27830 => x"C0C0C0A4F880B0C0",
 27831 => x"C0C0C0A4F880B0F9",
 27832 => x"C0C0C0A4F880B0A4",
 27833 => x"C0C0C0A4F880B0B0",
 27834 => x"C0C0C0A4F880B099",
 27835 => x"C0C0C0A4F880B092",
 27836 => x"C0C0C0A4F880B082",
 27837 => x"C0C0C0A4F880B0F8",
 27838 => x"C0C0C0A4F880B080",
 27839 => x"C0C0C0A4F880B090",
 27840 => x"C0C0C0A4F88099C0",
 27841 => x"C0C0C0A4F88099F9",
 27842 => x"C0C0C0A4F88099A4",
 27843 => x"C0C0C0A4F88099B0",
 27844 => x"C0C0C0A4F8809999",
 27845 => x"C0C0C0A4F8809992",
 27846 => x"C0C0C0A4F8809982",
 27847 => x"C0C0C0A4F88099F8",
 27848 => x"C0C0C0A4F8809980",
 27849 => x"C0C0C0A4F8809990",
 27850 => x"C0C0C0A4F88092C0",
 27851 => x"C0C0C0A4F88092F9",
 27852 => x"C0C0C0A4F88092A4",
 27853 => x"C0C0C0A4F88092B0",
 27854 => x"C0C0C0A4F8809299",
 27855 => x"C0C0C0A4F8809292",
 27856 => x"C0C0C0A4F8809282",
 27857 => x"C0C0C0A4F88092F8",
 27858 => x"C0C0C0A4F8809280",
 27859 => x"C0C0C0A4F8809290",
 27860 => x"C0C0C0A4F88082C0",
 27861 => x"C0C0C0A4F88082F9",
 27862 => x"C0C0C0A4F88082A4",
 27863 => x"C0C0C0A4F88082B0",
 27864 => x"C0C0C0A4F8808299",
 27865 => x"C0C0C0A4F8808292",
 27866 => x"C0C0C0A4F8808282",
 27867 => x"C0C0C0A4F88082F8",
 27868 => x"C0C0C0A4F8808280",
 27869 => x"C0C0C0A4F8808290",
 27870 => x"C0C0C0A4F880F8C0",
 27871 => x"C0C0C0A4F880F8F9",
 27872 => x"C0C0C0A4F880F8A4",
 27873 => x"C0C0C0A4F880F8B0",
 27874 => x"C0C0C0A4F880F899",
 27875 => x"C0C0C0A4F880F892",
 27876 => x"C0C0C0A4F880F882",
 27877 => x"C0C0C0A4F880F8F8",
 27878 => x"C0C0C0A4F880F880",
 27879 => x"C0C0C0A4F880F890",
 27880 => x"C0C0C0A4F88080C0",
 27881 => x"C0C0C0A4F88080F9",
 27882 => x"C0C0C0A4F88080A4",
 27883 => x"C0C0C0A4F88080B0",
 27884 => x"C0C0C0A4F8808099",
 27885 => x"C0C0C0A4F8808092",
 27886 => x"C0C0C0A4F8808082",
 27887 => x"C0C0C0A4F88080F8",
 27888 => x"C0C0C0A4F8808080",
 27889 => x"C0C0C0A4F8808090",
 27890 => x"C0C0C0A4F88090C0",
 27891 => x"C0C0C0A4F88090F9",
 27892 => x"C0C0C0A4F88090A4",
 27893 => x"C0C0C0A4F88090B0",
 27894 => x"C0C0C0A4F8809099",
 27895 => x"C0C0C0A4F8809092",
 27896 => x"C0C0C0A4F8809082",
 27897 => x"C0C0C0A4F88090F8",
 27898 => x"C0C0C0A4F8809080",
 27899 => x"C0C0C0A4F8809090",
 27900 => x"C0C0C0A4F890C0C0",
 27901 => x"C0C0C0A4F890C0F9",
 27902 => x"C0C0C0A4F890C0A4",
 27903 => x"C0C0C0A4F890C0B0",
 27904 => x"C0C0C0A4F890C099",
 27905 => x"C0C0C0A4F890C092",
 27906 => x"C0C0C0A4F890C082",
 27907 => x"C0C0C0A4F890C0F8",
 27908 => x"C0C0C0A4F890C080",
 27909 => x"C0C0C0A4F890C090",
 27910 => x"C0C0C0A4F890F9C0",
 27911 => x"C0C0C0A4F890F9F9",
 27912 => x"C0C0C0A4F890F9A4",
 27913 => x"C0C0C0A4F890F9B0",
 27914 => x"C0C0C0A4F890F999",
 27915 => x"C0C0C0A4F890F992",
 27916 => x"C0C0C0A4F890F982",
 27917 => x"C0C0C0A4F890F9F8",
 27918 => x"C0C0C0A4F890F980",
 27919 => x"C0C0C0A4F890F990",
 27920 => x"C0C0C0A4F890A4C0",
 27921 => x"C0C0C0A4F890A4F9",
 27922 => x"C0C0C0A4F890A4A4",
 27923 => x"C0C0C0A4F890A4B0",
 27924 => x"C0C0C0A4F890A499",
 27925 => x"C0C0C0A4F890A492",
 27926 => x"C0C0C0A4F890A482",
 27927 => x"C0C0C0A4F890A4F8",
 27928 => x"C0C0C0A4F890A480",
 27929 => x"C0C0C0A4F890A490",
 27930 => x"C0C0C0A4F890B0C0",
 27931 => x"C0C0C0A4F890B0F9",
 27932 => x"C0C0C0A4F890B0A4",
 27933 => x"C0C0C0A4F890B0B0",
 27934 => x"C0C0C0A4F890B099",
 27935 => x"C0C0C0A4F890B092",
 27936 => x"C0C0C0A4F890B082",
 27937 => x"C0C0C0A4F890B0F8",
 27938 => x"C0C0C0A4F890B080",
 27939 => x"C0C0C0A4F890B090",
 27940 => x"C0C0C0A4F89099C0",
 27941 => x"C0C0C0A4F89099F9",
 27942 => x"C0C0C0A4F89099A4",
 27943 => x"C0C0C0A4F89099B0",
 27944 => x"C0C0C0A4F8909999",
 27945 => x"C0C0C0A4F8909992",
 27946 => x"C0C0C0A4F8909982",
 27947 => x"C0C0C0A4F89099F8",
 27948 => x"C0C0C0A4F8909980",
 27949 => x"C0C0C0A4F8909990",
 27950 => x"C0C0C0A4F89092C0",
 27951 => x"C0C0C0A4F89092F9",
 27952 => x"C0C0C0A4F89092A4",
 27953 => x"C0C0C0A4F89092B0",
 27954 => x"C0C0C0A4F8909299",
 27955 => x"C0C0C0A4F8909292",
 27956 => x"C0C0C0A4F8909282",
 27957 => x"C0C0C0A4F89092F8",
 27958 => x"C0C0C0A4F8909280",
 27959 => x"C0C0C0A4F8909290",
 27960 => x"C0C0C0A4F89082C0",
 27961 => x"C0C0C0A4F89082F9",
 27962 => x"C0C0C0A4F89082A4",
 27963 => x"C0C0C0A4F89082B0",
 27964 => x"C0C0C0A4F8908299",
 27965 => x"C0C0C0A4F8908292",
 27966 => x"C0C0C0A4F8908282",
 27967 => x"C0C0C0A4F89082F8",
 27968 => x"C0C0C0A4F8908280",
 27969 => x"C0C0C0A4F8908290",
 27970 => x"C0C0C0A4F890F8C0",
 27971 => x"C0C0C0A4F890F8F9",
 27972 => x"C0C0C0A4F890F8A4",
 27973 => x"C0C0C0A4F890F8B0",
 27974 => x"C0C0C0A4F890F899",
 27975 => x"C0C0C0A4F890F892",
 27976 => x"C0C0C0A4F890F882",
 27977 => x"C0C0C0A4F890F8F8",
 27978 => x"C0C0C0A4F890F880",
 27979 => x"C0C0C0A4F890F890",
 27980 => x"C0C0C0A4F89080C0",
 27981 => x"C0C0C0A4F89080F9",
 27982 => x"C0C0C0A4F89080A4",
 27983 => x"C0C0C0A4F89080B0",
 27984 => x"C0C0C0A4F8908099",
 27985 => x"C0C0C0A4F8908092",
 27986 => x"C0C0C0A4F8908082",
 27987 => x"C0C0C0A4F89080F8",
 27988 => x"C0C0C0A4F8908080",
 27989 => x"C0C0C0A4F8908090",
 27990 => x"C0C0C0A4F89090C0",
 27991 => x"C0C0C0A4F89090F9",
 27992 => x"C0C0C0A4F89090A4",
 27993 => x"C0C0C0A4F89090B0",
 27994 => x"C0C0C0A4F8909099",
 27995 => x"C0C0C0A4F8909092",
 27996 => x"C0C0C0A4F8909082",
 27997 => x"C0C0C0A4F89090F8",
 27998 => x"C0C0C0A4F8909080",
 27999 => x"C0C0C0A4F8909090",
 28000 => x"C0C0C0A480C0C0C0",
 28001 => x"C0C0C0A480C0C0F9",
 28002 => x"C0C0C0A480C0C0A4",
 28003 => x"C0C0C0A480C0C0B0",
 28004 => x"C0C0C0A480C0C099",
 28005 => x"C0C0C0A480C0C092",
 28006 => x"C0C0C0A480C0C082",
 28007 => x"C0C0C0A480C0C0F8",
 28008 => x"C0C0C0A480C0C080",
 28009 => x"C0C0C0A480C0C090",
 28010 => x"C0C0C0A480C0F9C0",
 28011 => x"C0C0C0A480C0F9F9",
 28012 => x"C0C0C0A480C0F9A4",
 28013 => x"C0C0C0A480C0F9B0",
 28014 => x"C0C0C0A480C0F999",
 28015 => x"C0C0C0A480C0F992",
 28016 => x"C0C0C0A480C0F982",
 28017 => x"C0C0C0A480C0F9F8",
 28018 => x"C0C0C0A480C0F980",
 28019 => x"C0C0C0A480C0F990",
 28020 => x"C0C0C0A480C0A4C0",
 28021 => x"C0C0C0A480C0A4F9",
 28022 => x"C0C0C0A480C0A4A4",
 28023 => x"C0C0C0A480C0A4B0",
 28024 => x"C0C0C0A480C0A499",
 28025 => x"C0C0C0A480C0A492",
 28026 => x"C0C0C0A480C0A482",
 28027 => x"C0C0C0A480C0A4F8",
 28028 => x"C0C0C0A480C0A480",
 28029 => x"C0C0C0A480C0A490",
 28030 => x"C0C0C0A480C0B0C0",
 28031 => x"C0C0C0A480C0B0F9",
 28032 => x"C0C0C0A480C0B0A4",
 28033 => x"C0C0C0A480C0B0B0",
 28034 => x"C0C0C0A480C0B099",
 28035 => x"C0C0C0A480C0B092",
 28036 => x"C0C0C0A480C0B082",
 28037 => x"C0C0C0A480C0B0F8",
 28038 => x"C0C0C0A480C0B080",
 28039 => x"C0C0C0A480C0B090",
 28040 => x"C0C0C0A480C099C0",
 28041 => x"C0C0C0A480C099F9",
 28042 => x"C0C0C0A480C099A4",
 28043 => x"C0C0C0A480C099B0",
 28044 => x"C0C0C0A480C09999",
 28045 => x"C0C0C0A480C09992",
 28046 => x"C0C0C0A480C09982",
 28047 => x"C0C0C0A480C099F8",
 28048 => x"C0C0C0A480C09980",
 28049 => x"C0C0C0A480C09990",
 28050 => x"C0C0C0A480C092C0",
 28051 => x"C0C0C0A480C092F9",
 28052 => x"C0C0C0A480C092A4",
 28053 => x"C0C0C0A480C092B0",
 28054 => x"C0C0C0A480C09299",
 28055 => x"C0C0C0A480C09292",
 28056 => x"C0C0C0A480C09282",
 28057 => x"C0C0C0A480C092F8",
 28058 => x"C0C0C0A480C09280",
 28059 => x"C0C0C0A480C09290",
 28060 => x"C0C0C0A480C082C0",
 28061 => x"C0C0C0A480C082F9",
 28062 => x"C0C0C0A480C082A4",
 28063 => x"C0C0C0A480C082B0",
 28064 => x"C0C0C0A480C08299",
 28065 => x"C0C0C0A480C08292",
 28066 => x"C0C0C0A480C08282",
 28067 => x"C0C0C0A480C082F8",
 28068 => x"C0C0C0A480C08280",
 28069 => x"C0C0C0A480C08290",
 28070 => x"C0C0C0A480C0F8C0",
 28071 => x"C0C0C0A480C0F8F9",
 28072 => x"C0C0C0A480C0F8A4",
 28073 => x"C0C0C0A480C0F8B0",
 28074 => x"C0C0C0A480C0F899",
 28075 => x"C0C0C0A480C0F892",
 28076 => x"C0C0C0A480C0F882",
 28077 => x"C0C0C0A480C0F8F8",
 28078 => x"C0C0C0A480C0F880",
 28079 => x"C0C0C0A480C0F890",
 28080 => x"C0C0C0A480C080C0",
 28081 => x"C0C0C0A480C080F9",
 28082 => x"C0C0C0A480C080A4",
 28083 => x"C0C0C0A480C080B0",
 28084 => x"C0C0C0A480C08099",
 28085 => x"C0C0C0A480C08092",
 28086 => x"C0C0C0A480C08082",
 28087 => x"C0C0C0A480C080F8",
 28088 => x"C0C0C0A480C08080",
 28089 => x"C0C0C0A480C08090",
 28090 => x"C0C0C0A480C090C0",
 28091 => x"C0C0C0A480C090F9",
 28092 => x"C0C0C0A480C090A4",
 28093 => x"C0C0C0A480C090B0",
 28094 => x"C0C0C0A480C09099",
 28095 => x"C0C0C0A480C09092",
 28096 => x"C0C0C0A480C09082",
 28097 => x"C0C0C0A480C090F8",
 28098 => x"C0C0C0A480C09080",
 28099 => x"C0C0C0A480C09090",
 28100 => x"C0C0C0A480F9C0C0",
 28101 => x"C0C0C0A480F9C0F9",
 28102 => x"C0C0C0A480F9C0A4",
 28103 => x"C0C0C0A480F9C0B0",
 28104 => x"C0C0C0A480F9C099",
 28105 => x"C0C0C0A480F9C092",
 28106 => x"C0C0C0A480F9C082",
 28107 => x"C0C0C0A480F9C0F8",
 28108 => x"C0C0C0A480F9C080",
 28109 => x"C0C0C0A480F9C090",
 28110 => x"C0C0C0A480F9F9C0",
 28111 => x"C0C0C0A480F9F9F9",
 28112 => x"C0C0C0A480F9F9A4",
 28113 => x"C0C0C0A480F9F9B0",
 28114 => x"C0C0C0A480F9F999",
 28115 => x"C0C0C0A480F9F992",
 28116 => x"C0C0C0A480F9F982",
 28117 => x"C0C0C0A480F9F9F8",
 28118 => x"C0C0C0A480F9F980",
 28119 => x"C0C0C0A480F9F990",
 28120 => x"C0C0C0A480F9A4C0",
 28121 => x"C0C0C0A480F9A4F9",
 28122 => x"C0C0C0A480F9A4A4",
 28123 => x"C0C0C0A480F9A4B0",
 28124 => x"C0C0C0A480F9A499",
 28125 => x"C0C0C0A480F9A492",
 28126 => x"C0C0C0A480F9A482",
 28127 => x"C0C0C0A480F9A4F8",
 28128 => x"C0C0C0A480F9A480",
 28129 => x"C0C0C0A480F9A490",
 28130 => x"C0C0C0A480F9B0C0",
 28131 => x"C0C0C0A480F9B0F9",
 28132 => x"C0C0C0A480F9B0A4",
 28133 => x"C0C0C0A480F9B0B0",
 28134 => x"C0C0C0A480F9B099",
 28135 => x"C0C0C0A480F9B092",
 28136 => x"C0C0C0A480F9B082",
 28137 => x"C0C0C0A480F9B0F8",
 28138 => x"C0C0C0A480F9B080",
 28139 => x"C0C0C0A480F9B090",
 28140 => x"C0C0C0A480F999C0",
 28141 => x"C0C0C0A480F999F9",
 28142 => x"C0C0C0A480F999A4",
 28143 => x"C0C0C0A480F999B0",
 28144 => x"C0C0C0A480F99999",
 28145 => x"C0C0C0A480F99992",
 28146 => x"C0C0C0A480F99982",
 28147 => x"C0C0C0A480F999F8",
 28148 => x"C0C0C0A480F99980",
 28149 => x"C0C0C0A480F99990",
 28150 => x"C0C0C0A480F992C0",
 28151 => x"C0C0C0A480F992F9",
 28152 => x"C0C0C0A480F992A4",
 28153 => x"C0C0C0A480F992B0",
 28154 => x"C0C0C0A480F99299",
 28155 => x"C0C0C0A480F99292",
 28156 => x"C0C0C0A480F99282",
 28157 => x"C0C0C0A480F992F8",
 28158 => x"C0C0C0A480F99280",
 28159 => x"C0C0C0A480F99290",
 28160 => x"C0C0C0A480F982C0",
 28161 => x"C0C0C0A480F982F9",
 28162 => x"C0C0C0A480F982A4",
 28163 => x"C0C0C0A480F982B0",
 28164 => x"C0C0C0A480F98299",
 28165 => x"C0C0C0A480F98292",
 28166 => x"C0C0C0A480F98282",
 28167 => x"C0C0C0A480F982F8",
 28168 => x"C0C0C0A480F98280",
 28169 => x"C0C0C0A480F98290",
 28170 => x"C0C0C0A480F9F8C0",
 28171 => x"C0C0C0A480F9F8F9",
 28172 => x"C0C0C0A480F9F8A4",
 28173 => x"C0C0C0A480F9F8B0",
 28174 => x"C0C0C0A480F9F899",
 28175 => x"C0C0C0A480F9F892",
 28176 => x"C0C0C0A480F9F882",
 28177 => x"C0C0C0A480F9F8F8",
 28178 => x"C0C0C0A480F9F880",
 28179 => x"C0C0C0A480F9F890",
 28180 => x"C0C0C0A480F980C0",
 28181 => x"C0C0C0A480F980F9",
 28182 => x"C0C0C0A480F980A4",
 28183 => x"C0C0C0A480F980B0",
 28184 => x"C0C0C0A480F98099",
 28185 => x"C0C0C0A480F98092",
 28186 => x"C0C0C0A480F98082",
 28187 => x"C0C0C0A480F980F8",
 28188 => x"C0C0C0A480F98080",
 28189 => x"C0C0C0A480F98090",
 28190 => x"C0C0C0A480F990C0",
 28191 => x"C0C0C0A480F990F9",
 28192 => x"C0C0C0A480F990A4",
 28193 => x"C0C0C0A480F990B0",
 28194 => x"C0C0C0A480F99099",
 28195 => x"C0C0C0A480F99092",
 28196 => x"C0C0C0A480F99082",
 28197 => x"C0C0C0A480F990F8",
 28198 => x"C0C0C0A480F99080",
 28199 => x"C0C0C0A480F99090",
 28200 => x"C0C0C0A480A4C0C0",
 28201 => x"C0C0C0A480A4C0F9",
 28202 => x"C0C0C0A480A4C0A4",
 28203 => x"C0C0C0A480A4C0B0",
 28204 => x"C0C0C0A480A4C099",
 28205 => x"C0C0C0A480A4C092",
 28206 => x"C0C0C0A480A4C082",
 28207 => x"C0C0C0A480A4C0F8",
 28208 => x"C0C0C0A480A4C080",
 28209 => x"C0C0C0A480A4C090",
 28210 => x"C0C0C0A480A4F9C0",
 28211 => x"C0C0C0A480A4F9F9",
 28212 => x"C0C0C0A480A4F9A4",
 28213 => x"C0C0C0A480A4F9B0",
 28214 => x"C0C0C0A480A4F999",
 28215 => x"C0C0C0A480A4F992",
 28216 => x"C0C0C0A480A4F982",
 28217 => x"C0C0C0A480A4F9F8",
 28218 => x"C0C0C0A480A4F980",
 28219 => x"C0C0C0A480A4F990",
 28220 => x"C0C0C0A480A4A4C0",
 28221 => x"C0C0C0A480A4A4F9",
 28222 => x"C0C0C0A480A4A4A4",
 28223 => x"C0C0C0A480A4A4B0",
 28224 => x"C0C0C0A480A4A499",
 28225 => x"C0C0C0A480A4A492",
 28226 => x"C0C0C0A480A4A482",
 28227 => x"C0C0C0A480A4A4F8",
 28228 => x"C0C0C0A480A4A480",
 28229 => x"C0C0C0A480A4A490",
 28230 => x"C0C0C0A480A4B0C0",
 28231 => x"C0C0C0A480A4B0F9",
 28232 => x"C0C0C0A480A4B0A4",
 28233 => x"C0C0C0A480A4B0B0",
 28234 => x"C0C0C0A480A4B099",
 28235 => x"C0C0C0A480A4B092",
 28236 => x"C0C0C0A480A4B082",
 28237 => x"C0C0C0A480A4B0F8",
 28238 => x"C0C0C0A480A4B080",
 28239 => x"C0C0C0A480A4B090",
 28240 => x"C0C0C0A480A499C0",
 28241 => x"C0C0C0A480A499F9",
 28242 => x"C0C0C0A480A499A4",
 28243 => x"C0C0C0A480A499B0",
 28244 => x"C0C0C0A480A49999",
 28245 => x"C0C0C0A480A49992",
 28246 => x"C0C0C0A480A49982",
 28247 => x"C0C0C0A480A499F8",
 28248 => x"C0C0C0A480A49980",
 28249 => x"C0C0C0A480A49990",
 28250 => x"C0C0C0A480A492C0",
 28251 => x"C0C0C0A480A492F9",
 28252 => x"C0C0C0A480A492A4",
 28253 => x"C0C0C0A480A492B0",
 28254 => x"C0C0C0A480A49299",
 28255 => x"C0C0C0A480A49292",
 28256 => x"C0C0C0A480A49282",
 28257 => x"C0C0C0A480A492F8",
 28258 => x"C0C0C0A480A49280",
 28259 => x"C0C0C0A480A49290",
 28260 => x"C0C0C0A480A482C0",
 28261 => x"C0C0C0A480A482F9",
 28262 => x"C0C0C0A480A482A4",
 28263 => x"C0C0C0A480A482B0",
 28264 => x"C0C0C0A480A48299",
 28265 => x"C0C0C0A480A48292",
 28266 => x"C0C0C0A480A48282",
 28267 => x"C0C0C0A480A482F8",
 28268 => x"C0C0C0A480A48280",
 28269 => x"C0C0C0A480A48290",
 28270 => x"C0C0C0A480A4F8C0",
 28271 => x"C0C0C0A480A4F8F9",
 28272 => x"C0C0C0A480A4F8A4",
 28273 => x"C0C0C0A480A4F8B0",
 28274 => x"C0C0C0A480A4F899",
 28275 => x"C0C0C0A480A4F892",
 28276 => x"C0C0C0A480A4F882",
 28277 => x"C0C0C0A480A4F8F8",
 28278 => x"C0C0C0A480A4F880",
 28279 => x"C0C0C0A480A4F890",
 28280 => x"C0C0C0A480A480C0",
 28281 => x"C0C0C0A480A480F9",
 28282 => x"C0C0C0A480A480A4",
 28283 => x"C0C0C0A480A480B0",
 28284 => x"C0C0C0A480A48099",
 28285 => x"C0C0C0A480A48092",
 28286 => x"C0C0C0A480A48082",
 28287 => x"C0C0C0A480A480F8",
 28288 => x"C0C0C0A480A48080",
 28289 => x"C0C0C0A480A48090",
 28290 => x"C0C0C0A480A490C0",
 28291 => x"C0C0C0A480A490F9",
 28292 => x"C0C0C0A480A490A4",
 28293 => x"C0C0C0A480A490B0",
 28294 => x"C0C0C0A480A49099",
 28295 => x"C0C0C0A480A49092",
 28296 => x"C0C0C0A480A49082",
 28297 => x"C0C0C0A480A490F8",
 28298 => x"C0C0C0A480A49080",
 28299 => x"C0C0C0A480A49090",
 28300 => x"C0C0C0A480B0C0C0",
 28301 => x"C0C0C0A480B0C0F9",
 28302 => x"C0C0C0A480B0C0A4",
 28303 => x"C0C0C0A480B0C0B0",
 28304 => x"C0C0C0A480B0C099",
 28305 => x"C0C0C0A480B0C092",
 28306 => x"C0C0C0A480B0C082",
 28307 => x"C0C0C0A480B0C0F8",
 28308 => x"C0C0C0A480B0C080",
 28309 => x"C0C0C0A480B0C090",
 28310 => x"C0C0C0A480B0F9C0",
 28311 => x"C0C0C0A480B0F9F9",
 28312 => x"C0C0C0A480B0F9A4",
 28313 => x"C0C0C0A480B0F9B0",
 28314 => x"C0C0C0A480B0F999",
 28315 => x"C0C0C0A480B0F992",
 28316 => x"C0C0C0A480B0F982",
 28317 => x"C0C0C0A480B0F9F8",
 28318 => x"C0C0C0A480B0F980",
 28319 => x"C0C0C0A480B0F990",
 28320 => x"C0C0C0A480B0A4C0",
 28321 => x"C0C0C0A480B0A4F9",
 28322 => x"C0C0C0A480B0A4A4",
 28323 => x"C0C0C0A480B0A4B0",
 28324 => x"C0C0C0A480B0A499",
 28325 => x"C0C0C0A480B0A492",
 28326 => x"C0C0C0A480B0A482",
 28327 => x"C0C0C0A480B0A4F8",
 28328 => x"C0C0C0A480B0A480",
 28329 => x"C0C0C0A480B0A490",
 28330 => x"C0C0C0A480B0B0C0",
 28331 => x"C0C0C0A480B0B0F9",
 28332 => x"C0C0C0A480B0B0A4",
 28333 => x"C0C0C0A480B0B0B0",
 28334 => x"C0C0C0A480B0B099",
 28335 => x"C0C0C0A480B0B092",
 28336 => x"C0C0C0A480B0B082",
 28337 => x"C0C0C0A480B0B0F8",
 28338 => x"C0C0C0A480B0B080",
 28339 => x"C0C0C0A480B0B090",
 28340 => x"C0C0C0A480B099C0",
 28341 => x"C0C0C0A480B099F9",
 28342 => x"C0C0C0A480B099A4",
 28343 => x"C0C0C0A480B099B0",
 28344 => x"C0C0C0A480B09999",
 28345 => x"C0C0C0A480B09992",
 28346 => x"C0C0C0A480B09982",
 28347 => x"C0C0C0A480B099F8",
 28348 => x"C0C0C0A480B09980",
 28349 => x"C0C0C0A480B09990",
 28350 => x"C0C0C0A480B092C0",
 28351 => x"C0C0C0A480B092F9",
 28352 => x"C0C0C0A480B092A4",
 28353 => x"C0C0C0A480B092B0",
 28354 => x"C0C0C0A480B09299",
 28355 => x"C0C0C0A480B09292",
 28356 => x"C0C0C0A480B09282",
 28357 => x"C0C0C0A480B092F8",
 28358 => x"C0C0C0A480B09280",
 28359 => x"C0C0C0A480B09290",
 28360 => x"C0C0C0A480B082C0",
 28361 => x"C0C0C0A480B082F9",
 28362 => x"C0C0C0A480B082A4",
 28363 => x"C0C0C0A480B082B0",
 28364 => x"C0C0C0A480B08299",
 28365 => x"C0C0C0A480B08292",
 28366 => x"C0C0C0A480B08282",
 28367 => x"C0C0C0A480B082F8",
 28368 => x"C0C0C0A480B08280",
 28369 => x"C0C0C0A480B08290",
 28370 => x"C0C0C0A480B0F8C0",
 28371 => x"C0C0C0A480B0F8F9",
 28372 => x"C0C0C0A480B0F8A4",
 28373 => x"C0C0C0A480B0F8B0",
 28374 => x"C0C0C0A480B0F899",
 28375 => x"C0C0C0A480B0F892",
 28376 => x"C0C0C0A480B0F882",
 28377 => x"C0C0C0A480B0F8F8",
 28378 => x"C0C0C0A480B0F880",
 28379 => x"C0C0C0A480B0F890",
 28380 => x"C0C0C0A480B080C0",
 28381 => x"C0C0C0A480B080F9",
 28382 => x"C0C0C0A480B080A4",
 28383 => x"C0C0C0A480B080B0",
 28384 => x"C0C0C0A480B08099",
 28385 => x"C0C0C0A480B08092",
 28386 => x"C0C0C0A480B08082",
 28387 => x"C0C0C0A480B080F8",
 28388 => x"C0C0C0A480B08080",
 28389 => x"C0C0C0A480B08090",
 28390 => x"C0C0C0A480B090C0",
 28391 => x"C0C0C0A480B090F9",
 28392 => x"C0C0C0A480B090A4",
 28393 => x"C0C0C0A480B090B0",
 28394 => x"C0C0C0A480B09099",
 28395 => x"C0C0C0A480B09092",
 28396 => x"C0C0C0A480B09082",
 28397 => x"C0C0C0A480B090F8",
 28398 => x"C0C0C0A480B09080",
 28399 => x"C0C0C0A480B09090",
 28400 => x"C0C0C0A48099C0C0",
 28401 => x"C0C0C0A48099C0F9",
 28402 => x"C0C0C0A48099C0A4",
 28403 => x"C0C0C0A48099C0B0",
 28404 => x"C0C0C0A48099C099",
 28405 => x"C0C0C0A48099C092",
 28406 => x"C0C0C0A48099C082",
 28407 => x"C0C0C0A48099C0F8",
 28408 => x"C0C0C0A48099C080",
 28409 => x"C0C0C0A48099C090",
 28410 => x"C0C0C0A48099F9C0",
 28411 => x"C0C0C0A48099F9F9",
 28412 => x"C0C0C0A48099F9A4",
 28413 => x"C0C0C0A48099F9B0",
 28414 => x"C0C0C0A48099F999",
 28415 => x"C0C0C0A48099F992",
 28416 => x"C0C0C0A48099F982",
 28417 => x"C0C0C0A48099F9F8",
 28418 => x"C0C0C0A48099F980",
 28419 => x"C0C0C0A48099F990",
 28420 => x"C0C0C0A48099A4C0",
 28421 => x"C0C0C0A48099A4F9",
 28422 => x"C0C0C0A48099A4A4",
 28423 => x"C0C0C0A48099A4B0",
 28424 => x"C0C0C0A48099A499",
 28425 => x"C0C0C0A48099A492",
 28426 => x"C0C0C0A48099A482",
 28427 => x"C0C0C0A48099A4F8",
 28428 => x"C0C0C0A48099A480",
 28429 => x"C0C0C0A48099A490",
 28430 => x"C0C0C0A48099B0C0",
 28431 => x"C0C0C0A48099B0F9",
 28432 => x"C0C0C0A48099B0A4",
 28433 => x"C0C0C0A48099B0B0",
 28434 => x"C0C0C0A48099B099",
 28435 => x"C0C0C0A48099B092",
 28436 => x"C0C0C0A48099B082",
 28437 => x"C0C0C0A48099B0F8",
 28438 => x"C0C0C0A48099B080",
 28439 => x"C0C0C0A48099B090",
 28440 => x"C0C0C0A4809999C0",
 28441 => x"C0C0C0A4809999F9",
 28442 => x"C0C0C0A4809999A4",
 28443 => x"C0C0C0A4809999B0",
 28444 => x"C0C0C0A480999999",
 28445 => x"C0C0C0A480999992",
 28446 => x"C0C0C0A480999982",
 28447 => x"C0C0C0A4809999F8",
 28448 => x"C0C0C0A480999980",
 28449 => x"C0C0C0A480999990",
 28450 => x"C0C0C0A4809992C0",
 28451 => x"C0C0C0A4809992F9",
 28452 => x"C0C0C0A4809992A4",
 28453 => x"C0C0C0A4809992B0",
 28454 => x"C0C0C0A480999299",
 28455 => x"C0C0C0A480999292",
 28456 => x"C0C0C0A480999282",
 28457 => x"C0C0C0A4809992F8",
 28458 => x"C0C0C0A480999280",
 28459 => x"C0C0C0A480999290",
 28460 => x"C0C0C0A4809982C0",
 28461 => x"C0C0C0A4809982F9",
 28462 => x"C0C0C0A4809982A4",
 28463 => x"C0C0C0A4809982B0",
 28464 => x"C0C0C0A480998299",
 28465 => x"C0C0C0A480998292",
 28466 => x"C0C0C0A480998282",
 28467 => x"C0C0C0A4809982F8",
 28468 => x"C0C0C0A480998280",
 28469 => x"C0C0C0A480998290",
 28470 => x"C0C0C0A48099F8C0",
 28471 => x"C0C0C0A48099F8F9",
 28472 => x"C0C0C0A48099F8A4",
 28473 => x"C0C0C0A48099F8B0",
 28474 => x"C0C0C0A48099F899",
 28475 => x"C0C0C0A48099F892",
 28476 => x"C0C0C0A48099F882",
 28477 => x"C0C0C0A48099F8F8",
 28478 => x"C0C0C0A48099F880",
 28479 => x"C0C0C0A48099F890",
 28480 => x"C0C0C0A4809980C0",
 28481 => x"C0C0C0A4809980F9",
 28482 => x"C0C0C0A4809980A4",
 28483 => x"C0C0C0A4809980B0",
 28484 => x"C0C0C0A480998099",
 28485 => x"C0C0C0A480998092",
 28486 => x"C0C0C0A480998082",
 28487 => x"C0C0C0A4809980F8",
 28488 => x"C0C0C0A480998080",
 28489 => x"C0C0C0A480998090",
 28490 => x"C0C0C0A4809990C0",
 28491 => x"C0C0C0A4809990F9",
 28492 => x"C0C0C0A4809990A4",
 28493 => x"C0C0C0A4809990B0",
 28494 => x"C0C0C0A480999099",
 28495 => x"C0C0C0A480999092",
 28496 => x"C0C0C0A480999082",
 28497 => x"C0C0C0A4809990F8",
 28498 => x"C0C0C0A480999080",
 28499 => x"C0C0C0A480999090",
 28500 => x"C0C0C0A48092C0C0",
 28501 => x"C0C0C0A48092C0F9",
 28502 => x"C0C0C0A48092C0A4",
 28503 => x"C0C0C0A48092C0B0",
 28504 => x"C0C0C0A48092C099",
 28505 => x"C0C0C0A48092C092",
 28506 => x"C0C0C0A48092C082",
 28507 => x"C0C0C0A48092C0F8",
 28508 => x"C0C0C0A48092C080",
 28509 => x"C0C0C0A48092C090",
 28510 => x"C0C0C0A48092F9C0",
 28511 => x"C0C0C0A48092F9F9",
 28512 => x"C0C0C0A48092F9A4",
 28513 => x"C0C0C0A48092F9B0",
 28514 => x"C0C0C0A48092F999",
 28515 => x"C0C0C0A48092F992",
 28516 => x"C0C0C0A48092F982",
 28517 => x"C0C0C0A48092F9F8",
 28518 => x"C0C0C0A48092F980",
 28519 => x"C0C0C0A48092F990",
 28520 => x"C0C0C0A48092A4C0",
 28521 => x"C0C0C0A48092A4F9",
 28522 => x"C0C0C0A48092A4A4",
 28523 => x"C0C0C0A48092A4B0",
 28524 => x"C0C0C0A48092A499",
 28525 => x"C0C0C0A48092A492",
 28526 => x"C0C0C0A48092A482",
 28527 => x"C0C0C0A48092A4F8",
 28528 => x"C0C0C0A48092A480",
 28529 => x"C0C0C0A48092A490",
 28530 => x"C0C0C0A48092B0C0",
 28531 => x"C0C0C0A48092B0F9",
 28532 => x"C0C0C0A48092B0A4",
 28533 => x"C0C0C0A48092B0B0",
 28534 => x"C0C0C0A48092B099",
 28535 => x"C0C0C0A48092B092",
 28536 => x"C0C0C0A48092B082",
 28537 => x"C0C0C0A48092B0F8",
 28538 => x"C0C0C0A48092B080",
 28539 => x"C0C0C0A48092B090",
 28540 => x"C0C0C0A4809299C0",
 28541 => x"C0C0C0A4809299F9",
 28542 => x"C0C0C0A4809299A4",
 28543 => x"C0C0C0A4809299B0",
 28544 => x"C0C0C0A480929999",
 28545 => x"C0C0C0A480929992",
 28546 => x"C0C0C0A480929982",
 28547 => x"C0C0C0A4809299F8",
 28548 => x"C0C0C0A480929980",
 28549 => x"C0C0C0A480929990",
 28550 => x"C0C0C0A4809292C0",
 28551 => x"C0C0C0A4809292F9",
 28552 => x"C0C0C0A4809292A4",
 28553 => x"C0C0C0A4809292B0",
 28554 => x"C0C0C0A480929299",
 28555 => x"C0C0C0A480929292",
 28556 => x"C0C0C0A480929282",
 28557 => x"C0C0C0A4809292F8",
 28558 => x"C0C0C0A480929280",
 28559 => x"C0C0C0A480929290",
 28560 => x"C0C0C0A4809282C0",
 28561 => x"C0C0C0A4809282F9",
 28562 => x"C0C0C0A4809282A4",
 28563 => x"C0C0C0A4809282B0",
 28564 => x"C0C0C0A480928299",
 28565 => x"C0C0C0A480928292",
 28566 => x"C0C0C0A480928282",
 28567 => x"C0C0C0A4809282F8",
 28568 => x"C0C0C0A480928280",
 28569 => x"C0C0C0A480928290",
 28570 => x"C0C0C0A48092F8C0",
 28571 => x"C0C0C0A48092F8F9",
 28572 => x"C0C0C0A48092F8A4",
 28573 => x"C0C0C0A48092F8B0",
 28574 => x"C0C0C0A48092F899",
 28575 => x"C0C0C0A48092F892",
 28576 => x"C0C0C0A48092F882",
 28577 => x"C0C0C0A48092F8F8",
 28578 => x"C0C0C0A48092F880",
 28579 => x"C0C0C0A48092F890",
 28580 => x"C0C0C0A4809280C0",
 28581 => x"C0C0C0A4809280F9",
 28582 => x"C0C0C0A4809280A4",
 28583 => x"C0C0C0A4809280B0",
 28584 => x"C0C0C0A480928099",
 28585 => x"C0C0C0A480928092",
 28586 => x"C0C0C0A480928082",
 28587 => x"C0C0C0A4809280F8",
 28588 => x"C0C0C0A480928080",
 28589 => x"C0C0C0A480928090",
 28590 => x"C0C0C0A4809290C0",
 28591 => x"C0C0C0A4809290F9",
 28592 => x"C0C0C0A4809290A4",
 28593 => x"C0C0C0A4809290B0",
 28594 => x"C0C0C0A480929099",
 28595 => x"C0C0C0A480929092",
 28596 => x"C0C0C0A480929082",
 28597 => x"C0C0C0A4809290F8",
 28598 => x"C0C0C0A480929080",
 28599 => x"C0C0C0A480929090",
 28600 => x"C0C0C0A48082C0C0",
 28601 => x"C0C0C0A48082C0F9",
 28602 => x"C0C0C0A48082C0A4",
 28603 => x"C0C0C0A48082C0B0",
 28604 => x"C0C0C0A48082C099",
 28605 => x"C0C0C0A48082C092",
 28606 => x"C0C0C0A48082C082",
 28607 => x"C0C0C0A48082C0F8",
 28608 => x"C0C0C0A48082C080",
 28609 => x"C0C0C0A48082C090",
 28610 => x"C0C0C0A48082F9C0",
 28611 => x"C0C0C0A48082F9F9",
 28612 => x"C0C0C0A48082F9A4",
 28613 => x"C0C0C0A48082F9B0",
 28614 => x"C0C0C0A48082F999",
 28615 => x"C0C0C0A48082F992",
 28616 => x"C0C0C0A48082F982",
 28617 => x"C0C0C0A48082F9F8",
 28618 => x"C0C0C0A48082F980",
 28619 => x"C0C0C0A48082F990",
 28620 => x"C0C0C0A48082A4C0",
 28621 => x"C0C0C0A48082A4F9",
 28622 => x"C0C0C0A48082A4A4",
 28623 => x"C0C0C0A48082A4B0",
 28624 => x"C0C0C0A48082A499",
 28625 => x"C0C0C0A48082A492",
 28626 => x"C0C0C0A48082A482",
 28627 => x"C0C0C0A48082A4F8",
 28628 => x"C0C0C0A48082A480",
 28629 => x"C0C0C0A48082A490",
 28630 => x"C0C0C0A48082B0C0",
 28631 => x"C0C0C0A48082B0F9",
 28632 => x"C0C0C0A48082B0A4",
 28633 => x"C0C0C0A48082B0B0",
 28634 => x"C0C0C0A48082B099",
 28635 => x"C0C0C0A48082B092",
 28636 => x"C0C0C0A48082B082",
 28637 => x"C0C0C0A48082B0F8",
 28638 => x"C0C0C0A48082B080",
 28639 => x"C0C0C0A48082B090",
 28640 => x"C0C0C0A4808299C0",
 28641 => x"C0C0C0A4808299F9",
 28642 => x"C0C0C0A4808299A4",
 28643 => x"C0C0C0A4808299B0",
 28644 => x"C0C0C0A480829999",
 28645 => x"C0C0C0A480829992",
 28646 => x"C0C0C0A480829982",
 28647 => x"C0C0C0A4808299F8",
 28648 => x"C0C0C0A480829980",
 28649 => x"C0C0C0A480829990",
 28650 => x"C0C0C0A4808292C0",
 28651 => x"C0C0C0A4808292F9",
 28652 => x"C0C0C0A4808292A4",
 28653 => x"C0C0C0A4808292B0",
 28654 => x"C0C0C0A480829299",
 28655 => x"C0C0C0A480829292",
 28656 => x"C0C0C0A480829282",
 28657 => x"C0C0C0A4808292F8",
 28658 => x"C0C0C0A480829280",
 28659 => x"C0C0C0A480829290",
 28660 => x"C0C0C0A4808282C0",
 28661 => x"C0C0C0A4808282F9",
 28662 => x"C0C0C0A4808282A4",
 28663 => x"C0C0C0A4808282B0",
 28664 => x"C0C0C0A480828299",
 28665 => x"C0C0C0A480828292",
 28666 => x"C0C0C0A480828282",
 28667 => x"C0C0C0A4808282F8",
 28668 => x"C0C0C0A480828280",
 28669 => x"C0C0C0A480828290",
 28670 => x"C0C0C0A48082F8C0",
 28671 => x"C0C0C0A48082F8F9",
 28672 => x"C0C0C0A48082F8A4",
 28673 => x"C0C0C0A48082F8B0",
 28674 => x"C0C0C0A48082F899",
 28675 => x"C0C0C0A48082F892",
 28676 => x"C0C0C0A48082F882",
 28677 => x"C0C0C0A48082F8F8",
 28678 => x"C0C0C0A48082F880",
 28679 => x"C0C0C0A48082F890",
 28680 => x"C0C0C0A4808280C0",
 28681 => x"C0C0C0A4808280F9",
 28682 => x"C0C0C0A4808280A4",
 28683 => x"C0C0C0A4808280B0",
 28684 => x"C0C0C0A480828099",
 28685 => x"C0C0C0A480828092",
 28686 => x"C0C0C0A480828082",
 28687 => x"C0C0C0A4808280F8",
 28688 => x"C0C0C0A480828080",
 28689 => x"C0C0C0A480828090",
 28690 => x"C0C0C0A4808290C0",
 28691 => x"C0C0C0A4808290F9",
 28692 => x"C0C0C0A4808290A4",
 28693 => x"C0C0C0A4808290B0",
 28694 => x"C0C0C0A480829099",
 28695 => x"C0C0C0A480829092",
 28696 => x"C0C0C0A480829082",
 28697 => x"C0C0C0A4808290F8",
 28698 => x"C0C0C0A480829080",
 28699 => x"C0C0C0A480829090",
 28700 => x"C0C0C0A480F8C0C0",
 28701 => x"C0C0C0A480F8C0F9",
 28702 => x"C0C0C0A480F8C0A4",
 28703 => x"C0C0C0A480F8C0B0",
 28704 => x"C0C0C0A480F8C099",
 28705 => x"C0C0C0A480F8C092",
 28706 => x"C0C0C0A480F8C082",
 28707 => x"C0C0C0A480F8C0F8",
 28708 => x"C0C0C0A480F8C080",
 28709 => x"C0C0C0A480F8C090",
 28710 => x"C0C0C0A480F8F9C0",
 28711 => x"C0C0C0A480F8F9F9",
 28712 => x"C0C0C0A480F8F9A4",
 28713 => x"C0C0C0A480F8F9B0",
 28714 => x"C0C0C0A480F8F999",
 28715 => x"C0C0C0A480F8F992",
 28716 => x"C0C0C0A480F8F982",
 28717 => x"C0C0C0A480F8F9F8",
 28718 => x"C0C0C0A480F8F980",
 28719 => x"C0C0C0A480F8F990",
 28720 => x"C0C0C0A480F8A4C0",
 28721 => x"C0C0C0A480F8A4F9",
 28722 => x"C0C0C0A480F8A4A4",
 28723 => x"C0C0C0A480F8A4B0",
 28724 => x"C0C0C0A480F8A499",
 28725 => x"C0C0C0A480F8A492",
 28726 => x"C0C0C0A480F8A482",
 28727 => x"C0C0C0A480F8A4F8",
 28728 => x"C0C0C0A480F8A480",
 28729 => x"C0C0C0A480F8A490",
 28730 => x"C0C0C0A480F8B0C0",
 28731 => x"C0C0C0A480F8B0F9",
 28732 => x"C0C0C0A480F8B0A4",
 28733 => x"C0C0C0A480F8B0B0",
 28734 => x"C0C0C0A480F8B099",
 28735 => x"C0C0C0A480F8B092",
 28736 => x"C0C0C0A480F8B082",
 28737 => x"C0C0C0A480F8B0F8",
 28738 => x"C0C0C0A480F8B080",
 28739 => x"C0C0C0A480F8B090",
 28740 => x"C0C0C0A480F899C0",
 28741 => x"C0C0C0A480F899F9",
 28742 => x"C0C0C0A480F899A4",
 28743 => x"C0C0C0A480F899B0",
 28744 => x"C0C0C0A480F89999",
 28745 => x"C0C0C0A480F89992",
 28746 => x"C0C0C0A480F89982",
 28747 => x"C0C0C0A480F899F8",
 28748 => x"C0C0C0A480F89980",
 28749 => x"C0C0C0A480F89990",
 28750 => x"C0C0C0A480F892C0",
 28751 => x"C0C0C0A480F892F9",
 28752 => x"C0C0C0A480F892A4",
 28753 => x"C0C0C0A480F892B0",
 28754 => x"C0C0C0A480F89299",
 28755 => x"C0C0C0A480F89292",
 28756 => x"C0C0C0A480F89282",
 28757 => x"C0C0C0A480F892F8",
 28758 => x"C0C0C0A480F89280",
 28759 => x"C0C0C0A480F89290",
 28760 => x"C0C0C0A480F882C0",
 28761 => x"C0C0C0A480F882F9",
 28762 => x"C0C0C0A480F882A4",
 28763 => x"C0C0C0A480F882B0",
 28764 => x"C0C0C0A480F88299",
 28765 => x"C0C0C0A480F88292",
 28766 => x"C0C0C0A480F88282",
 28767 => x"C0C0C0A480F882F8",
 28768 => x"C0C0C0A480F88280",
 28769 => x"C0C0C0A480F88290",
 28770 => x"C0C0C0A480F8F8C0",
 28771 => x"C0C0C0A480F8F8F9",
 28772 => x"C0C0C0A480F8F8A4",
 28773 => x"C0C0C0A480F8F8B0",
 28774 => x"C0C0C0A480F8F899",
 28775 => x"C0C0C0A480F8F892",
 28776 => x"C0C0C0A480F8F882",
 28777 => x"C0C0C0A480F8F8F8",
 28778 => x"C0C0C0A480F8F880",
 28779 => x"C0C0C0A480F8F890",
 28780 => x"C0C0C0A480F880C0",
 28781 => x"C0C0C0A480F880F9",
 28782 => x"C0C0C0A480F880A4",
 28783 => x"C0C0C0A480F880B0",
 28784 => x"C0C0C0A480F88099",
 28785 => x"C0C0C0A480F88092",
 28786 => x"C0C0C0A480F88082",
 28787 => x"C0C0C0A480F880F8",
 28788 => x"C0C0C0A480F88080",
 28789 => x"C0C0C0A480F88090",
 28790 => x"C0C0C0A480F890C0",
 28791 => x"C0C0C0A480F890F9",
 28792 => x"C0C0C0A480F890A4",
 28793 => x"C0C0C0A480F890B0",
 28794 => x"C0C0C0A480F89099",
 28795 => x"C0C0C0A480F89092",
 28796 => x"C0C0C0A480F89082",
 28797 => x"C0C0C0A480F890F8",
 28798 => x"C0C0C0A480F89080",
 28799 => x"C0C0C0A480F89090",
 28800 => x"C0C0C0A48080C0C0",
 28801 => x"C0C0C0A48080C0F9",
 28802 => x"C0C0C0A48080C0A4",
 28803 => x"C0C0C0A48080C0B0",
 28804 => x"C0C0C0A48080C099",
 28805 => x"C0C0C0A48080C092",
 28806 => x"C0C0C0A48080C082",
 28807 => x"C0C0C0A48080C0F8",
 28808 => x"C0C0C0A48080C080",
 28809 => x"C0C0C0A48080C090",
 28810 => x"C0C0C0A48080F9C0",
 28811 => x"C0C0C0A48080F9F9",
 28812 => x"C0C0C0A48080F9A4",
 28813 => x"C0C0C0A48080F9B0",
 28814 => x"C0C0C0A48080F999",
 28815 => x"C0C0C0A48080F992",
 28816 => x"C0C0C0A48080F982",
 28817 => x"C0C0C0A48080F9F8",
 28818 => x"C0C0C0A48080F980",
 28819 => x"C0C0C0A48080F990",
 28820 => x"C0C0C0A48080A4C0",
 28821 => x"C0C0C0A48080A4F9",
 28822 => x"C0C0C0A48080A4A4",
 28823 => x"C0C0C0A48080A4B0",
 28824 => x"C0C0C0A48080A499",
 28825 => x"C0C0C0A48080A492",
 28826 => x"C0C0C0A48080A482",
 28827 => x"C0C0C0A48080A4F8",
 28828 => x"C0C0C0A48080A480",
 28829 => x"C0C0C0A48080A490",
 28830 => x"C0C0C0A48080B0C0",
 28831 => x"C0C0C0A48080B0F9",
 28832 => x"C0C0C0A48080B0A4",
 28833 => x"C0C0C0A48080B0B0",
 28834 => x"C0C0C0A48080B099",
 28835 => x"C0C0C0A48080B092",
 28836 => x"C0C0C0A48080B082",
 28837 => x"C0C0C0A48080B0F8",
 28838 => x"C0C0C0A48080B080",
 28839 => x"C0C0C0A48080B090",
 28840 => x"C0C0C0A4808099C0",
 28841 => x"C0C0C0A4808099F9",
 28842 => x"C0C0C0A4808099A4",
 28843 => x"C0C0C0A4808099B0",
 28844 => x"C0C0C0A480809999",
 28845 => x"C0C0C0A480809992",
 28846 => x"C0C0C0A480809982",
 28847 => x"C0C0C0A4808099F8",
 28848 => x"C0C0C0A480809980",
 28849 => x"C0C0C0A480809990",
 28850 => x"C0C0C0A4808092C0",
 28851 => x"C0C0C0A4808092F9",
 28852 => x"C0C0C0A4808092A4",
 28853 => x"C0C0C0A4808092B0",
 28854 => x"C0C0C0A480809299",
 28855 => x"C0C0C0A480809292",
 28856 => x"C0C0C0A480809282",
 28857 => x"C0C0C0A4808092F8",
 28858 => x"C0C0C0A480809280",
 28859 => x"C0C0C0A480809290",
 28860 => x"C0C0C0A4808082C0",
 28861 => x"C0C0C0A4808082F9",
 28862 => x"C0C0C0A4808082A4",
 28863 => x"C0C0C0A4808082B0",
 28864 => x"C0C0C0A480808299",
 28865 => x"C0C0C0A480808292",
 28866 => x"C0C0C0A480808282",
 28867 => x"C0C0C0A4808082F8",
 28868 => x"C0C0C0A480808280",
 28869 => x"C0C0C0A480808290",
 28870 => x"C0C0C0A48080F8C0",
 28871 => x"C0C0C0A48080F8F9",
 28872 => x"C0C0C0A48080F8A4",
 28873 => x"C0C0C0A48080F8B0",
 28874 => x"C0C0C0A48080F899",
 28875 => x"C0C0C0A48080F892",
 28876 => x"C0C0C0A48080F882",
 28877 => x"C0C0C0A48080F8F8",
 28878 => x"C0C0C0A48080F880",
 28879 => x"C0C0C0A48080F890",
 28880 => x"C0C0C0A4808080C0",
 28881 => x"C0C0C0A4808080F9",
 28882 => x"C0C0C0A4808080A4",
 28883 => x"C0C0C0A4808080B0",
 28884 => x"C0C0C0A480808099",
 28885 => x"C0C0C0A480808092",
 28886 => x"C0C0C0A480808082",
 28887 => x"C0C0C0A4808080F8",
 28888 => x"C0C0C0A480808080",
 28889 => x"C0C0C0A480808090",
 28890 => x"C0C0C0A4808090C0",
 28891 => x"C0C0C0A4808090F9",
 28892 => x"C0C0C0A4808090A4",
 28893 => x"C0C0C0A4808090B0",
 28894 => x"C0C0C0A480809099",
 28895 => x"C0C0C0A480809092",
 28896 => x"C0C0C0A480809082",
 28897 => x"C0C0C0A4808090F8",
 28898 => x"C0C0C0A480809080",
 28899 => x"C0C0C0A480809090",
 28900 => x"C0C0C0A48090C0C0",
 28901 => x"C0C0C0A48090C0F9",
 28902 => x"C0C0C0A48090C0A4",
 28903 => x"C0C0C0A48090C0B0",
 28904 => x"C0C0C0A48090C099",
 28905 => x"C0C0C0A48090C092",
 28906 => x"C0C0C0A48090C082",
 28907 => x"C0C0C0A48090C0F8",
 28908 => x"C0C0C0A48090C080",
 28909 => x"C0C0C0A48090C090",
 28910 => x"C0C0C0A48090F9C0",
 28911 => x"C0C0C0A48090F9F9",
 28912 => x"C0C0C0A48090F9A4",
 28913 => x"C0C0C0A48090F9B0",
 28914 => x"C0C0C0A48090F999",
 28915 => x"C0C0C0A48090F992",
 28916 => x"C0C0C0A48090F982",
 28917 => x"C0C0C0A48090F9F8",
 28918 => x"C0C0C0A48090F980",
 28919 => x"C0C0C0A48090F990",
 28920 => x"C0C0C0A48090A4C0",
 28921 => x"C0C0C0A48090A4F9",
 28922 => x"C0C0C0A48090A4A4",
 28923 => x"C0C0C0A48090A4B0",
 28924 => x"C0C0C0A48090A499",
 28925 => x"C0C0C0A48090A492",
 28926 => x"C0C0C0A48090A482",
 28927 => x"C0C0C0A48090A4F8",
 28928 => x"C0C0C0A48090A480",
 28929 => x"C0C0C0A48090A490",
 28930 => x"C0C0C0A48090B0C0",
 28931 => x"C0C0C0A48090B0F9",
 28932 => x"C0C0C0A48090B0A4",
 28933 => x"C0C0C0A48090B0B0",
 28934 => x"C0C0C0A48090B099",
 28935 => x"C0C0C0A48090B092",
 28936 => x"C0C0C0A48090B082",
 28937 => x"C0C0C0A48090B0F8",
 28938 => x"C0C0C0A48090B080",
 28939 => x"C0C0C0A48090B090",
 28940 => x"C0C0C0A4809099C0",
 28941 => x"C0C0C0A4809099F9",
 28942 => x"C0C0C0A4809099A4",
 28943 => x"C0C0C0A4809099B0",
 28944 => x"C0C0C0A480909999",
 28945 => x"C0C0C0A480909992",
 28946 => x"C0C0C0A480909982",
 28947 => x"C0C0C0A4809099F8",
 28948 => x"C0C0C0A480909980",
 28949 => x"C0C0C0A480909990",
 28950 => x"C0C0C0A4809092C0",
 28951 => x"C0C0C0A4809092F9",
 28952 => x"C0C0C0A4809092A4",
 28953 => x"C0C0C0A4809092B0",
 28954 => x"C0C0C0A480909299",
 28955 => x"C0C0C0A480909292",
 28956 => x"C0C0C0A480909282",
 28957 => x"C0C0C0A4809092F8",
 28958 => x"C0C0C0A480909280",
 28959 => x"C0C0C0A480909290",
 28960 => x"C0C0C0A4809082C0",
 28961 => x"C0C0C0A4809082F9",
 28962 => x"C0C0C0A4809082A4",
 28963 => x"C0C0C0A4809082B0",
 28964 => x"C0C0C0A480908299",
 28965 => x"C0C0C0A480908292",
 28966 => x"C0C0C0A480908282",
 28967 => x"C0C0C0A4809082F8",
 28968 => x"C0C0C0A480908280",
 28969 => x"C0C0C0A480908290",
 28970 => x"C0C0C0A48090F8C0",
 28971 => x"C0C0C0A48090F8F9",
 28972 => x"C0C0C0A48090F8A4",
 28973 => x"C0C0C0A48090F8B0",
 28974 => x"C0C0C0A48090F899",
 28975 => x"C0C0C0A48090F892",
 28976 => x"C0C0C0A48090F882",
 28977 => x"C0C0C0A48090F8F8",
 28978 => x"C0C0C0A48090F880",
 28979 => x"C0C0C0A48090F890",
 28980 => x"C0C0C0A4809080C0",
 28981 => x"C0C0C0A4809080F9",
 28982 => x"C0C0C0A4809080A4",
 28983 => x"C0C0C0A4809080B0",
 28984 => x"C0C0C0A480908099",
 28985 => x"C0C0C0A480908092",
 28986 => x"C0C0C0A480908082",
 28987 => x"C0C0C0A4809080F8",
 28988 => x"C0C0C0A480908080",
 28989 => x"C0C0C0A480908090",
 28990 => x"C0C0C0A4809090C0",
 28991 => x"C0C0C0A4809090F9",
 28992 => x"C0C0C0A4809090A4",
 28993 => x"C0C0C0A4809090B0",
 28994 => x"C0C0C0A480909099",
 28995 => x"C0C0C0A480909092",
 28996 => x"C0C0C0A480909082",
 28997 => x"C0C0C0A4809090F8",
 28998 => x"C0C0C0A480909080",
 28999 => x"C0C0C0A480909090",
 29000 => x"C0C0C0A490C0C0C0",
 29001 => x"C0C0C0A490C0C0F9",
 29002 => x"C0C0C0A490C0C0A4",
 29003 => x"C0C0C0A490C0C0B0",
 29004 => x"C0C0C0A490C0C099",
 29005 => x"C0C0C0A490C0C092",
 29006 => x"C0C0C0A490C0C082",
 29007 => x"C0C0C0A490C0C0F8",
 29008 => x"C0C0C0A490C0C080",
 29009 => x"C0C0C0A490C0C090",
 29010 => x"C0C0C0A490C0F9C0",
 29011 => x"C0C0C0A490C0F9F9",
 29012 => x"C0C0C0A490C0F9A4",
 29013 => x"C0C0C0A490C0F9B0",
 29014 => x"C0C0C0A490C0F999",
 29015 => x"C0C0C0A490C0F992",
 29016 => x"C0C0C0A490C0F982",
 29017 => x"C0C0C0A490C0F9F8",
 29018 => x"C0C0C0A490C0F980",
 29019 => x"C0C0C0A490C0F990",
 29020 => x"C0C0C0A490C0A4C0",
 29021 => x"C0C0C0A490C0A4F9",
 29022 => x"C0C0C0A490C0A4A4",
 29023 => x"C0C0C0A490C0A4B0",
 29024 => x"C0C0C0A490C0A499",
 29025 => x"C0C0C0A490C0A492",
 29026 => x"C0C0C0A490C0A482",
 29027 => x"C0C0C0A490C0A4F8",
 29028 => x"C0C0C0A490C0A480",
 29029 => x"C0C0C0A490C0A490",
 29030 => x"C0C0C0A490C0B0C0",
 29031 => x"C0C0C0A490C0B0F9",
 29032 => x"C0C0C0A490C0B0A4",
 29033 => x"C0C0C0A490C0B0B0",
 29034 => x"C0C0C0A490C0B099",
 29035 => x"C0C0C0A490C0B092",
 29036 => x"C0C0C0A490C0B082",
 29037 => x"C0C0C0A490C0B0F8",
 29038 => x"C0C0C0A490C0B080",
 29039 => x"C0C0C0A490C0B090",
 29040 => x"C0C0C0A490C099C0",
 29041 => x"C0C0C0A490C099F9",
 29042 => x"C0C0C0A490C099A4",
 29043 => x"C0C0C0A490C099B0",
 29044 => x"C0C0C0A490C09999",
 29045 => x"C0C0C0A490C09992",
 29046 => x"C0C0C0A490C09982",
 29047 => x"C0C0C0A490C099F8",
 29048 => x"C0C0C0A490C09980",
 29049 => x"C0C0C0A490C09990",
 29050 => x"C0C0C0A490C092C0",
 29051 => x"C0C0C0A490C092F9",
 29052 => x"C0C0C0A490C092A4",
 29053 => x"C0C0C0A490C092B0",
 29054 => x"C0C0C0A490C09299",
 29055 => x"C0C0C0A490C09292",
 29056 => x"C0C0C0A490C09282",
 29057 => x"C0C0C0A490C092F8",
 29058 => x"C0C0C0A490C09280",
 29059 => x"C0C0C0A490C09290",
 29060 => x"C0C0C0A490C082C0",
 29061 => x"C0C0C0A490C082F9",
 29062 => x"C0C0C0A490C082A4",
 29063 => x"C0C0C0A490C082B0",
 29064 => x"C0C0C0A490C08299",
 29065 => x"C0C0C0A490C08292",
 29066 => x"C0C0C0A490C08282",
 29067 => x"C0C0C0A490C082F8",
 29068 => x"C0C0C0A490C08280",
 29069 => x"C0C0C0A490C08290",
 29070 => x"C0C0C0A490C0F8C0",
 29071 => x"C0C0C0A490C0F8F9",
 29072 => x"C0C0C0A490C0F8A4",
 29073 => x"C0C0C0A490C0F8B0",
 29074 => x"C0C0C0A490C0F899",
 29075 => x"C0C0C0A490C0F892",
 29076 => x"C0C0C0A490C0F882",
 29077 => x"C0C0C0A490C0F8F8",
 29078 => x"C0C0C0A490C0F880",
 29079 => x"C0C0C0A490C0F890",
 29080 => x"C0C0C0A490C080C0",
 29081 => x"C0C0C0A490C080F9",
 29082 => x"C0C0C0A490C080A4",
 29083 => x"C0C0C0A490C080B0",
 29084 => x"C0C0C0A490C08099",
 29085 => x"C0C0C0A490C08092",
 29086 => x"C0C0C0A490C08082",
 29087 => x"C0C0C0A490C080F8",
 29088 => x"C0C0C0A490C08080",
 29089 => x"C0C0C0A490C08090",
 29090 => x"C0C0C0A490C090C0",
 29091 => x"C0C0C0A490C090F9",
 29092 => x"C0C0C0A490C090A4",
 29093 => x"C0C0C0A490C090B0",
 29094 => x"C0C0C0A490C09099",
 29095 => x"C0C0C0A490C09092",
 29096 => x"C0C0C0A490C09082",
 29097 => x"C0C0C0A490C090F8",
 29098 => x"C0C0C0A490C09080",
 29099 => x"C0C0C0A490C09090",
 29100 => x"C0C0C0A490F9C0C0",
 29101 => x"C0C0C0A490F9C0F9",
 29102 => x"C0C0C0A490F9C0A4",
 29103 => x"C0C0C0A490F9C0B0",
 29104 => x"C0C0C0A490F9C099",
 29105 => x"C0C0C0A490F9C092",
 29106 => x"C0C0C0A490F9C082",
 29107 => x"C0C0C0A490F9C0F8",
 29108 => x"C0C0C0A490F9C080",
 29109 => x"C0C0C0A490F9C090",
 29110 => x"C0C0C0A490F9F9C0",
 29111 => x"C0C0C0A490F9F9F9",
 29112 => x"C0C0C0A490F9F9A4",
 29113 => x"C0C0C0A490F9F9B0",
 29114 => x"C0C0C0A490F9F999",
 29115 => x"C0C0C0A490F9F992",
 29116 => x"C0C0C0A490F9F982",
 29117 => x"C0C0C0A490F9F9F8",
 29118 => x"C0C0C0A490F9F980",
 29119 => x"C0C0C0A490F9F990",
 29120 => x"C0C0C0A490F9A4C0",
 29121 => x"C0C0C0A490F9A4F9",
 29122 => x"C0C0C0A490F9A4A4",
 29123 => x"C0C0C0A490F9A4B0",
 29124 => x"C0C0C0A490F9A499",
 29125 => x"C0C0C0A490F9A492",
 29126 => x"C0C0C0A490F9A482",
 29127 => x"C0C0C0A490F9A4F8",
 29128 => x"C0C0C0A490F9A480",
 29129 => x"C0C0C0A490F9A490",
 29130 => x"C0C0C0A490F9B0C0",
 29131 => x"C0C0C0A490F9B0F9",
 29132 => x"C0C0C0A490F9B0A4",
 29133 => x"C0C0C0A490F9B0B0",
 29134 => x"C0C0C0A490F9B099",
 29135 => x"C0C0C0A490F9B092",
 29136 => x"C0C0C0A490F9B082",
 29137 => x"C0C0C0A490F9B0F8",
 29138 => x"C0C0C0A490F9B080",
 29139 => x"C0C0C0A490F9B090",
 29140 => x"C0C0C0A490F999C0",
 29141 => x"C0C0C0A490F999F9",
 29142 => x"C0C0C0A490F999A4",
 29143 => x"C0C0C0A490F999B0",
 29144 => x"C0C0C0A490F99999",
 29145 => x"C0C0C0A490F99992",
 29146 => x"C0C0C0A490F99982",
 29147 => x"C0C0C0A490F999F8",
 29148 => x"C0C0C0A490F99980",
 29149 => x"C0C0C0A490F99990",
 29150 => x"C0C0C0A490F992C0",
 29151 => x"C0C0C0A490F992F9",
 29152 => x"C0C0C0A490F992A4",
 29153 => x"C0C0C0A490F992B0",
 29154 => x"C0C0C0A490F99299",
 29155 => x"C0C0C0A490F99292",
 29156 => x"C0C0C0A490F99282",
 29157 => x"C0C0C0A490F992F8",
 29158 => x"C0C0C0A490F99280",
 29159 => x"C0C0C0A490F99290",
 29160 => x"C0C0C0A490F982C0",
 29161 => x"C0C0C0A490F982F9",
 29162 => x"C0C0C0A490F982A4",
 29163 => x"C0C0C0A490F982B0",
 29164 => x"C0C0C0A490F98299",
 29165 => x"C0C0C0A490F98292",
 29166 => x"C0C0C0A490F98282",
 29167 => x"C0C0C0A490F982F8",
 29168 => x"C0C0C0A490F98280",
 29169 => x"C0C0C0A490F98290",
 29170 => x"C0C0C0A490F9F8C0",
 29171 => x"C0C0C0A490F9F8F9",
 29172 => x"C0C0C0A490F9F8A4",
 29173 => x"C0C0C0A490F9F8B0",
 29174 => x"C0C0C0A490F9F899",
 29175 => x"C0C0C0A490F9F892",
 29176 => x"C0C0C0A490F9F882",
 29177 => x"C0C0C0A490F9F8F8",
 29178 => x"C0C0C0A490F9F880",
 29179 => x"C0C0C0A490F9F890",
 29180 => x"C0C0C0A490F980C0",
 29181 => x"C0C0C0A490F980F9",
 29182 => x"C0C0C0A490F980A4",
 29183 => x"C0C0C0A490F980B0",
 29184 => x"C0C0C0A490F98099",
 29185 => x"C0C0C0A490F98092",
 29186 => x"C0C0C0A490F98082",
 29187 => x"C0C0C0A490F980F8",
 29188 => x"C0C0C0A490F98080",
 29189 => x"C0C0C0A490F98090",
 29190 => x"C0C0C0A490F990C0",
 29191 => x"C0C0C0A490F990F9",
 29192 => x"C0C0C0A490F990A4",
 29193 => x"C0C0C0A490F990B0",
 29194 => x"C0C0C0A490F99099",
 29195 => x"C0C0C0A490F99092",
 29196 => x"C0C0C0A490F99082",
 29197 => x"C0C0C0A490F990F8",
 29198 => x"C0C0C0A490F99080",
 29199 => x"C0C0C0A490F99090",
 29200 => x"C0C0C0A490A4C0C0",
 29201 => x"C0C0C0A490A4C0F9",
 29202 => x"C0C0C0A490A4C0A4",
 29203 => x"C0C0C0A490A4C0B0",
 29204 => x"C0C0C0A490A4C099",
 29205 => x"C0C0C0A490A4C092",
 29206 => x"C0C0C0A490A4C082",
 29207 => x"C0C0C0A490A4C0F8",
 29208 => x"C0C0C0A490A4C080",
 29209 => x"C0C0C0A490A4C090",
 29210 => x"C0C0C0A490A4F9C0",
 29211 => x"C0C0C0A490A4F9F9",
 29212 => x"C0C0C0A490A4F9A4",
 29213 => x"C0C0C0A490A4F9B0",
 29214 => x"C0C0C0A490A4F999",
 29215 => x"C0C0C0A490A4F992",
 29216 => x"C0C0C0A490A4F982",
 29217 => x"C0C0C0A490A4F9F8",
 29218 => x"C0C0C0A490A4F980",
 29219 => x"C0C0C0A490A4F990",
 29220 => x"C0C0C0A490A4A4C0",
 29221 => x"C0C0C0A490A4A4F9",
 29222 => x"C0C0C0A490A4A4A4",
 29223 => x"C0C0C0A490A4A4B0",
 29224 => x"C0C0C0A490A4A499",
 29225 => x"C0C0C0A490A4A492",
 29226 => x"C0C0C0A490A4A482",
 29227 => x"C0C0C0A490A4A4F8",
 29228 => x"C0C0C0A490A4A480",
 29229 => x"C0C0C0A490A4A490",
 29230 => x"C0C0C0A490A4B0C0",
 29231 => x"C0C0C0A490A4B0F9",
 29232 => x"C0C0C0A490A4B0A4",
 29233 => x"C0C0C0A490A4B0B0",
 29234 => x"C0C0C0A490A4B099",
 29235 => x"C0C0C0A490A4B092",
 29236 => x"C0C0C0A490A4B082",
 29237 => x"C0C0C0A490A4B0F8",
 29238 => x"C0C0C0A490A4B080",
 29239 => x"C0C0C0A490A4B090",
 29240 => x"C0C0C0A490A499C0",
 29241 => x"C0C0C0A490A499F9",
 29242 => x"C0C0C0A490A499A4",
 29243 => x"C0C0C0A490A499B0",
 29244 => x"C0C0C0A490A49999",
 29245 => x"C0C0C0A490A49992",
 29246 => x"C0C0C0A490A49982",
 29247 => x"C0C0C0A490A499F8",
 29248 => x"C0C0C0A490A49980",
 29249 => x"C0C0C0A490A49990",
 29250 => x"C0C0C0A490A492C0",
 29251 => x"C0C0C0A490A492F9",
 29252 => x"C0C0C0A490A492A4",
 29253 => x"C0C0C0A490A492B0",
 29254 => x"C0C0C0A490A49299",
 29255 => x"C0C0C0A490A49292",
 29256 => x"C0C0C0A490A49282",
 29257 => x"C0C0C0A490A492F8",
 29258 => x"C0C0C0A490A49280",
 29259 => x"C0C0C0A490A49290",
 29260 => x"C0C0C0A490A482C0",
 29261 => x"C0C0C0A490A482F9",
 29262 => x"C0C0C0A490A482A4",
 29263 => x"C0C0C0A490A482B0",
 29264 => x"C0C0C0A490A48299",
 29265 => x"C0C0C0A490A48292",
 29266 => x"C0C0C0A490A48282",
 29267 => x"C0C0C0A490A482F8",
 29268 => x"C0C0C0A490A48280",
 29269 => x"C0C0C0A490A48290",
 29270 => x"C0C0C0A490A4F8C0",
 29271 => x"C0C0C0A490A4F8F9",
 29272 => x"C0C0C0A490A4F8A4",
 29273 => x"C0C0C0A490A4F8B0",
 29274 => x"C0C0C0A490A4F899",
 29275 => x"C0C0C0A490A4F892",
 29276 => x"C0C0C0A490A4F882",
 29277 => x"C0C0C0A490A4F8F8",
 29278 => x"C0C0C0A490A4F880",
 29279 => x"C0C0C0A490A4F890",
 29280 => x"C0C0C0A490A480C0",
 29281 => x"C0C0C0A490A480F9",
 29282 => x"C0C0C0A490A480A4",
 29283 => x"C0C0C0A490A480B0",
 29284 => x"C0C0C0A490A48099",
 29285 => x"C0C0C0A490A48092",
 29286 => x"C0C0C0A490A48082",
 29287 => x"C0C0C0A490A480F8",
 29288 => x"C0C0C0A490A48080",
 29289 => x"C0C0C0A490A48090",
 29290 => x"C0C0C0A490A490C0",
 29291 => x"C0C0C0A490A490F9",
 29292 => x"C0C0C0A490A490A4",
 29293 => x"C0C0C0A490A490B0",
 29294 => x"C0C0C0A490A49099",
 29295 => x"C0C0C0A490A49092",
 29296 => x"C0C0C0A490A49082",
 29297 => x"C0C0C0A490A490F8",
 29298 => x"C0C0C0A490A49080",
 29299 => x"C0C0C0A490A49090",
 29300 => x"C0C0C0A490B0C0C0",
 29301 => x"C0C0C0A490B0C0F9",
 29302 => x"C0C0C0A490B0C0A4",
 29303 => x"C0C0C0A490B0C0B0",
 29304 => x"C0C0C0A490B0C099",
 29305 => x"C0C0C0A490B0C092",
 29306 => x"C0C0C0A490B0C082",
 29307 => x"C0C0C0A490B0C0F8",
 29308 => x"C0C0C0A490B0C080",
 29309 => x"C0C0C0A490B0C090",
 29310 => x"C0C0C0A490B0F9C0",
 29311 => x"C0C0C0A490B0F9F9",
 29312 => x"C0C0C0A490B0F9A4",
 29313 => x"C0C0C0A490B0F9B0",
 29314 => x"C0C0C0A490B0F999",
 29315 => x"C0C0C0A490B0F992",
 29316 => x"C0C0C0A490B0F982",
 29317 => x"C0C0C0A490B0F9F8",
 29318 => x"C0C0C0A490B0F980",
 29319 => x"C0C0C0A490B0F990",
 29320 => x"C0C0C0A490B0A4C0",
 29321 => x"C0C0C0A490B0A4F9",
 29322 => x"C0C0C0A490B0A4A4",
 29323 => x"C0C0C0A490B0A4B0",
 29324 => x"C0C0C0A490B0A499",
 29325 => x"C0C0C0A490B0A492",
 29326 => x"C0C0C0A490B0A482",
 29327 => x"C0C0C0A490B0A4F8",
 29328 => x"C0C0C0A490B0A480",
 29329 => x"C0C0C0A490B0A490",
 29330 => x"C0C0C0A490B0B0C0",
 29331 => x"C0C0C0A490B0B0F9",
 29332 => x"C0C0C0A490B0B0A4",
 29333 => x"C0C0C0A490B0B0B0",
 29334 => x"C0C0C0A490B0B099",
 29335 => x"C0C0C0A490B0B092",
 29336 => x"C0C0C0A490B0B082",
 29337 => x"C0C0C0A490B0B0F8",
 29338 => x"C0C0C0A490B0B080",
 29339 => x"C0C0C0A490B0B090",
 29340 => x"C0C0C0A490B099C0",
 29341 => x"C0C0C0A490B099F9",
 29342 => x"C0C0C0A490B099A4",
 29343 => x"C0C0C0A490B099B0",
 29344 => x"C0C0C0A490B09999",
 29345 => x"C0C0C0A490B09992",
 29346 => x"C0C0C0A490B09982",
 29347 => x"C0C0C0A490B099F8",
 29348 => x"C0C0C0A490B09980",
 29349 => x"C0C0C0A490B09990",
 29350 => x"C0C0C0A490B092C0",
 29351 => x"C0C0C0A490B092F9",
 29352 => x"C0C0C0A490B092A4",
 29353 => x"C0C0C0A490B092B0",
 29354 => x"C0C0C0A490B09299",
 29355 => x"C0C0C0A490B09292",
 29356 => x"C0C0C0A490B09282",
 29357 => x"C0C0C0A490B092F8",
 29358 => x"C0C0C0A490B09280",
 29359 => x"C0C0C0A490B09290",
 29360 => x"C0C0C0A490B082C0",
 29361 => x"C0C0C0A490B082F9",
 29362 => x"C0C0C0A490B082A4",
 29363 => x"C0C0C0A490B082B0",
 29364 => x"C0C0C0A490B08299",
 29365 => x"C0C0C0A490B08292",
 29366 => x"C0C0C0A490B08282",
 29367 => x"C0C0C0A490B082F8",
 29368 => x"C0C0C0A490B08280",
 29369 => x"C0C0C0A490B08290",
 29370 => x"C0C0C0A490B0F8C0",
 29371 => x"C0C0C0A490B0F8F9",
 29372 => x"C0C0C0A490B0F8A4",
 29373 => x"C0C0C0A490B0F8B0",
 29374 => x"C0C0C0A490B0F899",
 29375 => x"C0C0C0A490B0F892",
 29376 => x"C0C0C0A490B0F882",
 29377 => x"C0C0C0A490B0F8F8",
 29378 => x"C0C0C0A490B0F880",
 29379 => x"C0C0C0A490B0F890",
 29380 => x"C0C0C0A490B080C0",
 29381 => x"C0C0C0A490B080F9",
 29382 => x"C0C0C0A490B080A4",
 29383 => x"C0C0C0A490B080B0",
 29384 => x"C0C0C0A490B08099",
 29385 => x"C0C0C0A490B08092",
 29386 => x"C0C0C0A490B08082",
 29387 => x"C0C0C0A490B080F8",
 29388 => x"C0C0C0A490B08080",
 29389 => x"C0C0C0A490B08090",
 29390 => x"C0C0C0A490B090C0",
 29391 => x"C0C0C0A490B090F9",
 29392 => x"C0C0C0A490B090A4",
 29393 => x"C0C0C0A490B090B0",
 29394 => x"C0C0C0A490B09099",
 29395 => x"C0C0C0A490B09092",
 29396 => x"C0C0C0A490B09082",
 29397 => x"C0C0C0A490B090F8",
 29398 => x"C0C0C0A490B09080",
 29399 => x"C0C0C0A490B09090",
 29400 => x"C0C0C0A49099C0C0",
 29401 => x"C0C0C0A49099C0F9",
 29402 => x"C0C0C0A49099C0A4",
 29403 => x"C0C0C0A49099C0B0",
 29404 => x"C0C0C0A49099C099",
 29405 => x"C0C0C0A49099C092",
 29406 => x"C0C0C0A49099C082",
 29407 => x"C0C0C0A49099C0F8",
 29408 => x"C0C0C0A49099C080",
 29409 => x"C0C0C0A49099C090",
 29410 => x"C0C0C0A49099F9C0",
 29411 => x"C0C0C0A49099F9F9",
 29412 => x"C0C0C0A49099F9A4",
 29413 => x"C0C0C0A49099F9B0",
 29414 => x"C0C0C0A49099F999",
 29415 => x"C0C0C0A49099F992",
 29416 => x"C0C0C0A49099F982",
 29417 => x"C0C0C0A49099F9F8",
 29418 => x"C0C0C0A49099F980",
 29419 => x"C0C0C0A49099F990",
 29420 => x"C0C0C0A49099A4C0",
 29421 => x"C0C0C0A49099A4F9",
 29422 => x"C0C0C0A49099A4A4",
 29423 => x"C0C0C0A49099A4B0",
 29424 => x"C0C0C0A49099A499",
 29425 => x"C0C0C0A49099A492",
 29426 => x"C0C0C0A49099A482",
 29427 => x"C0C0C0A49099A4F8",
 29428 => x"C0C0C0A49099A480",
 29429 => x"C0C0C0A49099A490",
 29430 => x"C0C0C0A49099B0C0",
 29431 => x"C0C0C0A49099B0F9",
 29432 => x"C0C0C0A49099B0A4",
 29433 => x"C0C0C0A49099B0B0",
 29434 => x"C0C0C0A49099B099",
 29435 => x"C0C0C0A49099B092",
 29436 => x"C0C0C0A49099B082",
 29437 => x"C0C0C0A49099B0F8",
 29438 => x"C0C0C0A49099B080",
 29439 => x"C0C0C0A49099B090",
 29440 => x"C0C0C0A4909999C0",
 29441 => x"C0C0C0A4909999F9",
 29442 => x"C0C0C0A4909999A4",
 29443 => x"C0C0C0A4909999B0",
 29444 => x"C0C0C0A490999999",
 29445 => x"C0C0C0A490999992",
 29446 => x"C0C0C0A490999982",
 29447 => x"C0C0C0A4909999F8",
 29448 => x"C0C0C0A490999980",
 29449 => x"C0C0C0A490999990",
 29450 => x"C0C0C0A4909992C0",
 29451 => x"C0C0C0A4909992F9",
 29452 => x"C0C0C0A4909992A4",
 29453 => x"C0C0C0A4909992B0",
 29454 => x"C0C0C0A490999299",
 29455 => x"C0C0C0A490999292",
 29456 => x"C0C0C0A490999282",
 29457 => x"C0C0C0A4909992F8",
 29458 => x"C0C0C0A490999280",
 29459 => x"C0C0C0A490999290",
 29460 => x"C0C0C0A4909982C0",
 29461 => x"C0C0C0A4909982F9",
 29462 => x"C0C0C0A4909982A4",
 29463 => x"C0C0C0A4909982B0",
 29464 => x"C0C0C0A490998299",
 29465 => x"C0C0C0A490998292",
 29466 => x"C0C0C0A490998282",
 29467 => x"C0C0C0A4909982F8",
 29468 => x"C0C0C0A490998280",
 29469 => x"C0C0C0A490998290",
 29470 => x"C0C0C0A49099F8C0",
 29471 => x"C0C0C0A49099F8F9",
 29472 => x"C0C0C0A49099F8A4",
 29473 => x"C0C0C0A49099F8B0",
 29474 => x"C0C0C0A49099F899",
 29475 => x"C0C0C0A49099F892",
 29476 => x"C0C0C0A49099F882",
 29477 => x"C0C0C0A49099F8F8",
 29478 => x"C0C0C0A49099F880",
 29479 => x"C0C0C0A49099F890",
 29480 => x"C0C0C0A4909980C0",
 29481 => x"C0C0C0A4909980F9",
 29482 => x"C0C0C0A4909980A4",
 29483 => x"C0C0C0A4909980B0",
 29484 => x"C0C0C0A490998099",
 29485 => x"C0C0C0A490998092",
 29486 => x"C0C0C0A490998082",
 29487 => x"C0C0C0A4909980F8",
 29488 => x"C0C0C0A490998080",
 29489 => x"C0C0C0A490998090",
 29490 => x"C0C0C0A4909990C0",
 29491 => x"C0C0C0A4909990F9",
 29492 => x"C0C0C0A4909990A4",
 29493 => x"C0C0C0A4909990B0",
 29494 => x"C0C0C0A490999099",
 29495 => x"C0C0C0A490999092",
 29496 => x"C0C0C0A490999082",
 29497 => x"C0C0C0A4909990F8",
 29498 => x"C0C0C0A490999080",
 29499 => x"C0C0C0A490999090",
 29500 => x"C0C0C0A49092C0C0",
 29501 => x"C0C0C0A49092C0F9",
 29502 => x"C0C0C0A49092C0A4",
 29503 => x"C0C0C0A49092C0B0",
 29504 => x"C0C0C0A49092C099",
 29505 => x"C0C0C0A49092C092",
 29506 => x"C0C0C0A49092C082",
 29507 => x"C0C0C0A49092C0F8",
 29508 => x"C0C0C0A49092C080",
 29509 => x"C0C0C0A49092C090",
 29510 => x"C0C0C0A49092F9C0",
 29511 => x"C0C0C0A49092F9F9",
 29512 => x"C0C0C0A49092F9A4",
 29513 => x"C0C0C0A49092F9B0",
 29514 => x"C0C0C0A49092F999",
 29515 => x"C0C0C0A49092F992",
 29516 => x"C0C0C0A49092F982",
 29517 => x"C0C0C0A49092F9F8",
 29518 => x"C0C0C0A49092F980",
 29519 => x"C0C0C0A49092F990",
 29520 => x"C0C0C0A49092A4C0",
 29521 => x"C0C0C0A49092A4F9",
 29522 => x"C0C0C0A49092A4A4",
 29523 => x"C0C0C0A49092A4B0",
 29524 => x"C0C0C0A49092A499",
 29525 => x"C0C0C0A49092A492",
 29526 => x"C0C0C0A49092A482",
 29527 => x"C0C0C0A49092A4F8",
 29528 => x"C0C0C0A49092A480",
 29529 => x"C0C0C0A49092A490",
 29530 => x"C0C0C0A49092B0C0",
 29531 => x"C0C0C0A49092B0F9",
 29532 => x"C0C0C0A49092B0A4",
 29533 => x"C0C0C0A49092B0B0",
 29534 => x"C0C0C0A49092B099",
 29535 => x"C0C0C0A49092B092",
 29536 => x"C0C0C0A49092B082",
 29537 => x"C0C0C0A49092B0F8",
 29538 => x"C0C0C0A49092B080",
 29539 => x"C0C0C0A49092B090",
 29540 => x"C0C0C0A4909299C0",
 29541 => x"C0C0C0A4909299F9",
 29542 => x"C0C0C0A4909299A4",
 29543 => x"C0C0C0A4909299B0",
 29544 => x"C0C0C0A490929999",
 29545 => x"C0C0C0A490929992",
 29546 => x"C0C0C0A490929982",
 29547 => x"C0C0C0A4909299F8",
 29548 => x"C0C0C0A490929980",
 29549 => x"C0C0C0A490929990",
 29550 => x"C0C0C0A4909292C0",
 29551 => x"C0C0C0A4909292F9",
 29552 => x"C0C0C0A4909292A4",
 29553 => x"C0C0C0A4909292B0",
 29554 => x"C0C0C0A490929299",
 29555 => x"C0C0C0A490929292",
 29556 => x"C0C0C0A490929282",
 29557 => x"C0C0C0A4909292F8",
 29558 => x"C0C0C0A490929280",
 29559 => x"C0C0C0A490929290",
 29560 => x"C0C0C0A4909282C0",
 29561 => x"C0C0C0A4909282F9",
 29562 => x"C0C0C0A4909282A4",
 29563 => x"C0C0C0A4909282B0",
 29564 => x"C0C0C0A490928299",
 29565 => x"C0C0C0A490928292",
 29566 => x"C0C0C0A490928282",
 29567 => x"C0C0C0A4909282F8",
 29568 => x"C0C0C0A490928280",
 29569 => x"C0C0C0A490928290",
 29570 => x"C0C0C0A49092F8C0",
 29571 => x"C0C0C0A49092F8F9",
 29572 => x"C0C0C0A49092F8A4",
 29573 => x"C0C0C0A49092F8B0",
 29574 => x"C0C0C0A49092F899",
 29575 => x"C0C0C0A49092F892",
 29576 => x"C0C0C0A49092F882",
 29577 => x"C0C0C0A49092F8F8",
 29578 => x"C0C0C0A49092F880",
 29579 => x"C0C0C0A49092F890",
 29580 => x"C0C0C0A4909280C0",
 29581 => x"C0C0C0A4909280F9",
 29582 => x"C0C0C0A4909280A4",
 29583 => x"C0C0C0A4909280B0",
 29584 => x"C0C0C0A490928099",
 29585 => x"C0C0C0A490928092",
 29586 => x"C0C0C0A490928082",
 29587 => x"C0C0C0A4909280F8",
 29588 => x"C0C0C0A490928080",
 29589 => x"C0C0C0A490928090",
 29590 => x"C0C0C0A4909290C0",
 29591 => x"C0C0C0A4909290F9",
 29592 => x"C0C0C0A4909290A4",
 29593 => x"C0C0C0A4909290B0",
 29594 => x"C0C0C0A490929099",
 29595 => x"C0C0C0A490929092",
 29596 => x"C0C0C0A490929082",
 29597 => x"C0C0C0A4909290F8",
 29598 => x"C0C0C0A490929080",
 29599 => x"C0C0C0A490929090",
 29600 => x"C0C0C0A49082C0C0",
 29601 => x"C0C0C0A49082C0F9",
 29602 => x"C0C0C0A49082C0A4",
 29603 => x"C0C0C0A49082C0B0",
 29604 => x"C0C0C0A49082C099",
 29605 => x"C0C0C0A49082C092",
 29606 => x"C0C0C0A49082C082",
 29607 => x"C0C0C0A49082C0F8",
 29608 => x"C0C0C0A49082C080",
 29609 => x"C0C0C0A49082C090",
 29610 => x"C0C0C0A49082F9C0",
 29611 => x"C0C0C0A49082F9F9",
 29612 => x"C0C0C0A49082F9A4",
 29613 => x"C0C0C0A49082F9B0",
 29614 => x"C0C0C0A49082F999",
 29615 => x"C0C0C0A49082F992",
 29616 => x"C0C0C0A49082F982",
 29617 => x"C0C0C0A49082F9F8",
 29618 => x"C0C0C0A49082F980",
 29619 => x"C0C0C0A49082F990",
 29620 => x"C0C0C0A49082A4C0",
 29621 => x"C0C0C0A49082A4F9",
 29622 => x"C0C0C0A49082A4A4",
 29623 => x"C0C0C0A49082A4B0",
 29624 => x"C0C0C0A49082A499",
 29625 => x"C0C0C0A49082A492",
 29626 => x"C0C0C0A49082A482",
 29627 => x"C0C0C0A49082A4F8",
 29628 => x"C0C0C0A49082A480",
 29629 => x"C0C0C0A49082A490",
 29630 => x"C0C0C0A49082B0C0",
 29631 => x"C0C0C0A49082B0F9",
 29632 => x"C0C0C0A49082B0A4",
 29633 => x"C0C0C0A49082B0B0",
 29634 => x"C0C0C0A49082B099",
 29635 => x"C0C0C0A49082B092",
 29636 => x"C0C0C0A49082B082",
 29637 => x"C0C0C0A49082B0F8",
 29638 => x"C0C0C0A49082B080",
 29639 => x"C0C0C0A49082B090",
 29640 => x"C0C0C0A4908299C0",
 29641 => x"C0C0C0A4908299F9",
 29642 => x"C0C0C0A4908299A4",
 29643 => x"C0C0C0A4908299B0",
 29644 => x"C0C0C0A490829999",
 29645 => x"C0C0C0A490829992",
 29646 => x"C0C0C0A490829982",
 29647 => x"C0C0C0A4908299F8",
 29648 => x"C0C0C0A490829980",
 29649 => x"C0C0C0A490829990",
 29650 => x"C0C0C0A4908292C0",
 29651 => x"C0C0C0A4908292F9",
 29652 => x"C0C0C0A4908292A4",
 29653 => x"C0C0C0A4908292B0",
 29654 => x"C0C0C0A490829299",
 29655 => x"C0C0C0A490829292",
 29656 => x"C0C0C0A490829282",
 29657 => x"C0C0C0A4908292F8",
 29658 => x"C0C0C0A490829280",
 29659 => x"C0C0C0A490829290",
 29660 => x"C0C0C0A4908282C0",
 29661 => x"C0C0C0A4908282F9",
 29662 => x"C0C0C0A4908282A4",
 29663 => x"C0C0C0A4908282B0",
 29664 => x"C0C0C0A490828299",
 29665 => x"C0C0C0A490828292",
 29666 => x"C0C0C0A490828282",
 29667 => x"C0C0C0A4908282F8",
 29668 => x"C0C0C0A490828280",
 29669 => x"C0C0C0A490828290",
 29670 => x"C0C0C0A49082F8C0",
 29671 => x"C0C0C0A49082F8F9",
 29672 => x"C0C0C0A49082F8A4",
 29673 => x"C0C0C0A49082F8B0",
 29674 => x"C0C0C0A49082F899",
 29675 => x"C0C0C0A49082F892",
 29676 => x"C0C0C0A49082F882",
 29677 => x"C0C0C0A49082F8F8",
 29678 => x"C0C0C0A49082F880",
 29679 => x"C0C0C0A49082F890",
 29680 => x"C0C0C0A4908280C0",
 29681 => x"C0C0C0A4908280F9",
 29682 => x"C0C0C0A4908280A4",
 29683 => x"C0C0C0A4908280B0",
 29684 => x"C0C0C0A490828099",
 29685 => x"C0C0C0A490828092",
 29686 => x"C0C0C0A490828082",
 29687 => x"C0C0C0A4908280F8",
 29688 => x"C0C0C0A490828080",
 29689 => x"C0C0C0A490828090",
 29690 => x"C0C0C0A4908290C0",
 29691 => x"C0C0C0A4908290F9",
 29692 => x"C0C0C0A4908290A4",
 29693 => x"C0C0C0A4908290B0",
 29694 => x"C0C0C0A490829099",
 29695 => x"C0C0C0A490829092",
 29696 => x"C0C0C0A490829082",
 29697 => x"C0C0C0A4908290F8",
 29698 => x"C0C0C0A490829080",
 29699 => x"C0C0C0A490829090",
 29700 => x"C0C0C0A490F8C0C0",
 29701 => x"C0C0C0A490F8C0F9",
 29702 => x"C0C0C0A490F8C0A4",
 29703 => x"C0C0C0A490F8C0B0",
 29704 => x"C0C0C0A490F8C099",
 29705 => x"C0C0C0A490F8C092",
 29706 => x"C0C0C0A490F8C082",
 29707 => x"C0C0C0A490F8C0F8",
 29708 => x"C0C0C0A490F8C080",
 29709 => x"C0C0C0A490F8C090",
 29710 => x"C0C0C0A490F8F9C0",
 29711 => x"C0C0C0A490F8F9F9",
 29712 => x"C0C0C0A490F8F9A4",
 29713 => x"C0C0C0A490F8F9B0",
 29714 => x"C0C0C0A490F8F999",
 29715 => x"C0C0C0A490F8F992",
 29716 => x"C0C0C0A490F8F982",
 29717 => x"C0C0C0A490F8F9F8",
 29718 => x"C0C0C0A490F8F980",
 29719 => x"C0C0C0A490F8F990",
 29720 => x"C0C0C0A490F8A4C0",
 29721 => x"C0C0C0A490F8A4F9",
 29722 => x"C0C0C0A490F8A4A4",
 29723 => x"C0C0C0A490F8A4B0",
 29724 => x"C0C0C0A490F8A499",
 29725 => x"C0C0C0A490F8A492",
 29726 => x"C0C0C0A490F8A482",
 29727 => x"C0C0C0A490F8A4F8",
 29728 => x"C0C0C0A490F8A480",
 29729 => x"C0C0C0A490F8A490",
 29730 => x"C0C0C0A490F8B0C0",
 29731 => x"C0C0C0A490F8B0F9",
 29732 => x"C0C0C0A490F8B0A4",
 29733 => x"C0C0C0A490F8B0B0",
 29734 => x"C0C0C0A490F8B099",
 29735 => x"C0C0C0A490F8B092",
 29736 => x"C0C0C0A490F8B082",
 29737 => x"C0C0C0A490F8B0F8",
 29738 => x"C0C0C0A490F8B080",
 29739 => x"C0C0C0A490F8B090",
 29740 => x"C0C0C0A490F899C0",
 29741 => x"C0C0C0A490F899F9",
 29742 => x"C0C0C0A490F899A4",
 29743 => x"C0C0C0A490F899B0",
 29744 => x"C0C0C0A490F89999",
 29745 => x"C0C0C0A490F89992",
 29746 => x"C0C0C0A490F89982",
 29747 => x"C0C0C0A490F899F8",
 29748 => x"C0C0C0A490F89980",
 29749 => x"C0C0C0A490F89990",
 29750 => x"C0C0C0A490F892C0",
 29751 => x"C0C0C0A490F892F9",
 29752 => x"C0C0C0A490F892A4",
 29753 => x"C0C0C0A490F892B0",
 29754 => x"C0C0C0A490F89299",
 29755 => x"C0C0C0A490F89292",
 29756 => x"C0C0C0A490F89282",
 29757 => x"C0C0C0A490F892F8",
 29758 => x"C0C0C0A490F89280",
 29759 => x"C0C0C0A490F89290",
 29760 => x"C0C0C0A490F882C0",
 29761 => x"C0C0C0A490F882F9",
 29762 => x"C0C0C0A490F882A4",
 29763 => x"C0C0C0A490F882B0",
 29764 => x"C0C0C0A490F88299",
 29765 => x"C0C0C0A490F88292",
 29766 => x"C0C0C0A490F88282",
 29767 => x"C0C0C0A490F882F8",
 29768 => x"C0C0C0A490F88280",
 29769 => x"C0C0C0A490F88290",
 29770 => x"C0C0C0A490F8F8C0",
 29771 => x"C0C0C0A490F8F8F9",
 29772 => x"C0C0C0A490F8F8A4",
 29773 => x"C0C0C0A490F8F8B0",
 29774 => x"C0C0C0A490F8F899",
 29775 => x"C0C0C0A490F8F892",
 29776 => x"C0C0C0A490F8F882",
 29777 => x"C0C0C0A490F8F8F8",
 29778 => x"C0C0C0A490F8F880",
 29779 => x"C0C0C0A490F8F890",
 29780 => x"C0C0C0A490F880C0",
 29781 => x"C0C0C0A490F880F9",
 29782 => x"C0C0C0A490F880A4",
 29783 => x"C0C0C0A490F880B0",
 29784 => x"C0C0C0A490F88099",
 29785 => x"C0C0C0A490F88092",
 29786 => x"C0C0C0A490F88082",
 29787 => x"C0C0C0A490F880F8",
 29788 => x"C0C0C0A490F88080",
 29789 => x"C0C0C0A490F88090",
 29790 => x"C0C0C0A490F890C0",
 29791 => x"C0C0C0A490F890F9",
 29792 => x"C0C0C0A490F890A4",
 29793 => x"C0C0C0A490F890B0",
 29794 => x"C0C0C0A490F89099",
 29795 => x"C0C0C0A490F89092",
 29796 => x"C0C0C0A490F89082",
 29797 => x"C0C0C0A490F890F8",
 29798 => x"C0C0C0A490F89080",
 29799 => x"C0C0C0A490F89090",
 29800 => x"C0C0C0A49080C0C0",
 29801 => x"C0C0C0A49080C0F9",
 29802 => x"C0C0C0A49080C0A4",
 29803 => x"C0C0C0A49080C0B0",
 29804 => x"C0C0C0A49080C099",
 29805 => x"C0C0C0A49080C092",
 29806 => x"C0C0C0A49080C082",
 29807 => x"C0C0C0A49080C0F8",
 29808 => x"C0C0C0A49080C080",
 29809 => x"C0C0C0A49080C090",
 29810 => x"C0C0C0A49080F9C0",
 29811 => x"C0C0C0A49080F9F9",
 29812 => x"C0C0C0A49080F9A4",
 29813 => x"C0C0C0A49080F9B0",
 29814 => x"C0C0C0A49080F999",
 29815 => x"C0C0C0A49080F992",
 29816 => x"C0C0C0A49080F982",
 29817 => x"C0C0C0A49080F9F8",
 29818 => x"C0C0C0A49080F980",
 29819 => x"C0C0C0A49080F990",
 29820 => x"C0C0C0A49080A4C0",
 29821 => x"C0C0C0A49080A4F9",
 29822 => x"C0C0C0A49080A4A4",
 29823 => x"C0C0C0A49080A4B0",
 29824 => x"C0C0C0A49080A499",
 29825 => x"C0C0C0A49080A492",
 29826 => x"C0C0C0A49080A482",
 29827 => x"C0C0C0A49080A4F8",
 29828 => x"C0C0C0A49080A480",
 29829 => x"C0C0C0A49080A490",
 29830 => x"C0C0C0A49080B0C0",
 29831 => x"C0C0C0A49080B0F9",
 29832 => x"C0C0C0A49080B0A4",
 29833 => x"C0C0C0A49080B0B0",
 29834 => x"C0C0C0A49080B099",
 29835 => x"C0C0C0A49080B092",
 29836 => x"C0C0C0A49080B082",
 29837 => x"C0C0C0A49080B0F8",
 29838 => x"C0C0C0A49080B080",
 29839 => x"C0C0C0A49080B090",
 29840 => x"C0C0C0A4908099C0",
 29841 => x"C0C0C0A4908099F9",
 29842 => x"C0C0C0A4908099A4",
 29843 => x"C0C0C0A4908099B0",
 29844 => x"C0C0C0A490809999",
 29845 => x"C0C0C0A490809992",
 29846 => x"C0C0C0A490809982",
 29847 => x"C0C0C0A4908099F8",
 29848 => x"C0C0C0A490809980",
 29849 => x"C0C0C0A490809990",
 29850 => x"C0C0C0A4908092C0",
 29851 => x"C0C0C0A4908092F9",
 29852 => x"C0C0C0A4908092A4",
 29853 => x"C0C0C0A4908092B0",
 29854 => x"C0C0C0A490809299",
 29855 => x"C0C0C0A490809292",
 29856 => x"C0C0C0A490809282",
 29857 => x"C0C0C0A4908092F8",
 29858 => x"C0C0C0A490809280",
 29859 => x"C0C0C0A490809290",
 29860 => x"C0C0C0A4908082C0",
 29861 => x"C0C0C0A4908082F9",
 29862 => x"C0C0C0A4908082A4",
 29863 => x"C0C0C0A4908082B0",
 29864 => x"C0C0C0A490808299",
 29865 => x"C0C0C0A490808292",
 29866 => x"C0C0C0A490808282",
 29867 => x"C0C0C0A4908082F8",
 29868 => x"C0C0C0A490808280",
 29869 => x"C0C0C0A490808290",
 29870 => x"C0C0C0A49080F8C0",
 29871 => x"C0C0C0A49080F8F9",
 29872 => x"C0C0C0A49080F8A4",
 29873 => x"C0C0C0A49080F8B0",
 29874 => x"C0C0C0A49080F899",
 29875 => x"C0C0C0A49080F892",
 29876 => x"C0C0C0A49080F882",
 29877 => x"C0C0C0A49080F8F8",
 29878 => x"C0C0C0A49080F880",
 29879 => x"C0C0C0A49080F890",
 29880 => x"C0C0C0A4908080C0",
 29881 => x"C0C0C0A4908080F9",
 29882 => x"C0C0C0A4908080A4",
 29883 => x"C0C0C0A4908080B0",
 29884 => x"C0C0C0A490808099",
 29885 => x"C0C0C0A490808092",
 29886 => x"C0C0C0A490808082",
 29887 => x"C0C0C0A4908080F8",
 29888 => x"C0C0C0A490808080",
 29889 => x"C0C0C0A490808090",
 29890 => x"C0C0C0A4908090C0",
 29891 => x"C0C0C0A4908090F9",
 29892 => x"C0C0C0A4908090A4",
 29893 => x"C0C0C0A4908090B0",
 29894 => x"C0C0C0A490809099",
 29895 => x"C0C0C0A490809092",
 29896 => x"C0C0C0A490809082",
 29897 => x"C0C0C0A4908090F8",
 29898 => x"C0C0C0A490809080",
 29899 => x"C0C0C0A490809090",
 29900 => x"C0C0C0A49090C0C0",
 29901 => x"C0C0C0A49090C0F9",
 29902 => x"C0C0C0A49090C0A4",
 29903 => x"C0C0C0A49090C0B0",
 29904 => x"C0C0C0A49090C099",
 29905 => x"C0C0C0A49090C092",
 29906 => x"C0C0C0A49090C082",
 29907 => x"C0C0C0A49090C0F8",
 29908 => x"C0C0C0A49090C080",
 29909 => x"C0C0C0A49090C090",
 29910 => x"C0C0C0A49090F9C0",
 29911 => x"C0C0C0A49090F9F9",
 29912 => x"C0C0C0A49090F9A4",
 29913 => x"C0C0C0A49090F9B0",
 29914 => x"C0C0C0A49090F999",
 29915 => x"C0C0C0A49090F992",
 29916 => x"C0C0C0A49090F982",
 29917 => x"C0C0C0A49090F9F8",
 29918 => x"C0C0C0A49090F980",
 29919 => x"C0C0C0A49090F990",
 29920 => x"C0C0C0A49090A4C0",
 29921 => x"C0C0C0A49090A4F9",
 29922 => x"C0C0C0A49090A4A4",
 29923 => x"C0C0C0A49090A4B0",
 29924 => x"C0C0C0A49090A499",
 29925 => x"C0C0C0A49090A492",
 29926 => x"C0C0C0A49090A482",
 29927 => x"C0C0C0A49090A4F8",
 29928 => x"C0C0C0A49090A480",
 29929 => x"C0C0C0A49090A490",
 29930 => x"C0C0C0A49090B0C0",
 29931 => x"C0C0C0A49090B0F9",
 29932 => x"C0C0C0A49090B0A4",
 29933 => x"C0C0C0A49090B0B0",
 29934 => x"C0C0C0A49090B099",
 29935 => x"C0C0C0A49090B092",
 29936 => x"C0C0C0A49090B082",
 29937 => x"C0C0C0A49090B0F8",
 29938 => x"C0C0C0A49090B080",
 29939 => x"C0C0C0A49090B090",
 29940 => x"C0C0C0A4909099C0",
 29941 => x"C0C0C0A4909099F9",
 29942 => x"C0C0C0A4909099A4",
 29943 => x"C0C0C0A4909099B0",
 29944 => x"C0C0C0A490909999",
 29945 => x"C0C0C0A490909992",
 29946 => x"C0C0C0A490909982",
 29947 => x"C0C0C0A4909099F8",
 29948 => x"C0C0C0A490909980",
 29949 => x"C0C0C0A490909990",
 29950 => x"C0C0C0A4909092C0",
 29951 => x"C0C0C0A4909092F9",
 29952 => x"C0C0C0A4909092A4",
 29953 => x"C0C0C0A4909092B0",
 29954 => x"C0C0C0A490909299",
 29955 => x"C0C0C0A490909292",
 29956 => x"C0C0C0A490909282",
 29957 => x"C0C0C0A4909092F8",
 29958 => x"C0C0C0A490909280",
 29959 => x"C0C0C0A490909290",
 29960 => x"C0C0C0A4909082C0",
 29961 => x"C0C0C0A4909082F9",
 29962 => x"C0C0C0A4909082A4",
 29963 => x"C0C0C0A4909082B0",
 29964 => x"C0C0C0A490908299",
 29965 => x"C0C0C0A490908292",
 29966 => x"C0C0C0A490908282",
 29967 => x"C0C0C0A4909082F8",
 29968 => x"C0C0C0A490908280",
 29969 => x"C0C0C0A490908290",
 29970 => x"C0C0C0A49090F8C0",
 29971 => x"C0C0C0A49090F8F9",
 29972 => x"C0C0C0A49090F8A4",
 29973 => x"C0C0C0A49090F8B0",
 29974 => x"C0C0C0A49090F899",
 29975 => x"C0C0C0A49090F892",
 29976 => x"C0C0C0A49090F882",
 29977 => x"C0C0C0A49090F8F8",
 29978 => x"C0C0C0A49090F880",
 29979 => x"C0C0C0A49090F890",
 29980 => x"C0C0C0A4909080C0",
 29981 => x"C0C0C0A4909080F9",
 29982 => x"C0C0C0A4909080A4",
 29983 => x"C0C0C0A4909080B0",
 29984 => x"C0C0C0A490908099",
 29985 => x"C0C0C0A490908092",
 29986 => x"C0C0C0A490908082",
 29987 => x"C0C0C0A4909080F8",
 29988 => x"C0C0C0A490908080",
 29989 => x"C0C0C0A490908090",
 29990 => x"C0C0C0A4909090C0",
 29991 => x"C0C0C0A4909090F9",
 29992 => x"C0C0C0A4909090A4",
 29993 => x"C0C0C0A4909090B0",
 29994 => x"C0C0C0A490909099",
 29995 => x"C0C0C0A490909092",
 29996 => x"C0C0C0A490909082",
 29997 => x"C0C0C0A4909090F8",
 29998 => x"C0C0C0A490909080",
 29999 => x"C0C0C0A490909090",
 30000 => x"C0C0C0B0C0C0C0C0",
 30001 => x"C0C0C0B0C0C0C0F9",
 30002 => x"C0C0C0B0C0C0C0A4",
 30003 => x"C0C0C0B0C0C0C0B0",
 30004 => x"C0C0C0B0C0C0C099",
 30005 => x"C0C0C0B0C0C0C092",
 30006 => x"C0C0C0B0C0C0C082",
 30007 => x"C0C0C0B0C0C0C0F8",
 30008 => x"C0C0C0B0C0C0C080",
 30009 => x"C0C0C0B0C0C0C090",
 30010 => x"C0C0C0B0C0C0F9C0",
 30011 => x"C0C0C0B0C0C0F9F9",
 30012 => x"C0C0C0B0C0C0F9A4",
 30013 => x"C0C0C0B0C0C0F9B0",
 30014 => x"C0C0C0B0C0C0F999",
 30015 => x"C0C0C0B0C0C0F992",
 30016 => x"C0C0C0B0C0C0F982",
 30017 => x"C0C0C0B0C0C0F9F8",
 30018 => x"C0C0C0B0C0C0F980",
 30019 => x"C0C0C0B0C0C0F990",
 30020 => x"C0C0C0B0C0C0A4C0",
 30021 => x"C0C0C0B0C0C0A4F9",
 30022 => x"C0C0C0B0C0C0A4A4",
 30023 => x"C0C0C0B0C0C0A4B0",
 30024 => x"C0C0C0B0C0C0A499",
 30025 => x"C0C0C0B0C0C0A492",
 30026 => x"C0C0C0B0C0C0A482",
 30027 => x"C0C0C0B0C0C0A4F8",
 30028 => x"C0C0C0B0C0C0A480",
 30029 => x"C0C0C0B0C0C0A490",
 30030 => x"C0C0C0B0C0C0B0C0",
 30031 => x"C0C0C0B0C0C0B0F9",
 30032 => x"C0C0C0B0C0C0B0A4",
 30033 => x"C0C0C0B0C0C0B0B0",
 30034 => x"C0C0C0B0C0C0B099",
 30035 => x"C0C0C0B0C0C0B092",
 30036 => x"C0C0C0B0C0C0B082",
 30037 => x"C0C0C0B0C0C0B0F8",
 30038 => x"C0C0C0B0C0C0B080",
 30039 => x"C0C0C0B0C0C0B090",
 30040 => x"C0C0C0B0C0C099C0",
 30041 => x"C0C0C0B0C0C099F9",
 30042 => x"C0C0C0B0C0C099A4",
 30043 => x"C0C0C0B0C0C099B0",
 30044 => x"C0C0C0B0C0C09999",
 30045 => x"C0C0C0B0C0C09992",
 30046 => x"C0C0C0B0C0C09982",
 30047 => x"C0C0C0B0C0C099F8",
 30048 => x"C0C0C0B0C0C09980",
 30049 => x"C0C0C0B0C0C09990",
 30050 => x"C0C0C0B0C0C092C0",
 30051 => x"C0C0C0B0C0C092F9",
 30052 => x"C0C0C0B0C0C092A4",
 30053 => x"C0C0C0B0C0C092B0",
 30054 => x"C0C0C0B0C0C09299",
 30055 => x"C0C0C0B0C0C09292",
 30056 => x"C0C0C0B0C0C09282",
 30057 => x"C0C0C0B0C0C092F8",
 30058 => x"C0C0C0B0C0C09280",
 30059 => x"C0C0C0B0C0C09290",
 30060 => x"C0C0C0B0C0C082C0",
 30061 => x"C0C0C0B0C0C082F9",
 30062 => x"C0C0C0B0C0C082A4",
 30063 => x"C0C0C0B0C0C082B0",
 30064 => x"C0C0C0B0C0C08299",
 30065 => x"C0C0C0B0C0C08292",
 30066 => x"C0C0C0B0C0C08282",
 30067 => x"C0C0C0B0C0C082F8",
 30068 => x"C0C0C0B0C0C08280",
 30069 => x"C0C0C0B0C0C08290",
 30070 => x"C0C0C0B0C0C0F8C0",
 30071 => x"C0C0C0B0C0C0F8F9",
 30072 => x"C0C0C0B0C0C0F8A4",
 30073 => x"C0C0C0B0C0C0F8B0",
 30074 => x"C0C0C0B0C0C0F899",
 30075 => x"C0C0C0B0C0C0F892",
 30076 => x"C0C0C0B0C0C0F882",
 30077 => x"C0C0C0B0C0C0F8F8",
 30078 => x"C0C0C0B0C0C0F880",
 30079 => x"C0C0C0B0C0C0F890",
 30080 => x"C0C0C0B0C0C080C0",
 30081 => x"C0C0C0B0C0C080F9",
 30082 => x"C0C0C0B0C0C080A4",
 30083 => x"C0C0C0B0C0C080B0",
 30084 => x"C0C0C0B0C0C08099",
 30085 => x"C0C0C0B0C0C08092",
 30086 => x"C0C0C0B0C0C08082",
 30087 => x"C0C0C0B0C0C080F8",
 30088 => x"C0C0C0B0C0C08080",
 30089 => x"C0C0C0B0C0C08090",
 30090 => x"C0C0C0B0C0C090C0",
 30091 => x"C0C0C0B0C0C090F9",
 30092 => x"C0C0C0B0C0C090A4",
 30093 => x"C0C0C0B0C0C090B0",
 30094 => x"C0C0C0B0C0C09099",
 30095 => x"C0C0C0B0C0C09092",
 30096 => x"C0C0C0B0C0C09082",
 30097 => x"C0C0C0B0C0C090F8",
 30098 => x"C0C0C0B0C0C09080",
 30099 => x"C0C0C0B0C0C09090",
 30100 => x"C0C0C0B0C0F9C0C0",
 30101 => x"C0C0C0B0C0F9C0F9",
 30102 => x"C0C0C0B0C0F9C0A4",
 30103 => x"C0C0C0B0C0F9C0B0",
 30104 => x"C0C0C0B0C0F9C099",
 30105 => x"C0C0C0B0C0F9C092",
 30106 => x"C0C0C0B0C0F9C082",
 30107 => x"C0C0C0B0C0F9C0F8",
 30108 => x"C0C0C0B0C0F9C080",
 30109 => x"C0C0C0B0C0F9C090",
 30110 => x"C0C0C0B0C0F9F9C0",
 30111 => x"C0C0C0B0C0F9F9F9",
 30112 => x"C0C0C0B0C0F9F9A4",
 30113 => x"C0C0C0B0C0F9F9B0",
 30114 => x"C0C0C0B0C0F9F999",
 30115 => x"C0C0C0B0C0F9F992",
 30116 => x"C0C0C0B0C0F9F982",
 30117 => x"C0C0C0B0C0F9F9F8",
 30118 => x"C0C0C0B0C0F9F980",
 30119 => x"C0C0C0B0C0F9F990",
 30120 => x"C0C0C0B0C0F9A4C0",
 30121 => x"C0C0C0B0C0F9A4F9",
 30122 => x"C0C0C0B0C0F9A4A4",
 30123 => x"C0C0C0B0C0F9A4B0",
 30124 => x"C0C0C0B0C0F9A499",
 30125 => x"C0C0C0B0C0F9A492",
 30126 => x"C0C0C0B0C0F9A482",
 30127 => x"C0C0C0B0C0F9A4F8",
 30128 => x"C0C0C0B0C0F9A480",
 30129 => x"C0C0C0B0C0F9A490",
 30130 => x"C0C0C0B0C0F9B0C0",
 30131 => x"C0C0C0B0C0F9B0F9",
 30132 => x"C0C0C0B0C0F9B0A4",
 30133 => x"C0C0C0B0C0F9B0B0",
 30134 => x"C0C0C0B0C0F9B099",
 30135 => x"C0C0C0B0C0F9B092",
 30136 => x"C0C0C0B0C0F9B082",
 30137 => x"C0C0C0B0C0F9B0F8",
 30138 => x"C0C0C0B0C0F9B080",
 30139 => x"C0C0C0B0C0F9B090",
 30140 => x"C0C0C0B0C0F999C0",
 30141 => x"C0C0C0B0C0F999F9",
 30142 => x"C0C0C0B0C0F999A4",
 30143 => x"C0C0C0B0C0F999B0",
 30144 => x"C0C0C0B0C0F99999",
 30145 => x"C0C0C0B0C0F99992",
 30146 => x"C0C0C0B0C0F99982",
 30147 => x"C0C0C0B0C0F999F8",
 30148 => x"C0C0C0B0C0F99980",
 30149 => x"C0C0C0B0C0F99990",
 30150 => x"C0C0C0B0C0F992C0",
 30151 => x"C0C0C0B0C0F992F9",
 30152 => x"C0C0C0B0C0F992A4",
 30153 => x"C0C0C0B0C0F992B0",
 30154 => x"C0C0C0B0C0F99299",
 30155 => x"C0C0C0B0C0F99292",
 30156 => x"C0C0C0B0C0F99282",
 30157 => x"C0C0C0B0C0F992F8",
 30158 => x"C0C0C0B0C0F99280",
 30159 => x"C0C0C0B0C0F99290",
 30160 => x"C0C0C0B0C0F982C0",
 30161 => x"C0C0C0B0C0F982F9",
 30162 => x"C0C0C0B0C0F982A4",
 30163 => x"C0C0C0B0C0F982B0",
 30164 => x"C0C0C0B0C0F98299",
 30165 => x"C0C0C0B0C0F98292",
 30166 => x"C0C0C0B0C0F98282",
 30167 => x"C0C0C0B0C0F982F8",
 30168 => x"C0C0C0B0C0F98280",
 30169 => x"C0C0C0B0C0F98290",
 30170 => x"C0C0C0B0C0F9F8C0",
 30171 => x"C0C0C0B0C0F9F8F9",
 30172 => x"C0C0C0B0C0F9F8A4",
 30173 => x"C0C0C0B0C0F9F8B0",
 30174 => x"C0C0C0B0C0F9F899",
 30175 => x"C0C0C0B0C0F9F892",
 30176 => x"C0C0C0B0C0F9F882",
 30177 => x"C0C0C0B0C0F9F8F8",
 30178 => x"C0C0C0B0C0F9F880",
 30179 => x"C0C0C0B0C0F9F890",
 30180 => x"C0C0C0B0C0F980C0",
 30181 => x"C0C0C0B0C0F980F9",
 30182 => x"C0C0C0B0C0F980A4",
 30183 => x"C0C0C0B0C0F980B0",
 30184 => x"C0C0C0B0C0F98099",
 30185 => x"C0C0C0B0C0F98092",
 30186 => x"C0C0C0B0C0F98082",
 30187 => x"C0C0C0B0C0F980F8",
 30188 => x"C0C0C0B0C0F98080",
 30189 => x"C0C0C0B0C0F98090",
 30190 => x"C0C0C0B0C0F990C0",
 30191 => x"C0C0C0B0C0F990F9",
 30192 => x"C0C0C0B0C0F990A4",
 30193 => x"C0C0C0B0C0F990B0",
 30194 => x"C0C0C0B0C0F99099",
 30195 => x"C0C0C0B0C0F99092",
 30196 => x"C0C0C0B0C0F99082",
 30197 => x"C0C0C0B0C0F990F8",
 30198 => x"C0C0C0B0C0F99080",
 30199 => x"C0C0C0B0C0F99090",
 30200 => x"C0C0C0B0C0A4C0C0",
 30201 => x"C0C0C0B0C0A4C0F9",
 30202 => x"C0C0C0B0C0A4C0A4",
 30203 => x"C0C0C0B0C0A4C0B0",
 30204 => x"C0C0C0B0C0A4C099",
 30205 => x"C0C0C0B0C0A4C092",
 30206 => x"C0C0C0B0C0A4C082",
 30207 => x"C0C0C0B0C0A4C0F8",
 30208 => x"C0C0C0B0C0A4C080",
 30209 => x"C0C0C0B0C0A4C090",
 30210 => x"C0C0C0B0C0A4F9C0",
 30211 => x"C0C0C0B0C0A4F9F9",
 30212 => x"C0C0C0B0C0A4F9A4",
 30213 => x"C0C0C0B0C0A4F9B0",
 30214 => x"C0C0C0B0C0A4F999",
 30215 => x"C0C0C0B0C0A4F992",
 30216 => x"C0C0C0B0C0A4F982",
 30217 => x"C0C0C0B0C0A4F9F8",
 30218 => x"C0C0C0B0C0A4F980",
 30219 => x"C0C0C0B0C0A4F990",
 30220 => x"C0C0C0B0C0A4A4C0",
 30221 => x"C0C0C0B0C0A4A4F9",
 30222 => x"C0C0C0B0C0A4A4A4",
 30223 => x"C0C0C0B0C0A4A4B0",
 30224 => x"C0C0C0B0C0A4A499",
 30225 => x"C0C0C0B0C0A4A492",
 30226 => x"C0C0C0B0C0A4A482",
 30227 => x"C0C0C0B0C0A4A4F8",
 30228 => x"C0C0C0B0C0A4A480",
 30229 => x"C0C0C0B0C0A4A490",
 30230 => x"C0C0C0B0C0A4B0C0",
 30231 => x"C0C0C0B0C0A4B0F9",
 30232 => x"C0C0C0B0C0A4B0A4",
 30233 => x"C0C0C0B0C0A4B0B0",
 30234 => x"C0C0C0B0C0A4B099",
 30235 => x"C0C0C0B0C0A4B092",
 30236 => x"C0C0C0B0C0A4B082",
 30237 => x"C0C0C0B0C0A4B0F8",
 30238 => x"C0C0C0B0C0A4B080",
 30239 => x"C0C0C0B0C0A4B090",
 30240 => x"C0C0C0B0C0A499C0",
 30241 => x"C0C0C0B0C0A499F9",
 30242 => x"C0C0C0B0C0A499A4",
 30243 => x"C0C0C0B0C0A499B0",
 30244 => x"C0C0C0B0C0A49999",
 30245 => x"C0C0C0B0C0A49992",
 30246 => x"C0C0C0B0C0A49982",
 30247 => x"C0C0C0B0C0A499F8",
 30248 => x"C0C0C0B0C0A49980",
 30249 => x"C0C0C0B0C0A49990",
 30250 => x"C0C0C0B0C0A492C0",
 30251 => x"C0C0C0B0C0A492F9",
 30252 => x"C0C0C0B0C0A492A4",
 30253 => x"C0C0C0B0C0A492B0",
 30254 => x"C0C0C0B0C0A49299",
 30255 => x"C0C0C0B0C0A49292",
 30256 => x"C0C0C0B0C0A49282",
 30257 => x"C0C0C0B0C0A492F8",
 30258 => x"C0C0C0B0C0A49280",
 30259 => x"C0C0C0B0C0A49290",
 30260 => x"C0C0C0B0C0A482C0",
 30261 => x"C0C0C0B0C0A482F9",
 30262 => x"C0C0C0B0C0A482A4",
 30263 => x"C0C0C0B0C0A482B0",
 30264 => x"C0C0C0B0C0A48299",
 30265 => x"C0C0C0B0C0A48292",
 30266 => x"C0C0C0B0C0A48282",
 30267 => x"C0C0C0B0C0A482F8",
 30268 => x"C0C0C0B0C0A48280",
 30269 => x"C0C0C0B0C0A48290",
 30270 => x"C0C0C0B0C0A4F8C0",
 30271 => x"C0C0C0B0C0A4F8F9",
 30272 => x"C0C0C0B0C0A4F8A4",
 30273 => x"C0C0C0B0C0A4F8B0",
 30274 => x"C0C0C0B0C0A4F899",
 30275 => x"C0C0C0B0C0A4F892",
 30276 => x"C0C0C0B0C0A4F882",
 30277 => x"C0C0C0B0C0A4F8F8",
 30278 => x"C0C0C0B0C0A4F880",
 30279 => x"C0C0C0B0C0A4F890",
 30280 => x"C0C0C0B0C0A480C0",
 30281 => x"C0C0C0B0C0A480F9",
 30282 => x"C0C0C0B0C0A480A4",
 30283 => x"C0C0C0B0C0A480B0",
 30284 => x"C0C0C0B0C0A48099",
 30285 => x"C0C0C0B0C0A48092",
 30286 => x"C0C0C0B0C0A48082",
 30287 => x"C0C0C0B0C0A480F8",
 30288 => x"C0C0C0B0C0A48080",
 30289 => x"C0C0C0B0C0A48090",
 30290 => x"C0C0C0B0C0A490C0",
 30291 => x"C0C0C0B0C0A490F9",
 30292 => x"C0C0C0B0C0A490A4",
 30293 => x"C0C0C0B0C0A490B0",
 30294 => x"C0C0C0B0C0A49099",
 30295 => x"C0C0C0B0C0A49092",
 30296 => x"C0C0C0B0C0A49082",
 30297 => x"C0C0C0B0C0A490F8",
 30298 => x"C0C0C0B0C0A49080",
 30299 => x"C0C0C0B0C0A49090",
 30300 => x"C0C0C0B0C0B0C0C0",
 30301 => x"C0C0C0B0C0B0C0F9",
 30302 => x"C0C0C0B0C0B0C0A4",
 30303 => x"C0C0C0B0C0B0C0B0",
 30304 => x"C0C0C0B0C0B0C099",
 30305 => x"C0C0C0B0C0B0C092",
 30306 => x"C0C0C0B0C0B0C082",
 30307 => x"C0C0C0B0C0B0C0F8",
 30308 => x"C0C0C0B0C0B0C080",
 30309 => x"C0C0C0B0C0B0C090",
 30310 => x"C0C0C0B0C0B0F9C0",
 30311 => x"C0C0C0B0C0B0F9F9",
 30312 => x"C0C0C0B0C0B0F9A4",
 30313 => x"C0C0C0B0C0B0F9B0",
 30314 => x"C0C0C0B0C0B0F999",
 30315 => x"C0C0C0B0C0B0F992",
 30316 => x"C0C0C0B0C0B0F982",
 30317 => x"C0C0C0B0C0B0F9F8",
 30318 => x"C0C0C0B0C0B0F980",
 30319 => x"C0C0C0B0C0B0F990",
 30320 => x"C0C0C0B0C0B0A4C0",
 30321 => x"C0C0C0B0C0B0A4F9",
 30322 => x"C0C0C0B0C0B0A4A4",
 30323 => x"C0C0C0B0C0B0A4B0",
 30324 => x"C0C0C0B0C0B0A499",
 30325 => x"C0C0C0B0C0B0A492",
 30326 => x"C0C0C0B0C0B0A482",
 30327 => x"C0C0C0B0C0B0A4F8",
 30328 => x"C0C0C0B0C0B0A480",
 30329 => x"C0C0C0B0C0B0A490",
 30330 => x"C0C0C0B0C0B0B0C0",
 30331 => x"C0C0C0B0C0B0B0F9",
 30332 => x"C0C0C0B0C0B0B0A4",
 30333 => x"C0C0C0B0C0B0B0B0",
 30334 => x"C0C0C0B0C0B0B099",
 30335 => x"C0C0C0B0C0B0B092",
 30336 => x"C0C0C0B0C0B0B082",
 30337 => x"C0C0C0B0C0B0B0F8",
 30338 => x"C0C0C0B0C0B0B080",
 30339 => x"C0C0C0B0C0B0B090",
 30340 => x"C0C0C0B0C0B099C0",
 30341 => x"C0C0C0B0C0B099F9",
 30342 => x"C0C0C0B0C0B099A4",
 30343 => x"C0C0C0B0C0B099B0",
 30344 => x"C0C0C0B0C0B09999",
 30345 => x"C0C0C0B0C0B09992",
 30346 => x"C0C0C0B0C0B09982",
 30347 => x"C0C0C0B0C0B099F8",
 30348 => x"C0C0C0B0C0B09980",
 30349 => x"C0C0C0B0C0B09990",
 30350 => x"C0C0C0B0C0B092C0",
 30351 => x"C0C0C0B0C0B092F9",
 30352 => x"C0C0C0B0C0B092A4",
 30353 => x"C0C0C0B0C0B092B0",
 30354 => x"C0C0C0B0C0B09299",
 30355 => x"C0C0C0B0C0B09292",
 30356 => x"C0C0C0B0C0B09282",
 30357 => x"C0C0C0B0C0B092F8",
 30358 => x"C0C0C0B0C0B09280",
 30359 => x"C0C0C0B0C0B09290",
 30360 => x"C0C0C0B0C0B082C0",
 30361 => x"C0C0C0B0C0B082F9",
 30362 => x"C0C0C0B0C0B082A4",
 30363 => x"C0C0C0B0C0B082B0",
 30364 => x"C0C0C0B0C0B08299",
 30365 => x"C0C0C0B0C0B08292",
 30366 => x"C0C0C0B0C0B08282",
 30367 => x"C0C0C0B0C0B082F8",
 30368 => x"C0C0C0B0C0B08280",
 30369 => x"C0C0C0B0C0B08290",
 30370 => x"C0C0C0B0C0B0F8C0",
 30371 => x"C0C0C0B0C0B0F8F9",
 30372 => x"C0C0C0B0C0B0F8A4",
 30373 => x"C0C0C0B0C0B0F8B0",
 30374 => x"C0C0C0B0C0B0F899",
 30375 => x"C0C0C0B0C0B0F892",
 30376 => x"C0C0C0B0C0B0F882",
 30377 => x"C0C0C0B0C0B0F8F8",
 30378 => x"C0C0C0B0C0B0F880",
 30379 => x"C0C0C0B0C0B0F890",
 30380 => x"C0C0C0B0C0B080C0",
 30381 => x"C0C0C0B0C0B080F9",
 30382 => x"C0C0C0B0C0B080A4",
 30383 => x"C0C0C0B0C0B080B0",
 30384 => x"C0C0C0B0C0B08099",
 30385 => x"C0C0C0B0C0B08092",
 30386 => x"C0C0C0B0C0B08082",
 30387 => x"C0C0C0B0C0B080F8",
 30388 => x"C0C0C0B0C0B08080",
 30389 => x"C0C0C0B0C0B08090",
 30390 => x"C0C0C0B0C0B090C0",
 30391 => x"C0C0C0B0C0B090F9",
 30392 => x"C0C0C0B0C0B090A4",
 30393 => x"C0C0C0B0C0B090B0",
 30394 => x"C0C0C0B0C0B09099",
 30395 => x"C0C0C0B0C0B09092",
 30396 => x"C0C0C0B0C0B09082",
 30397 => x"C0C0C0B0C0B090F8",
 30398 => x"C0C0C0B0C0B09080",
 30399 => x"C0C0C0B0C0B09090",
 30400 => x"C0C0C0B0C099C0C0",
 30401 => x"C0C0C0B0C099C0F9",
 30402 => x"C0C0C0B0C099C0A4",
 30403 => x"C0C0C0B0C099C0B0",
 30404 => x"C0C0C0B0C099C099",
 30405 => x"C0C0C0B0C099C092",
 30406 => x"C0C0C0B0C099C082",
 30407 => x"C0C0C0B0C099C0F8",
 30408 => x"C0C0C0B0C099C080",
 30409 => x"C0C0C0B0C099C090",
 30410 => x"C0C0C0B0C099F9C0",
 30411 => x"C0C0C0B0C099F9F9",
 30412 => x"C0C0C0B0C099F9A4",
 30413 => x"C0C0C0B0C099F9B0",
 30414 => x"C0C0C0B0C099F999",
 30415 => x"C0C0C0B0C099F992",
 30416 => x"C0C0C0B0C099F982",
 30417 => x"C0C0C0B0C099F9F8",
 30418 => x"C0C0C0B0C099F980",
 30419 => x"C0C0C0B0C099F990",
 30420 => x"C0C0C0B0C099A4C0",
 30421 => x"C0C0C0B0C099A4F9",
 30422 => x"C0C0C0B0C099A4A4",
 30423 => x"C0C0C0B0C099A4B0",
 30424 => x"C0C0C0B0C099A499",
 30425 => x"C0C0C0B0C099A492",
 30426 => x"C0C0C0B0C099A482",
 30427 => x"C0C0C0B0C099A4F8",
 30428 => x"C0C0C0B0C099A480",
 30429 => x"C0C0C0B0C099A490",
 30430 => x"C0C0C0B0C099B0C0",
 30431 => x"C0C0C0B0C099B0F9",
 30432 => x"C0C0C0B0C099B0A4",
 30433 => x"C0C0C0B0C099B0B0",
 30434 => x"C0C0C0B0C099B099",
 30435 => x"C0C0C0B0C099B092",
 30436 => x"C0C0C0B0C099B082",
 30437 => x"C0C0C0B0C099B0F8",
 30438 => x"C0C0C0B0C099B080",
 30439 => x"C0C0C0B0C099B090",
 30440 => x"C0C0C0B0C09999C0",
 30441 => x"C0C0C0B0C09999F9",
 30442 => x"C0C0C0B0C09999A4",
 30443 => x"C0C0C0B0C09999B0",
 30444 => x"C0C0C0B0C0999999",
 30445 => x"C0C0C0B0C0999992",
 30446 => x"C0C0C0B0C0999982",
 30447 => x"C0C0C0B0C09999F8",
 30448 => x"C0C0C0B0C0999980",
 30449 => x"C0C0C0B0C0999990",
 30450 => x"C0C0C0B0C09992C0",
 30451 => x"C0C0C0B0C09992F9",
 30452 => x"C0C0C0B0C09992A4",
 30453 => x"C0C0C0B0C09992B0",
 30454 => x"C0C0C0B0C0999299",
 30455 => x"C0C0C0B0C0999292",
 30456 => x"C0C0C0B0C0999282",
 30457 => x"C0C0C0B0C09992F8",
 30458 => x"C0C0C0B0C0999280",
 30459 => x"C0C0C0B0C0999290",
 30460 => x"C0C0C0B0C09982C0",
 30461 => x"C0C0C0B0C09982F9",
 30462 => x"C0C0C0B0C09982A4",
 30463 => x"C0C0C0B0C09982B0",
 30464 => x"C0C0C0B0C0998299",
 30465 => x"C0C0C0B0C0998292",
 30466 => x"C0C0C0B0C0998282",
 30467 => x"C0C0C0B0C09982F8",
 30468 => x"C0C0C0B0C0998280",
 30469 => x"C0C0C0B0C0998290",
 30470 => x"C0C0C0B0C099F8C0",
 30471 => x"C0C0C0B0C099F8F9",
 30472 => x"C0C0C0B0C099F8A4",
 30473 => x"C0C0C0B0C099F8B0",
 30474 => x"C0C0C0B0C099F899",
 30475 => x"C0C0C0B0C099F892",
 30476 => x"C0C0C0B0C099F882",
 30477 => x"C0C0C0B0C099F8F8",
 30478 => x"C0C0C0B0C099F880",
 30479 => x"C0C0C0B0C099F890",
 30480 => x"C0C0C0B0C09980C0",
 30481 => x"C0C0C0B0C09980F9",
 30482 => x"C0C0C0B0C09980A4",
 30483 => x"C0C0C0B0C09980B0",
 30484 => x"C0C0C0B0C0998099",
 30485 => x"C0C0C0B0C0998092",
 30486 => x"C0C0C0B0C0998082",
 30487 => x"C0C0C0B0C09980F8",
 30488 => x"C0C0C0B0C0998080",
 30489 => x"C0C0C0B0C0998090",
 30490 => x"C0C0C0B0C09990C0",
 30491 => x"C0C0C0B0C09990F9",
 30492 => x"C0C0C0B0C09990A4",
 30493 => x"C0C0C0B0C09990B0",
 30494 => x"C0C0C0B0C0999099",
 30495 => x"C0C0C0B0C0999092",
 30496 => x"C0C0C0B0C0999082",
 30497 => x"C0C0C0B0C09990F8",
 30498 => x"C0C0C0B0C0999080",
 30499 => x"C0C0C0B0C0999090",
 30500 => x"C0C0C0B0C092C0C0",
 30501 => x"C0C0C0B0C092C0F9",
 30502 => x"C0C0C0B0C092C0A4",
 30503 => x"C0C0C0B0C092C0B0",
 30504 => x"C0C0C0B0C092C099",
 30505 => x"C0C0C0B0C092C092",
 30506 => x"C0C0C0B0C092C082",
 30507 => x"C0C0C0B0C092C0F8",
 30508 => x"C0C0C0B0C092C080",
 30509 => x"C0C0C0B0C092C090",
 30510 => x"C0C0C0B0C092F9C0",
 30511 => x"C0C0C0B0C092F9F9",
 30512 => x"C0C0C0B0C092F9A4",
 30513 => x"C0C0C0B0C092F9B0",
 30514 => x"C0C0C0B0C092F999",
 30515 => x"C0C0C0B0C092F992",
 30516 => x"C0C0C0B0C092F982",
 30517 => x"C0C0C0B0C092F9F8",
 30518 => x"C0C0C0B0C092F980",
 30519 => x"C0C0C0B0C092F990",
 30520 => x"C0C0C0B0C092A4C0",
 30521 => x"C0C0C0B0C092A4F9",
 30522 => x"C0C0C0B0C092A4A4",
 30523 => x"C0C0C0B0C092A4B0",
 30524 => x"C0C0C0B0C092A499",
 30525 => x"C0C0C0B0C092A492",
 30526 => x"C0C0C0B0C092A482",
 30527 => x"C0C0C0B0C092A4F8",
 30528 => x"C0C0C0B0C092A480",
 30529 => x"C0C0C0B0C092A490",
 30530 => x"C0C0C0B0C092B0C0",
 30531 => x"C0C0C0B0C092B0F9",
 30532 => x"C0C0C0B0C092B0A4",
 30533 => x"C0C0C0B0C092B0B0",
 30534 => x"C0C0C0B0C092B099",
 30535 => x"C0C0C0B0C092B092",
 30536 => x"C0C0C0B0C092B082",
 30537 => x"C0C0C0B0C092B0F8",
 30538 => x"C0C0C0B0C092B080",
 30539 => x"C0C0C0B0C092B090",
 30540 => x"C0C0C0B0C09299C0",
 30541 => x"C0C0C0B0C09299F9",
 30542 => x"C0C0C0B0C09299A4",
 30543 => x"C0C0C0B0C09299B0",
 30544 => x"C0C0C0B0C0929999",
 30545 => x"C0C0C0B0C0929992",
 30546 => x"C0C0C0B0C0929982",
 30547 => x"C0C0C0B0C09299F8",
 30548 => x"C0C0C0B0C0929980",
 30549 => x"C0C0C0B0C0929990",
 30550 => x"C0C0C0B0C09292C0",
 30551 => x"C0C0C0B0C09292F9",
 30552 => x"C0C0C0B0C09292A4",
 30553 => x"C0C0C0B0C09292B0",
 30554 => x"C0C0C0B0C0929299",
 30555 => x"C0C0C0B0C0929292",
 30556 => x"C0C0C0B0C0929282",
 30557 => x"C0C0C0B0C09292F8",
 30558 => x"C0C0C0B0C0929280",
 30559 => x"C0C0C0B0C0929290",
 30560 => x"C0C0C0B0C09282C0",
 30561 => x"C0C0C0B0C09282F9",
 30562 => x"C0C0C0B0C09282A4",
 30563 => x"C0C0C0B0C09282B0",
 30564 => x"C0C0C0B0C0928299",
 30565 => x"C0C0C0B0C0928292",
 30566 => x"C0C0C0B0C0928282",
 30567 => x"C0C0C0B0C09282F8",
 30568 => x"C0C0C0B0C0928280",
 30569 => x"C0C0C0B0C0928290",
 30570 => x"C0C0C0B0C092F8C0",
 30571 => x"C0C0C0B0C092F8F9",
 30572 => x"C0C0C0B0C092F8A4",
 30573 => x"C0C0C0B0C092F8B0",
 30574 => x"C0C0C0B0C092F899",
 30575 => x"C0C0C0B0C092F892",
 30576 => x"C0C0C0B0C092F882",
 30577 => x"C0C0C0B0C092F8F8",
 30578 => x"C0C0C0B0C092F880",
 30579 => x"C0C0C0B0C092F890",
 30580 => x"C0C0C0B0C09280C0",
 30581 => x"C0C0C0B0C09280F9",
 30582 => x"C0C0C0B0C09280A4",
 30583 => x"C0C0C0B0C09280B0",
 30584 => x"C0C0C0B0C0928099",
 30585 => x"C0C0C0B0C0928092",
 30586 => x"C0C0C0B0C0928082",
 30587 => x"C0C0C0B0C09280F8",
 30588 => x"C0C0C0B0C0928080",
 30589 => x"C0C0C0B0C0928090",
 30590 => x"C0C0C0B0C09290C0",
 30591 => x"C0C0C0B0C09290F9",
 30592 => x"C0C0C0B0C09290A4",
 30593 => x"C0C0C0B0C09290B0",
 30594 => x"C0C0C0B0C0929099",
 30595 => x"C0C0C0B0C0929092",
 30596 => x"C0C0C0B0C0929082",
 30597 => x"C0C0C0B0C09290F8",
 30598 => x"C0C0C0B0C0929080",
 30599 => x"C0C0C0B0C0929090",
 30600 => x"C0C0C0B0C082C0C0",
 30601 => x"C0C0C0B0C082C0F9",
 30602 => x"C0C0C0B0C082C0A4",
 30603 => x"C0C0C0B0C082C0B0",
 30604 => x"C0C0C0B0C082C099",
 30605 => x"C0C0C0B0C082C092",
 30606 => x"C0C0C0B0C082C082",
 30607 => x"C0C0C0B0C082C0F8",
 30608 => x"C0C0C0B0C082C080",
 30609 => x"C0C0C0B0C082C090",
 30610 => x"C0C0C0B0C082F9C0",
 30611 => x"C0C0C0B0C082F9F9",
 30612 => x"C0C0C0B0C082F9A4",
 30613 => x"C0C0C0B0C082F9B0",
 30614 => x"C0C0C0B0C082F999",
 30615 => x"C0C0C0B0C082F992",
 30616 => x"C0C0C0B0C082F982",
 30617 => x"C0C0C0B0C082F9F8",
 30618 => x"C0C0C0B0C082F980",
 30619 => x"C0C0C0B0C082F990",
 30620 => x"C0C0C0B0C082A4C0",
 30621 => x"C0C0C0B0C082A4F9",
 30622 => x"C0C0C0B0C082A4A4",
 30623 => x"C0C0C0B0C082A4B0",
 30624 => x"C0C0C0B0C082A499",
 30625 => x"C0C0C0B0C082A492",
 30626 => x"C0C0C0B0C082A482",
 30627 => x"C0C0C0B0C082A4F8",
 30628 => x"C0C0C0B0C082A480",
 30629 => x"C0C0C0B0C082A490",
 30630 => x"C0C0C0B0C082B0C0",
 30631 => x"C0C0C0B0C082B0F9",
 30632 => x"C0C0C0B0C082B0A4",
 30633 => x"C0C0C0B0C082B0B0",
 30634 => x"C0C0C0B0C082B099",
 30635 => x"C0C0C0B0C082B092",
 30636 => x"C0C0C0B0C082B082",
 30637 => x"C0C0C0B0C082B0F8",
 30638 => x"C0C0C0B0C082B080",
 30639 => x"C0C0C0B0C082B090",
 30640 => x"C0C0C0B0C08299C0",
 30641 => x"C0C0C0B0C08299F9",
 30642 => x"C0C0C0B0C08299A4",
 30643 => x"C0C0C0B0C08299B0",
 30644 => x"C0C0C0B0C0829999",
 30645 => x"C0C0C0B0C0829992",
 30646 => x"C0C0C0B0C0829982",
 30647 => x"C0C0C0B0C08299F8",
 30648 => x"C0C0C0B0C0829980",
 30649 => x"C0C0C0B0C0829990",
 30650 => x"C0C0C0B0C08292C0",
 30651 => x"C0C0C0B0C08292F9",
 30652 => x"C0C0C0B0C08292A4",
 30653 => x"C0C0C0B0C08292B0",
 30654 => x"C0C0C0B0C0829299",
 30655 => x"C0C0C0B0C0829292",
 30656 => x"C0C0C0B0C0829282",
 30657 => x"C0C0C0B0C08292F8",
 30658 => x"C0C0C0B0C0829280",
 30659 => x"C0C0C0B0C0829290",
 30660 => x"C0C0C0B0C08282C0",
 30661 => x"C0C0C0B0C08282F9",
 30662 => x"C0C0C0B0C08282A4",
 30663 => x"C0C0C0B0C08282B0",
 30664 => x"C0C0C0B0C0828299",
 30665 => x"C0C0C0B0C0828292",
 30666 => x"C0C0C0B0C0828282",
 30667 => x"C0C0C0B0C08282F8",
 30668 => x"C0C0C0B0C0828280",
 30669 => x"C0C0C0B0C0828290",
 30670 => x"C0C0C0B0C082F8C0",
 30671 => x"C0C0C0B0C082F8F9",
 30672 => x"C0C0C0B0C082F8A4",
 30673 => x"C0C0C0B0C082F8B0",
 30674 => x"C0C0C0B0C082F899",
 30675 => x"C0C0C0B0C082F892",
 30676 => x"C0C0C0B0C082F882",
 30677 => x"C0C0C0B0C082F8F8",
 30678 => x"C0C0C0B0C082F880",
 30679 => x"C0C0C0B0C082F890",
 30680 => x"C0C0C0B0C08280C0",
 30681 => x"C0C0C0B0C08280F9",
 30682 => x"C0C0C0B0C08280A4",
 30683 => x"C0C0C0B0C08280B0",
 30684 => x"C0C0C0B0C0828099",
 30685 => x"C0C0C0B0C0828092",
 30686 => x"C0C0C0B0C0828082",
 30687 => x"C0C0C0B0C08280F8",
 30688 => x"C0C0C0B0C0828080",
 30689 => x"C0C0C0B0C0828090",
 30690 => x"C0C0C0B0C08290C0",
 30691 => x"C0C0C0B0C08290F9",
 30692 => x"C0C0C0B0C08290A4",
 30693 => x"C0C0C0B0C08290B0",
 30694 => x"C0C0C0B0C0829099",
 30695 => x"C0C0C0B0C0829092",
 30696 => x"C0C0C0B0C0829082",
 30697 => x"C0C0C0B0C08290F8",
 30698 => x"C0C0C0B0C0829080",
 30699 => x"C0C0C0B0C0829090",
 30700 => x"C0C0C0B0C0F8C0C0",
 30701 => x"C0C0C0B0C0F8C0F9",
 30702 => x"C0C0C0B0C0F8C0A4",
 30703 => x"C0C0C0B0C0F8C0B0",
 30704 => x"C0C0C0B0C0F8C099",
 30705 => x"C0C0C0B0C0F8C092",
 30706 => x"C0C0C0B0C0F8C082",
 30707 => x"C0C0C0B0C0F8C0F8",
 30708 => x"C0C0C0B0C0F8C080",
 30709 => x"C0C0C0B0C0F8C090",
 30710 => x"C0C0C0B0C0F8F9C0",
 30711 => x"C0C0C0B0C0F8F9F9",
 30712 => x"C0C0C0B0C0F8F9A4",
 30713 => x"C0C0C0B0C0F8F9B0",
 30714 => x"C0C0C0B0C0F8F999",
 30715 => x"C0C0C0B0C0F8F992",
 30716 => x"C0C0C0B0C0F8F982",
 30717 => x"C0C0C0B0C0F8F9F8",
 30718 => x"C0C0C0B0C0F8F980",
 30719 => x"C0C0C0B0C0F8F990",
 30720 => x"C0C0C0B0C0F8A4C0",
 30721 => x"C0C0C0B0C0F8A4F9",
 30722 => x"C0C0C0B0C0F8A4A4",
 30723 => x"C0C0C0B0C0F8A4B0",
 30724 => x"C0C0C0B0C0F8A499",
 30725 => x"C0C0C0B0C0F8A492",
 30726 => x"C0C0C0B0C0F8A482",
 30727 => x"C0C0C0B0C0F8A4F8",
 30728 => x"C0C0C0B0C0F8A480",
 30729 => x"C0C0C0B0C0F8A490",
 30730 => x"C0C0C0B0C0F8B0C0",
 30731 => x"C0C0C0B0C0F8B0F9",
 30732 => x"C0C0C0B0C0F8B0A4",
 30733 => x"C0C0C0B0C0F8B0B0",
 30734 => x"C0C0C0B0C0F8B099",
 30735 => x"C0C0C0B0C0F8B092",
 30736 => x"C0C0C0B0C0F8B082",
 30737 => x"C0C0C0B0C0F8B0F8",
 30738 => x"C0C0C0B0C0F8B080",
 30739 => x"C0C0C0B0C0F8B090",
 30740 => x"C0C0C0B0C0F899C0",
 30741 => x"C0C0C0B0C0F899F9",
 30742 => x"C0C0C0B0C0F899A4",
 30743 => x"C0C0C0B0C0F899B0",
 30744 => x"C0C0C0B0C0F89999",
 30745 => x"C0C0C0B0C0F89992",
 30746 => x"C0C0C0B0C0F89982",
 30747 => x"C0C0C0B0C0F899F8",
 30748 => x"C0C0C0B0C0F89980",
 30749 => x"C0C0C0B0C0F89990",
 30750 => x"C0C0C0B0C0F892C0",
 30751 => x"C0C0C0B0C0F892F9",
 30752 => x"C0C0C0B0C0F892A4",
 30753 => x"C0C0C0B0C0F892B0",
 30754 => x"C0C0C0B0C0F89299",
 30755 => x"C0C0C0B0C0F89292",
 30756 => x"C0C0C0B0C0F89282",
 30757 => x"C0C0C0B0C0F892F8",
 30758 => x"C0C0C0B0C0F89280",
 30759 => x"C0C0C0B0C0F89290",
 30760 => x"C0C0C0B0C0F882C0",
 30761 => x"C0C0C0B0C0F882F9",
 30762 => x"C0C0C0B0C0F882A4",
 30763 => x"C0C0C0B0C0F882B0",
 30764 => x"C0C0C0B0C0F88299",
 30765 => x"C0C0C0B0C0F88292",
 30766 => x"C0C0C0B0C0F88282",
 30767 => x"C0C0C0B0C0F882F8",
 30768 => x"C0C0C0B0C0F88280",
 30769 => x"C0C0C0B0C0F88290",
 30770 => x"C0C0C0B0C0F8F8C0",
 30771 => x"C0C0C0B0C0F8F8F9",
 30772 => x"C0C0C0B0C0F8F8A4",
 30773 => x"C0C0C0B0C0F8F8B0",
 30774 => x"C0C0C0B0C0F8F899",
 30775 => x"C0C0C0B0C0F8F892",
 30776 => x"C0C0C0B0C0F8F882",
 30777 => x"C0C0C0B0C0F8F8F8",
 30778 => x"C0C0C0B0C0F8F880",
 30779 => x"C0C0C0B0C0F8F890",
 30780 => x"C0C0C0B0C0F880C0",
 30781 => x"C0C0C0B0C0F880F9",
 30782 => x"C0C0C0B0C0F880A4",
 30783 => x"C0C0C0B0C0F880B0",
 30784 => x"C0C0C0B0C0F88099",
 30785 => x"C0C0C0B0C0F88092",
 30786 => x"C0C0C0B0C0F88082",
 30787 => x"C0C0C0B0C0F880F8",
 30788 => x"C0C0C0B0C0F88080",
 30789 => x"C0C0C0B0C0F88090",
 30790 => x"C0C0C0B0C0F890C0",
 30791 => x"C0C0C0B0C0F890F9",
 30792 => x"C0C0C0B0C0F890A4",
 30793 => x"C0C0C0B0C0F890B0",
 30794 => x"C0C0C0B0C0F89099",
 30795 => x"C0C0C0B0C0F89092",
 30796 => x"C0C0C0B0C0F89082",
 30797 => x"C0C0C0B0C0F890F8",
 30798 => x"C0C0C0B0C0F89080",
 30799 => x"C0C0C0B0C0F89090",
 30800 => x"C0C0C0B0C080C0C0",
 30801 => x"C0C0C0B0C080C0F9",
 30802 => x"C0C0C0B0C080C0A4",
 30803 => x"C0C0C0B0C080C0B0",
 30804 => x"C0C0C0B0C080C099",
 30805 => x"C0C0C0B0C080C092",
 30806 => x"C0C0C0B0C080C082",
 30807 => x"C0C0C0B0C080C0F8",
 30808 => x"C0C0C0B0C080C080",
 30809 => x"C0C0C0B0C080C090",
 30810 => x"C0C0C0B0C080F9C0",
 30811 => x"C0C0C0B0C080F9F9",
 30812 => x"C0C0C0B0C080F9A4",
 30813 => x"C0C0C0B0C080F9B0",
 30814 => x"C0C0C0B0C080F999",
 30815 => x"C0C0C0B0C080F992",
 30816 => x"C0C0C0B0C080F982",
 30817 => x"C0C0C0B0C080F9F8",
 30818 => x"C0C0C0B0C080F980",
 30819 => x"C0C0C0B0C080F990",
 30820 => x"C0C0C0B0C080A4C0",
 30821 => x"C0C0C0B0C080A4F9",
 30822 => x"C0C0C0B0C080A4A4",
 30823 => x"C0C0C0B0C080A4B0",
 30824 => x"C0C0C0B0C080A499",
 30825 => x"C0C0C0B0C080A492",
 30826 => x"C0C0C0B0C080A482",
 30827 => x"C0C0C0B0C080A4F8",
 30828 => x"C0C0C0B0C080A480",
 30829 => x"C0C0C0B0C080A490",
 30830 => x"C0C0C0B0C080B0C0",
 30831 => x"C0C0C0B0C080B0F9",
 30832 => x"C0C0C0B0C080B0A4",
 30833 => x"C0C0C0B0C080B0B0",
 30834 => x"C0C0C0B0C080B099",
 30835 => x"C0C0C0B0C080B092",
 30836 => x"C0C0C0B0C080B082",
 30837 => x"C0C0C0B0C080B0F8",
 30838 => x"C0C0C0B0C080B080",
 30839 => x"C0C0C0B0C080B090",
 30840 => x"C0C0C0B0C08099C0",
 30841 => x"C0C0C0B0C08099F9",
 30842 => x"C0C0C0B0C08099A4",
 30843 => x"C0C0C0B0C08099B0",
 30844 => x"C0C0C0B0C0809999",
 30845 => x"C0C0C0B0C0809992",
 30846 => x"C0C0C0B0C0809982",
 30847 => x"C0C0C0B0C08099F8",
 30848 => x"C0C0C0B0C0809980",
 30849 => x"C0C0C0B0C0809990",
 30850 => x"C0C0C0B0C08092C0",
 30851 => x"C0C0C0B0C08092F9",
 30852 => x"C0C0C0B0C08092A4",
 30853 => x"C0C0C0B0C08092B0",
 30854 => x"C0C0C0B0C0809299",
 30855 => x"C0C0C0B0C0809292",
 30856 => x"C0C0C0B0C0809282",
 30857 => x"C0C0C0B0C08092F8",
 30858 => x"C0C0C0B0C0809280",
 30859 => x"C0C0C0B0C0809290",
 30860 => x"C0C0C0B0C08082C0",
 30861 => x"C0C0C0B0C08082F9",
 30862 => x"C0C0C0B0C08082A4",
 30863 => x"C0C0C0B0C08082B0",
 30864 => x"C0C0C0B0C0808299",
 30865 => x"C0C0C0B0C0808292",
 30866 => x"C0C0C0B0C0808282",
 30867 => x"C0C0C0B0C08082F8",
 30868 => x"C0C0C0B0C0808280",
 30869 => x"C0C0C0B0C0808290",
 30870 => x"C0C0C0B0C080F8C0",
 30871 => x"C0C0C0B0C080F8F9",
 30872 => x"C0C0C0B0C080F8A4",
 30873 => x"C0C0C0B0C080F8B0",
 30874 => x"C0C0C0B0C080F899",
 30875 => x"C0C0C0B0C080F892",
 30876 => x"C0C0C0B0C080F882",
 30877 => x"C0C0C0B0C080F8F8",
 30878 => x"C0C0C0B0C080F880",
 30879 => x"C0C0C0B0C080F890",
 30880 => x"C0C0C0B0C08080C0",
 30881 => x"C0C0C0B0C08080F9",
 30882 => x"C0C0C0B0C08080A4",
 30883 => x"C0C0C0B0C08080B0",
 30884 => x"C0C0C0B0C0808099",
 30885 => x"C0C0C0B0C0808092",
 30886 => x"C0C0C0B0C0808082",
 30887 => x"C0C0C0B0C08080F8",
 30888 => x"C0C0C0B0C0808080",
 30889 => x"C0C0C0B0C0808090",
 30890 => x"C0C0C0B0C08090C0",
 30891 => x"C0C0C0B0C08090F9",
 30892 => x"C0C0C0B0C08090A4",
 30893 => x"C0C0C0B0C08090B0",
 30894 => x"C0C0C0B0C0809099",
 30895 => x"C0C0C0B0C0809092",
 30896 => x"C0C0C0B0C0809082",
 30897 => x"C0C0C0B0C08090F8",
 30898 => x"C0C0C0B0C0809080",
 30899 => x"C0C0C0B0C0809090",
 30900 => x"C0C0C0B0C090C0C0",
 30901 => x"C0C0C0B0C090C0F9",
 30902 => x"C0C0C0B0C090C0A4",
 30903 => x"C0C0C0B0C090C0B0",
 30904 => x"C0C0C0B0C090C099",
 30905 => x"C0C0C0B0C090C092",
 30906 => x"C0C0C0B0C090C082",
 30907 => x"C0C0C0B0C090C0F8",
 30908 => x"C0C0C0B0C090C080",
 30909 => x"C0C0C0B0C090C090",
 30910 => x"C0C0C0B0C090F9C0",
 30911 => x"C0C0C0B0C090F9F9",
 30912 => x"C0C0C0B0C090F9A4",
 30913 => x"C0C0C0B0C090F9B0",
 30914 => x"C0C0C0B0C090F999",
 30915 => x"C0C0C0B0C090F992",
 30916 => x"C0C0C0B0C090F982",
 30917 => x"C0C0C0B0C090F9F8",
 30918 => x"C0C0C0B0C090F980",
 30919 => x"C0C0C0B0C090F990",
 30920 => x"C0C0C0B0C090A4C0",
 30921 => x"C0C0C0B0C090A4F9",
 30922 => x"C0C0C0B0C090A4A4",
 30923 => x"C0C0C0B0C090A4B0",
 30924 => x"C0C0C0B0C090A499",
 30925 => x"C0C0C0B0C090A492",
 30926 => x"C0C0C0B0C090A482",
 30927 => x"C0C0C0B0C090A4F8",
 30928 => x"C0C0C0B0C090A480",
 30929 => x"C0C0C0B0C090A490",
 30930 => x"C0C0C0B0C090B0C0",
 30931 => x"C0C0C0B0C090B0F9",
 30932 => x"C0C0C0B0C090B0A4",
 30933 => x"C0C0C0B0C090B0B0",
 30934 => x"C0C0C0B0C090B099",
 30935 => x"C0C0C0B0C090B092",
 30936 => x"C0C0C0B0C090B082",
 30937 => x"C0C0C0B0C090B0F8",
 30938 => x"C0C0C0B0C090B080",
 30939 => x"C0C0C0B0C090B090",
 30940 => x"C0C0C0B0C09099C0",
 30941 => x"C0C0C0B0C09099F9",
 30942 => x"C0C0C0B0C09099A4",
 30943 => x"C0C0C0B0C09099B0",
 30944 => x"C0C0C0B0C0909999",
 30945 => x"C0C0C0B0C0909992",
 30946 => x"C0C0C0B0C0909982",
 30947 => x"C0C0C0B0C09099F8",
 30948 => x"C0C0C0B0C0909980",
 30949 => x"C0C0C0B0C0909990",
 30950 => x"C0C0C0B0C09092C0",
 30951 => x"C0C0C0B0C09092F9",
 30952 => x"C0C0C0B0C09092A4",
 30953 => x"C0C0C0B0C09092B0",
 30954 => x"C0C0C0B0C0909299",
 30955 => x"C0C0C0B0C0909292",
 30956 => x"C0C0C0B0C0909282",
 30957 => x"C0C0C0B0C09092F8",
 30958 => x"C0C0C0B0C0909280",
 30959 => x"C0C0C0B0C0909290",
 30960 => x"C0C0C0B0C09082C0",
 30961 => x"C0C0C0B0C09082F9",
 30962 => x"C0C0C0B0C09082A4",
 30963 => x"C0C0C0B0C09082B0",
 30964 => x"C0C0C0B0C0908299",
 30965 => x"C0C0C0B0C0908292",
 30966 => x"C0C0C0B0C0908282",
 30967 => x"C0C0C0B0C09082F8",
 30968 => x"C0C0C0B0C0908280",
 30969 => x"C0C0C0B0C0908290",
 30970 => x"C0C0C0B0C090F8C0",
 30971 => x"C0C0C0B0C090F8F9",
 30972 => x"C0C0C0B0C090F8A4",
 30973 => x"C0C0C0B0C090F8B0",
 30974 => x"C0C0C0B0C090F899",
 30975 => x"C0C0C0B0C090F892",
 30976 => x"C0C0C0B0C090F882",
 30977 => x"C0C0C0B0C090F8F8",
 30978 => x"C0C0C0B0C090F880",
 30979 => x"C0C0C0B0C090F890",
 30980 => x"C0C0C0B0C09080C0",
 30981 => x"C0C0C0B0C09080F9",
 30982 => x"C0C0C0B0C09080A4",
 30983 => x"C0C0C0B0C09080B0",
 30984 => x"C0C0C0B0C0908099",
 30985 => x"C0C0C0B0C0908092",
 30986 => x"C0C0C0B0C0908082",
 30987 => x"C0C0C0B0C09080F8",
 30988 => x"C0C0C0B0C0908080",
 30989 => x"C0C0C0B0C0908090",
 30990 => x"C0C0C0B0C09090C0",
 30991 => x"C0C0C0B0C09090F9",
 30992 => x"C0C0C0B0C09090A4",
 30993 => x"C0C0C0B0C09090B0",
 30994 => x"C0C0C0B0C0909099",
 30995 => x"C0C0C0B0C0909092",
 30996 => x"C0C0C0B0C0909082",
 30997 => x"C0C0C0B0C09090F8",
 30998 => x"C0C0C0B0C0909080",
 30999 => x"C0C0C0B0C0909090",
 31000 => x"C0C0C0B0F9C0C0C0",
 31001 => x"C0C0C0B0F9C0C0F9",
 31002 => x"C0C0C0B0F9C0C0A4",
 31003 => x"C0C0C0B0F9C0C0B0",
 31004 => x"C0C0C0B0F9C0C099",
 31005 => x"C0C0C0B0F9C0C092",
 31006 => x"C0C0C0B0F9C0C082",
 31007 => x"C0C0C0B0F9C0C0F8",
 31008 => x"C0C0C0B0F9C0C080",
 31009 => x"C0C0C0B0F9C0C090",
 31010 => x"C0C0C0B0F9C0F9C0",
 31011 => x"C0C0C0B0F9C0F9F9",
 31012 => x"C0C0C0B0F9C0F9A4",
 31013 => x"C0C0C0B0F9C0F9B0",
 31014 => x"C0C0C0B0F9C0F999",
 31015 => x"C0C0C0B0F9C0F992",
 31016 => x"C0C0C0B0F9C0F982",
 31017 => x"C0C0C0B0F9C0F9F8",
 31018 => x"C0C0C0B0F9C0F980",
 31019 => x"C0C0C0B0F9C0F990",
 31020 => x"C0C0C0B0F9C0A4C0",
 31021 => x"C0C0C0B0F9C0A4F9",
 31022 => x"C0C0C0B0F9C0A4A4",
 31023 => x"C0C0C0B0F9C0A4B0",
 31024 => x"C0C0C0B0F9C0A499",
 31025 => x"C0C0C0B0F9C0A492",
 31026 => x"C0C0C0B0F9C0A482",
 31027 => x"C0C0C0B0F9C0A4F8",
 31028 => x"C0C0C0B0F9C0A480",
 31029 => x"C0C0C0B0F9C0A490",
 31030 => x"C0C0C0B0F9C0B0C0",
 31031 => x"C0C0C0B0F9C0B0F9",
 31032 => x"C0C0C0B0F9C0B0A4",
 31033 => x"C0C0C0B0F9C0B0B0",
 31034 => x"C0C0C0B0F9C0B099",
 31035 => x"C0C0C0B0F9C0B092",
 31036 => x"C0C0C0B0F9C0B082",
 31037 => x"C0C0C0B0F9C0B0F8",
 31038 => x"C0C0C0B0F9C0B080",
 31039 => x"C0C0C0B0F9C0B090",
 31040 => x"C0C0C0B0F9C099C0",
 31041 => x"C0C0C0B0F9C099F9",
 31042 => x"C0C0C0B0F9C099A4",
 31043 => x"C0C0C0B0F9C099B0",
 31044 => x"C0C0C0B0F9C09999",
 31045 => x"C0C0C0B0F9C09992",
 31046 => x"C0C0C0B0F9C09982",
 31047 => x"C0C0C0B0F9C099F8",
 31048 => x"C0C0C0B0F9C09980",
 31049 => x"C0C0C0B0F9C09990",
 31050 => x"C0C0C0B0F9C092C0",
 31051 => x"C0C0C0B0F9C092F9",
 31052 => x"C0C0C0B0F9C092A4",
 31053 => x"C0C0C0B0F9C092B0",
 31054 => x"C0C0C0B0F9C09299",
 31055 => x"C0C0C0B0F9C09292",
 31056 => x"C0C0C0B0F9C09282",
 31057 => x"C0C0C0B0F9C092F8",
 31058 => x"C0C0C0B0F9C09280",
 31059 => x"C0C0C0B0F9C09290",
 31060 => x"C0C0C0B0F9C082C0",
 31061 => x"C0C0C0B0F9C082F9",
 31062 => x"C0C0C0B0F9C082A4",
 31063 => x"C0C0C0B0F9C082B0",
 31064 => x"C0C0C0B0F9C08299",
 31065 => x"C0C0C0B0F9C08292",
 31066 => x"C0C0C0B0F9C08282",
 31067 => x"C0C0C0B0F9C082F8",
 31068 => x"C0C0C0B0F9C08280",
 31069 => x"C0C0C0B0F9C08290",
 31070 => x"C0C0C0B0F9C0F8C0",
 31071 => x"C0C0C0B0F9C0F8F9",
 31072 => x"C0C0C0B0F9C0F8A4",
 31073 => x"C0C0C0B0F9C0F8B0",
 31074 => x"C0C0C0B0F9C0F899",
 31075 => x"C0C0C0B0F9C0F892",
 31076 => x"C0C0C0B0F9C0F882",
 31077 => x"C0C0C0B0F9C0F8F8",
 31078 => x"C0C0C0B0F9C0F880",
 31079 => x"C0C0C0B0F9C0F890",
 31080 => x"C0C0C0B0F9C080C0",
 31081 => x"C0C0C0B0F9C080F9",
 31082 => x"C0C0C0B0F9C080A4",
 31083 => x"C0C0C0B0F9C080B0",
 31084 => x"C0C0C0B0F9C08099",
 31085 => x"C0C0C0B0F9C08092",
 31086 => x"C0C0C0B0F9C08082",
 31087 => x"C0C0C0B0F9C080F8",
 31088 => x"C0C0C0B0F9C08080",
 31089 => x"C0C0C0B0F9C08090",
 31090 => x"C0C0C0B0F9C090C0",
 31091 => x"C0C0C0B0F9C090F9",
 31092 => x"C0C0C0B0F9C090A4",
 31093 => x"C0C0C0B0F9C090B0",
 31094 => x"C0C0C0B0F9C09099",
 31095 => x"C0C0C0B0F9C09092",
 31096 => x"C0C0C0B0F9C09082",
 31097 => x"C0C0C0B0F9C090F8",
 31098 => x"C0C0C0B0F9C09080",
 31099 => x"C0C0C0B0F9C09090",
 31100 => x"C0C0C0B0F9F9C0C0",
 31101 => x"C0C0C0B0F9F9C0F9",
 31102 => x"C0C0C0B0F9F9C0A4",
 31103 => x"C0C0C0B0F9F9C0B0",
 31104 => x"C0C0C0B0F9F9C099",
 31105 => x"C0C0C0B0F9F9C092",
 31106 => x"C0C0C0B0F9F9C082",
 31107 => x"C0C0C0B0F9F9C0F8",
 31108 => x"C0C0C0B0F9F9C080",
 31109 => x"C0C0C0B0F9F9C090",
 31110 => x"C0C0C0B0F9F9F9C0",
 31111 => x"C0C0C0B0F9F9F9F9",
 31112 => x"C0C0C0B0F9F9F9A4",
 31113 => x"C0C0C0B0F9F9F9B0",
 31114 => x"C0C0C0B0F9F9F999",
 31115 => x"C0C0C0B0F9F9F992",
 31116 => x"C0C0C0B0F9F9F982",
 31117 => x"C0C0C0B0F9F9F9F8",
 31118 => x"C0C0C0B0F9F9F980",
 31119 => x"C0C0C0B0F9F9F990",
 31120 => x"C0C0C0B0F9F9A4C0",
 31121 => x"C0C0C0B0F9F9A4F9",
 31122 => x"C0C0C0B0F9F9A4A4",
 31123 => x"C0C0C0B0F9F9A4B0",
 31124 => x"C0C0C0B0F9F9A499",
 31125 => x"C0C0C0B0F9F9A492",
 31126 => x"C0C0C0B0F9F9A482",
 31127 => x"C0C0C0B0F9F9A4F8",
 31128 => x"C0C0C0B0F9F9A480",
 31129 => x"C0C0C0B0F9F9A490",
 31130 => x"C0C0C0B0F9F9B0C0",
 31131 => x"C0C0C0B0F9F9B0F9",
 31132 => x"C0C0C0B0F9F9B0A4",
 31133 => x"C0C0C0B0F9F9B0B0",
 31134 => x"C0C0C0B0F9F9B099",
 31135 => x"C0C0C0B0F9F9B092",
 31136 => x"C0C0C0B0F9F9B082",
 31137 => x"C0C0C0B0F9F9B0F8",
 31138 => x"C0C0C0B0F9F9B080",
 31139 => x"C0C0C0B0F9F9B090",
 31140 => x"C0C0C0B0F9F999C0",
 31141 => x"C0C0C0B0F9F999F9",
 31142 => x"C0C0C0B0F9F999A4",
 31143 => x"C0C0C0B0F9F999B0",
 31144 => x"C0C0C0B0F9F99999",
 31145 => x"C0C0C0B0F9F99992",
 31146 => x"C0C0C0B0F9F99982",
 31147 => x"C0C0C0B0F9F999F8",
 31148 => x"C0C0C0B0F9F99980",
 31149 => x"C0C0C0B0F9F99990",
 31150 => x"C0C0C0B0F9F992C0",
 31151 => x"C0C0C0B0F9F992F9",
 31152 => x"C0C0C0B0F9F992A4",
 31153 => x"C0C0C0B0F9F992B0",
 31154 => x"C0C0C0B0F9F99299",
 31155 => x"C0C0C0B0F9F99292",
 31156 => x"C0C0C0B0F9F99282",
 31157 => x"C0C0C0B0F9F992F8",
 31158 => x"C0C0C0B0F9F99280",
 31159 => x"C0C0C0B0F9F99290",
 31160 => x"C0C0C0B0F9F982C0",
 31161 => x"C0C0C0B0F9F982F9",
 31162 => x"C0C0C0B0F9F982A4",
 31163 => x"C0C0C0B0F9F982B0",
 31164 => x"C0C0C0B0F9F98299",
 31165 => x"C0C0C0B0F9F98292",
 31166 => x"C0C0C0B0F9F98282",
 31167 => x"C0C0C0B0F9F982F8",
 31168 => x"C0C0C0B0F9F98280",
 31169 => x"C0C0C0B0F9F98290",
 31170 => x"C0C0C0B0F9F9F8C0",
 31171 => x"C0C0C0B0F9F9F8F9",
 31172 => x"C0C0C0B0F9F9F8A4",
 31173 => x"C0C0C0B0F9F9F8B0",
 31174 => x"C0C0C0B0F9F9F899",
 31175 => x"C0C0C0B0F9F9F892",
 31176 => x"C0C0C0B0F9F9F882",
 31177 => x"C0C0C0B0F9F9F8F8",
 31178 => x"C0C0C0B0F9F9F880",
 31179 => x"C0C0C0B0F9F9F890",
 31180 => x"C0C0C0B0F9F980C0",
 31181 => x"C0C0C0B0F9F980F9",
 31182 => x"C0C0C0B0F9F980A4",
 31183 => x"C0C0C0B0F9F980B0",
 31184 => x"C0C0C0B0F9F98099",
 31185 => x"C0C0C0B0F9F98092",
 31186 => x"C0C0C0B0F9F98082",
 31187 => x"C0C0C0B0F9F980F8",
 31188 => x"C0C0C0B0F9F98080",
 31189 => x"C0C0C0B0F9F98090",
 31190 => x"C0C0C0B0F9F990C0",
 31191 => x"C0C0C0B0F9F990F9",
 31192 => x"C0C0C0B0F9F990A4",
 31193 => x"C0C0C0B0F9F990B0",
 31194 => x"C0C0C0B0F9F99099",
 31195 => x"C0C0C0B0F9F99092",
 31196 => x"C0C0C0B0F9F99082",
 31197 => x"C0C0C0B0F9F990F8",
 31198 => x"C0C0C0B0F9F99080",
 31199 => x"C0C0C0B0F9F99090",
 31200 => x"C0C0C0B0F9A4C0C0",
 31201 => x"C0C0C0B0F9A4C0F9",
 31202 => x"C0C0C0B0F9A4C0A4",
 31203 => x"C0C0C0B0F9A4C0B0",
 31204 => x"C0C0C0B0F9A4C099",
 31205 => x"C0C0C0B0F9A4C092",
 31206 => x"C0C0C0B0F9A4C082",
 31207 => x"C0C0C0B0F9A4C0F8",
 31208 => x"C0C0C0B0F9A4C080",
 31209 => x"C0C0C0B0F9A4C090",
 31210 => x"C0C0C0B0F9A4F9C0",
 31211 => x"C0C0C0B0F9A4F9F9",
 31212 => x"C0C0C0B0F9A4F9A4",
 31213 => x"C0C0C0B0F9A4F9B0",
 31214 => x"C0C0C0B0F9A4F999",
 31215 => x"C0C0C0B0F9A4F992",
 31216 => x"C0C0C0B0F9A4F982",
 31217 => x"C0C0C0B0F9A4F9F8",
 31218 => x"C0C0C0B0F9A4F980",
 31219 => x"C0C0C0B0F9A4F990",
 31220 => x"C0C0C0B0F9A4A4C0",
 31221 => x"C0C0C0B0F9A4A4F9",
 31222 => x"C0C0C0B0F9A4A4A4",
 31223 => x"C0C0C0B0F9A4A4B0",
 31224 => x"C0C0C0B0F9A4A499",
 31225 => x"C0C0C0B0F9A4A492",
 31226 => x"C0C0C0B0F9A4A482",
 31227 => x"C0C0C0B0F9A4A4F8",
 31228 => x"C0C0C0B0F9A4A480",
 31229 => x"C0C0C0B0F9A4A490",
 31230 => x"C0C0C0B0F9A4B0C0",
 31231 => x"C0C0C0B0F9A4B0F9",
 31232 => x"C0C0C0B0F9A4B0A4",
 31233 => x"C0C0C0B0F9A4B0B0",
 31234 => x"C0C0C0B0F9A4B099",
 31235 => x"C0C0C0B0F9A4B092",
 31236 => x"C0C0C0B0F9A4B082",
 31237 => x"C0C0C0B0F9A4B0F8",
 31238 => x"C0C0C0B0F9A4B080",
 31239 => x"C0C0C0B0F9A4B090",
 31240 => x"C0C0C0B0F9A499C0",
 31241 => x"C0C0C0B0F9A499F9",
 31242 => x"C0C0C0B0F9A499A4",
 31243 => x"C0C0C0B0F9A499B0",
 31244 => x"C0C0C0B0F9A49999",
 31245 => x"C0C0C0B0F9A49992",
 31246 => x"C0C0C0B0F9A49982",
 31247 => x"C0C0C0B0F9A499F8",
 31248 => x"C0C0C0B0F9A49980",
 31249 => x"C0C0C0B0F9A49990",
 31250 => x"C0C0C0B0F9A492C0",
 31251 => x"C0C0C0B0F9A492F9",
 31252 => x"C0C0C0B0F9A492A4",
 31253 => x"C0C0C0B0F9A492B0",
 31254 => x"C0C0C0B0F9A49299",
 31255 => x"C0C0C0B0F9A49292",
 31256 => x"C0C0C0B0F9A49282",
 31257 => x"C0C0C0B0F9A492F8",
 31258 => x"C0C0C0B0F9A49280",
 31259 => x"C0C0C0B0F9A49290",
 31260 => x"C0C0C0B0F9A482C0",
 31261 => x"C0C0C0B0F9A482F9",
 31262 => x"C0C0C0B0F9A482A4",
 31263 => x"C0C0C0B0F9A482B0",
 31264 => x"C0C0C0B0F9A48299",
 31265 => x"C0C0C0B0F9A48292",
 31266 => x"C0C0C0B0F9A48282",
 31267 => x"C0C0C0B0F9A482F8",
 31268 => x"C0C0C0B0F9A48280",
 31269 => x"C0C0C0B0F9A48290",
 31270 => x"C0C0C0B0F9A4F8C0",
 31271 => x"C0C0C0B0F9A4F8F9",
 31272 => x"C0C0C0B0F9A4F8A4",
 31273 => x"C0C0C0B0F9A4F8B0",
 31274 => x"C0C0C0B0F9A4F899",
 31275 => x"C0C0C0B0F9A4F892",
 31276 => x"C0C0C0B0F9A4F882",
 31277 => x"C0C0C0B0F9A4F8F8",
 31278 => x"C0C0C0B0F9A4F880",
 31279 => x"C0C0C0B0F9A4F890",
 31280 => x"C0C0C0B0F9A480C0",
 31281 => x"C0C0C0B0F9A480F9",
 31282 => x"C0C0C0B0F9A480A4",
 31283 => x"C0C0C0B0F9A480B0",
 31284 => x"C0C0C0B0F9A48099",
 31285 => x"C0C0C0B0F9A48092",
 31286 => x"C0C0C0B0F9A48082",
 31287 => x"C0C0C0B0F9A480F8",
 31288 => x"C0C0C0B0F9A48080",
 31289 => x"C0C0C0B0F9A48090",
 31290 => x"C0C0C0B0F9A490C0",
 31291 => x"C0C0C0B0F9A490F9",
 31292 => x"C0C0C0B0F9A490A4",
 31293 => x"C0C0C0B0F9A490B0",
 31294 => x"C0C0C0B0F9A49099",
 31295 => x"C0C0C0B0F9A49092",
 31296 => x"C0C0C0B0F9A49082",
 31297 => x"C0C0C0B0F9A490F8",
 31298 => x"C0C0C0B0F9A49080",
 31299 => x"C0C0C0B0F9A49090",
 31300 => x"C0C0C0B0F9B0C0C0",
 31301 => x"C0C0C0B0F9B0C0F9",
 31302 => x"C0C0C0B0F9B0C0A4",
 31303 => x"C0C0C0B0F9B0C0B0",
 31304 => x"C0C0C0B0F9B0C099",
 31305 => x"C0C0C0B0F9B0C092",
 31306 => x"C0C0C0B0F9B0C082",
 31307 => x"C0C0C0B0F9B0C0F8",
 31308 => x"C0C0C0B0F9B0C080",
 31309 => x"C0C0C0B0F9B0C090",
 31310 => x"C0C0C0B0F9B0F9C0",
 31311 => x"C0C0C0B0F9B0F9F9",
 31312 => x"C0C0C0B0F9B0F9A4",
 31313 => x"C0C0C0B0F9B0F9B0",
 31314 => x"C0C0C0B0F9B0F999",
 31315 => x"C0C0C0B0F9B0F992",
 31316 => x"C0C0C0B0F9B0F982",
 31317 => x"C0C0C0B0F9B0F9F8",
 31318 => x"C0C0C0B0F9B0F980",
 31319 => x"C0C0C0B0F9B0F990",
 31320 => x"C0C0C0B0F9B0A4C0",
 31321 => x"C0C0C0B0F9B0A4F9",
 31322 => x"C0C0C0B0F9B0A4A4",
 31323 => x"C0C0C0B0F9B0A4B0",
 31324 => x"C0C0C0B0F9B0A499",
 31325 => x"C0C0C0B0F9B0A492",
 31326 => x"C0C0C0B0F9B0A482",
 31327 => x"C0C0C0B0F9B0A4F8",
 31328 => x"C0C0C0B0F9B0A480",
 31329 => x"C0C0C0B0F9B0A490",
 31330 => x"C0C0C0B0F9B0B0C0",
 31331 => x"C0C0C0B0F9B0B0F9",
 31332 => x"C0C0C0B0F9B0B0A4",
 31333 => x"C0C0C0B0F9B0B0B0",
 31334 => x"C0C0C0B0F9B0B099",
 31335 => x"C0C0C0B0F9B0B092",
 31336 => x"C0C0C0B0F9B0B082",
 31337 => x"C0C0C0B0F9B0B0F8",
 31338 => x"C0C0C0B0F9B0B080",
 31339 => x"C0C0C0B0F9B0B090",
 31340 => x"C0C0C0B0F9B099C0",
 31341 => x"C0C0C0B0F9B099F9",
 31342 => x"C0C0C0B0F9B099A4",
 31343 => x"C0C0C0B0F9B099B0",
 31344 => x"C0C0C0B0F9B09999",
 31345 => x"C0C0C0B0F9B09992",
 31346 => x"C0C0C0B0F9B09982",
 31347 => x"C0C0C0B0F9B099F8",
 31348 => x"C0C0C0B0F9B09980",
 31349 => x"C0C0C0B0F9B09990",
 31350 => x"C0C0C0B0F9B092C0",
 31351 => x"C0C0C0B0F9B092F9",
 31352 => x"C0C0C0B0F9B092A4",
 31353 => x"C0C0C0B0F9B092B0",
 31354 => x"C0C0C0B0F9B09299",
 31355 => x"C0C0C0B0F9B09292",
 31356 => x"C0C0C0B0F9B09282",
 31357 => x"C0C0C0B0F9B092F8",
 31358 => x"C0C0C0B0F9B09280",
 31359 => x"C0C0C0B0F9B09290",
 31360 => x"C0C0C0B0F9B082C0",
 31361 => x"C0C0C0B0F9B082F9",
 31362 => x"C0C0C0B0F9B082A4",
 31363 => x"C0C0C0B0F9B082B0",
 31364 => x"C0C0C0B0F9B08299",
 31365 => x"C0C0C0B0F9B08292",
 31366 => x"C0C0C0B0F9B08282",
 31367 => x"C0C0C0B0F9B082F8",
 31368 => x"C0C0C0B0F9B08280",
 31369 => x"C0C0C0B0F9B08290",
 31370 => x"C0C0C0B0F9B0F8C0",
 31371 => x"C0C0C0B0F9B0F8F9",
 31372 => x"C0C0C0B0F9B0F8A4",
 31373 => x"C0C0C0B0F9B0F8B0",
 31374 => x"C0C0C0B0F9B0F899",
 31375 => x"C0C0C0B0F9B0F892",
 31376 => x"C0C0C0B0F9B0F882",
 31377 => x"C0C0C0B0F9B0F8F8",
 31378 => x"C0C0C0B0F9B0F880",
 31379 => x"C0C0C0B0F9B0F890",
 31380 => x"C0C0C0B0F9B080C0",
 31381 => x"C0C0C0B0F9B080F9",
 31382 => x"C0C0C0B0F9B080A4",
 31383 => x"C0C0C0B0F9B080B0",
 31384 => x"C0C0C0B0F9B08099",
 31385 => x"C0C0C0B0F9B08092",
 31386 => x"C0C0C0B0F9B08082",
 31387 => x"C0C0C0B0F9B080F8",
 31388 => x"C0C0C0B0F9B08080",
 31389 => x"C0C0C0B0F9B08090",
 31390 => x"C0C0C0B0F9B090C0",
 31391 => x"C0C0C0B0F9B090F9",
 31392 => x"C0C0C0B0F9B090A4",
 31393 => x"C0C0C0B0F9B090B0",
 31394 => x"C0C0C0B0F9B09099",
 31395 => x"C0C0C0B0F9B09092",
 31396 => x"C0C0C0B0F9B09082",
 31397 => x"C0C0C0B0F9B090F8",
 31398 => x"C0C0C0B0F9B09080",
 31399 => x"C0C0C0B0F9B09090",
 31400 => x"C0C0C0B0F999C0C0",
 31401 => x"C0C0C0B0F999C0F9",
 31402 => x"C0C0C0B0F999C0A4",
 31403 => x"C0C0C0B0F999C0B0",
 31404 => x"C0C0C0B0F999C099",
 31405 => x"C0C0C0B0F999C092",
 31406 => x"C0C0C0B0F999C082",
 31407 => x"C0C0C0B0F999C0F8",
 31408 => x"C0C0C0B0F999C080",
 31409 => x"C0C0C0B0F999C090",
 31410 => x"C0C0C0B0F999F9C0",
 31411 => x"C0C0C0B0F999F9F9",
 31412 => x"C0C0C0B0F999F9A4",
 31413 => x"C0C0C0B0F999F9B0",
 31414 => x"C0C0C0B0F999F999",
 31415 => x"C0C0C0B0F999F992",
 31416 => x"C0C0C0B0F999F982",
 31417 => x"C0C0C0B0F999F9F8",
 31418 => x"C0C0C0B0F999F980",
 31419 => x"C0C0C0B0F999F990",
 31420 => x"C0C0C0B0F999A4C0",
 31421 => x"C0C0C0B0F999A4F9",
 31422 => x"C0C0C0B0F999A4A4",
 31423 => x"C0C0C0B0F999A4B0",
 31424 => x"C0C0C0B0F999A499",
 31425 => x"C0C0C0B0F999A492",
 31426 => x"C0C0C0B0F999A482",
 31427 => x"C0C0C0B0F999A4F8",
 31428 => x"C0C0C0B0F999A480",
 31429 => x"C0C0C0B0F999A490",
 31430 => x"C0C0C0B0F999B0C0",
 31431 => x"C0C0C0B0F999B0F9",
 31432 => x"C0C0C0B0F999B0A4",
 31433 => x"C0C0C0B0F999B0B0",
 31434 => x"C0C0C0B0F999B099",
 31435 => x"C0C0C0B0F999B092",
 31436 => x"C0C0C0B0F999B082",
 31437 => x"C0C0C0B0F999B0F8",
 31438 => x"C0C0C0B0F999B080",
 31439 => x"C0C0C0B0F999B090",
 31440 => x"C0C0C0B0F99999C0",
 31441 => x"C0C0C0B0F99999F9",
 31442 => x"C0C0C0B0F99999A4",
 31443 => x"C0C0C0B0F99999B0",
 31444 => x"C0C0C0B0F9999999",
 31445 => x"C0C0C0B0F9999992",
 31446 => x"C0C0C0B0F9999982",
 31447 => x"C0C0C0B0F99999F8",
 31448 => x"C0C0C0B0F9999980",
 31449 => x"C0C0C0B0F9999990",
 31450 => x"C0C0C0B0F99992C0",
 31451 => x"C0C0C0B0F99992F9",
 31452 => x"C0C0C0B0F99992A4",
 31453 => x"C0C0C0B0F99992B0",
 31454 => x"C0C0C0B0F9999299",
 31455 => x"C0C0C0B0F9999292",
 31456 => x"C0C0C0B0F9999282",
 31457 => x"C0C0C0B0F99992F8",
 31458 => x"C0C0C0B0F9999280",
 31459 => x"C0C0C0B0F9999290",
 31460 => x"C0C0C0B0F99982C0",
 31461 => x"C0C0C0B0F99982F9",
 31462 => x"C0C0C0B0F99982A4",
 31463 => x"C0C0C0B0F99982B0",
 31464 => x"C0C0C0B0F9998299",
 31465 => x"C0C0C0B0F9998292",
 31466 => x"C0C0C0B0F9998282",
 31467 => x"C0C0C0B0F99982F8",
 31468 => x"C0C0C0B0F9998280",
 31469 => x"C0C0C0B0F9998290",
 31470 => x"C0C0C0B0F999F8C0",
 31471 => x"C0C0C0B0F999F8F9",
 31472 => x"C0C0C0B0F999F8A4",
 31473 => x"C0C0C0B0F999F8B0",
 31474 => x"C0C0C0B0F999F899",
 31475 => x"C0C0C0B0F999F892",
 31476 => x"C0C0C0B0F999F882",
 31477 => x"C0C0C0B0F999F8F8",
 31478 => x"C0C0C0B0F999F880",
 31479 => x"C0C0C0B0F999F890",
 31480 => x"C0C0C0B0F99980C0",
 31481 => x"C0C0C0B0F99980F9",
 31482 => x"C0C0C0B0F99980A4",
 31483 => x"C0C0C0B0F99980B0",
 31484 => x"C0C0C0B0F9998099",
 31485 => x"C0C0C0B0F9998092",
 31486 => x"C0C0C0B0F9998082",
 31487 => x"C0C0C0B0F99980F8",
 31488 => x"C0C0C0B0F9998080",
 31489 => x"C0C0C0B0F9998090",
 31490 => x"C0C0C0B0F99990C0",
 31491 => x"C0C0C0B0F99990F9",
 31492 => x"C0C0C0B0F99990A4",
 31493 => x"C0C0C0B0F99990B0",
 31494 => x"C0C0C0B0F9999099",
 31495 => x"C0C0C0B0F9999092",
 31496 => x"C0C0C0B0F9999082",
 31497 => x"C0C0C0B0F99990F8",
 31498 => x"C0C0C0B0F9999080",
 31499 => x"C0C0C0B0F9999090",
 31500 => x"C0C0C0B0F992C0C0",
 31501 => x"C0C0C0B0F992C0F9",
 31502 => x"C0C0C0B0F992C0A4",
 31503 => x"C0C0C0B0F992C0B0",
 31504 => x"C0C0C0B0F992C099",
 31505 => x"C0C0C0B0F992C092",
 31506 => x"C0C0C0B0F992C082",
 31507 => x"C0C0C0B0F992C0F8",
 31508 => x"C0C0C0B0F992C080",
 31509 => x"C0C0C0B0F992C090",
 31510 => x"C0C0C0B0F992F9C0",
 31511 => x"C0C0C0B0F992F9F9",
 31512 => x"C0C0C0B0F992F9A4",
 31513 => x"C0C0C0B0F992F9B0",
 31514 => x"C0C0C0B0F992F999",
 31515 => x"C0C0C0B0F992F992",
 31516 => x"C0C0C0B0F992F982",
 31517 => x"C0C0C0B0F992F9F8",
 31518 => x"C0C0C0B0F992F980",
 31519 => x"C0C0C0B0F992F990",
 31520 => x"C0C0C0B0F992A4C0",
 31521 => x"C0C0C0B0F992A4F9",
 31522 => x"C0C0C0B0F992A4A4",
 31523 => x"C0C0C0B0F992A4B0",
 31524 => x"C0C0C0B0F992A499",
 31525 => x"C0C0C0B0F992A492",
 31526 => x"C0C0C0B0F992A482",
 31527 => x"C0C0C0B0F992A4F8",
 31528 => x"C0C0C0B0F992A480",
 31529 => x"C0C0C0B0F992A490",
 31530 => x"C0C0C0B0F992B0C0",
 31531 => x"C0C0C0B0F992B0F9",
 31532 => x"C0C0C0B0F992B0A4",
 31533 => x"C0C0C0B0F992B0B0",
 31534 => x"C0C0C0B0F992B099",
 31535 => x"C0C0C0B0F992B092",
 31536 => x"C0C0C0B0F992B082",
 31537 => x"C0C0C0B0F992B0F8",
 31538 => x"C0C0C0B0F992B080",
 31539 => x"C0C0C0B0F992B090",
 31540 => x"C0C0C0B0F99299C0",
 31541 => x"C0C0C0B0F99299F9",
 31542 => x"C0C0C0B0F99299A4",
 31543 => x"C0C0C0B0F99299B0",
 31544 => x"C0C0C0B0F9929999",
 31545 => x"C0C0C0B0F9929992",
 31546 => x"C0C0C0B0F9929982",
 31547 => x"C0C0C0B0F99299F8",
 31548 => x"C0C0C0B0F9929980",
 31549 => x"C0C0C0B0F9929990",
 31550 => x"C0C0C0B0F99292C0",
 31551 => x"C0C0C0B0F99292F9",
 31552 => x"C0C0C0B0F99292A4",
 31553 => x"C0C0C0B0F99292B0",
 31554 => x"C0C0C0B0F9929299",
 31555 => x"C0C0C0B0F9929292",
 31556 => x"C0C0C0B0F9929282",
 31557 => x"C0C0C0B0F99292F8",
 31558 => x"C0C0C0B0F9929280",
 31559 => x"C0C0C0B0F9929290",
 31560 => x"C0C0C0B0F99282C0",
 31561 => x"C0C0C0B0F99282F9",
 31562 => x"C0C0C0B0F99282A4",
 31563 => x"C0C0C0B0F99282B0",
 31564 => x"C0C0C0B0F9928299",
 31565 => x"C0C0C0B0F9928292",
 31566 => x"C0C0C0B0F9928282",
 31567 => x"C0C0C0B0F99282F8",
 31568 => x"C0C0C0B0F9928280",
 31569 => x"C0C0C0B0F9928290",
 31570 => x"C0C0C0B0F992F8C0",
 31571 => x"C0C0C0B0F992F8F9",
 31572 => x"C0C0C0B0F992F8A4",
 31573 => x"C0C0C0B0F992F8B0",
 31574 => x"C0C0C0B0F992F899",
 31575 => x"C0C0C0B0F992F892",
 31576 => x"C0C0C0B0F992F882",
 31577 => x"C0C0C0B0F992F8F8",
 31578 => x"C0C0C0B0F992F880",
 31579 => x"C0C0C0B0F992F890",
 31580 => x"C0C0C0B0F99280C0",
 31581 => x"C0C0C0B0F99280F9",
 31582 => x"C0C0C0B0F99280A4",
 31583 => x"C0C0C0B0F99280B0",
 31584 => x"C0C0C0B0F9928099",
 31585 => x"C0C0C0B0F9928092",
 31586 => x"C0C0C0B0F9928082",
 31587 => x"C0C0C0B0F99280F8",
 31588 => x"C0C0C0B0F9928080",
 31589 => x"C0C0C0B0F9928090",
 31590 => x"C0C0C0B0F99290C0",
 31591 => x"C0C0C0B0F99290F9",
 31592 => x"C0C0C0B0F99290A4",
 31593 => x"C0C0C0B0F99290B0",
 31594 => x"C0C0C0B0F9929099",
 31595 => x"C0C0C0B0F9929092",
 31596 => x"C0C0C0B0F9929082",
 31597 => x"C0C0C0B0F99290F8",
 31598 => x"C0C0C0B0F9929080",
 31599 => x"C0C0C0B0F9929090",
 31600 => x"C0C0C0B0F982C0C0",
 31601 => x"C0C0C0B0F982C0F9",
 31602 => x"C0C0C0B0F982C0A4",
 31603 => x"C0C0C0B0F982C0B0",
 31604 => x"C0C0C0B0F982C099",
 31605 => x"C0C0C0B0F982C092",
 31606 => x"C0C0C0B0F982C082",
 31607 => x"C0C0C0B0F982C0F8",
 31608 => x"C0C0C0B0F982C080",
 31609 => x"C0C0C0B0F982C090",
 31610 => x"C0C0C0B0F982F9C0",
 31611 => x"C0C0C0B0F982F9F9",
 31612 => x"C0C0C0B0F982F9A4",
 31613 => x"C0C0C0B0F982F9B0",
 31614 => x"C0C0C0B0F982F999",
 31615 => x"C0C0C0B0F982F992",
 31616 => x"C0C0C0B0F982F982",
 31617 => x"C0C0C0B0F982F9F8",
 31618 => x"C0C0C0B0F982F980",
 31619 => x"C0C0C0B0F982F990",
 31620 => x"C0C0C0B0F982A4C0",
 31621 => x"C0C0C0B0F982A4F9",
 31622 => x"C0C0C0B0F982A4A4",
 31623 => x"C0C0C0B0F982A4B0",
 31624 => x"C0C0C0B0F982A499",
 31625 => x"C0C0C0B0F982A492",
 31626 => x"C0C0C0B0F982A482",
 31627 => x"C0C0C0B0F982A4F8",
 31628 => x"C0C0C0B0F982A480",
 31629 => x"C0C0C0B0F982A490",
 31630 => x"C0C0C0B0F982B0C0",
 31631 => x"C0C0C0B0F982B0F9",
 31632 => x"C0C0C0B0F982B0A4",
 31633 => x"C0C0C0B0F982B0B0",
 31634 => x"C0C0C0B0F982B099",
 31635 => x"C0C0C0B0F982B092",
 31636 => x"C0C0C0B0F982B082",
 31637 => x"C0C0C0B0F982B0F8",
 31638 => x"C0C0C0B0F982B080",
 31639 => x"C0C0C0B0F982B090",
 31640 => x"C0C0C0B0F98299C0",
 31641 => x"C0C0C0B0F98299F9",
 31642 => x"C0C0C0B0F98299A4",
 31643 => x"C0C0C0B0F98299B0",
 31644 => x"C0C0C0B0F9829999",
 31645 => x"C0C0C0B0F9829992",
 31646 => x"C0C0C0B0F9829982",
 31647 => x"C0C0C0B0F98299F8",
 31648 => x"C0C0C0B0F9829980",
 31649 => x"C0C0C0B0F9829990",
 31650 => x"C0C0C0B0F98292C0",
 31651 => x"C0C0C0B0F98292F9",
 31652 => x"C0C0C0B0F98292A4",
 31653 => x"C0C0C0B0F98292B0",
 31654 => x"C0C0C0B0F9829299",
 31655 => x"C0C0C0B0F9829292",
 31656 => x"C0C0C0B0F9829282",
 31657 => x"C0C0C0B0F98292F8",
 31658 => x"C0C0C0B0F9829280",
 31659 => x"C0C0C0B0F9829290",
 31660 => x"C0C0C0B0F98282C0",
 31661 => x"C0C0C0B0F98282F9",
 31662 => x"C0C0C0B0F98282A4",
 31663 => x"C0C0C0B0F98282B0",
 31664 => x"C0C0C0B0F9828299",
 31665 => x"C0C0C0B0F9828292",
 31666 => x"C0C0C0B0F9828282",
 31667 => x"C0C0C0B0F98282F8",
 31668 => x"C0C0C0B0F9828280",
 31669 => x"C0C0C0B0F9828290",
 31670 => x"C0C0C0B0F982F8C0",
 31671 => x"C0C0C0B0F982F8F9",
 31672 => x"C0C0C0B0F982F8A4",
 31673 => x"C0C0C0B0F982F8B0",
 31674 => x"C0C0C0B0F982F899",
 31675 => x"C0C0C0B0F982F892",
 31676 => x"C0C0C0B0F982F882",
 31677 => x"C0C0C0B0F982F8F8",
 31678 => x"C0C0C0B0F982F880",
 31679 => x"C0C0C0B0F982F890",
 31680 => x"C0C0C0B0F98280C0",
 31681 => x"C0C0C0B0F98280F9",
 31682 => x"C0C0C0B0F98280A4",
 31683 => x"C0C0C0B0F98280B0",
 31684 => x"C0C0C0B0F9828099",
 31685 => x"C0C0C0B0F9828092",
 31686 => x"C0C0C0B0F9828082",
 31687 => x"C0C0C0B0F98280F8",
 31688 => x"C0C0C0B0F9828080",
 31689 => x"C0C0C0B0F9828090",
 31690 => x"C0C0C0B0F98290C0",
 31691 => x"C0C0C0B0F98290F9",
 31692 => x"C0C0C0B0F98290A4",
 31693 => x"C0C0C0B0F98290B0",
 31694 => x"C0C0C0B0F9829099",
 31695 => x"C0C0C0B0F9829092",
 31696 => x"C0C0C0B0F9829082",
 31697 => x"C0C0C0B0F98290F8",
 31698 => x"C0C0C0B0F9829080",
 31699 => x"C0C0C0B0F9829090",
 31700 => x"C0C0C0B0F9F8C0C0",
 31701 => x"C0C0C0B0F9F8C0F9",
 31702 => x"C0C0C0B0F9F8C0A4",
 31703 => x"C0C0C0B0F9F8C0B0",
 31704 => x"C0C0C0B0F9F8C099",
 31705 => x"C0C0C0B0F9F8C092",
 31706 => x"C0C0C0B0F9F8C082",
 31707 => x"C0C0C0B0F9F8C0F8",
 31708 => x"C0C0C0B0F9F8C080",
 31709 => x"C0C0C0B0F9F8C090",
 31710 => x"C0C0C0B0F9F8F9C0",
 31711 => x"C0C0C0B0F9F8F9F9",
 31712 => x"C0C0C0B0F9F8F9A4",
 31713 => x"C0C0C0B0F9F8F9B0",
 31714 => x"C0C0C0B0F9F8F999",
 31715 => x"C0C0C0B0F9F8F992",
 31716 => x"C0C0C0B0F9F8F982",
 31717 => x"C0C0C0B0F9F8F9F8",
 31718 => x"C0C0C0B0F9F8F980",
 31719 => x"C0C0C0B0F9F8F990",
 31720 => x"C0C0C0B0F9F8A4C0",
 31721 => x"C0C0C0B0F9F8A4F9",
 31722 => x"C0C0C0B0F9F8A4A4",
 31723 => x"C0C0C0B0F9F8A4B0",
 31724 => x"C0C0C0B0F9F8A499",
 31725 => x"C0C0C0B0F9F8A492",
 31726 => x"C0C0C0B0F9F8A482",
 31727 => x"C0C0C0B0F9F8A4F8",
 31728 => x"C0C0C0B0F9F8A480",
 31729 => x"C0C0C0B0F9F8A490",
 31730 => x"C0C0C0B0F9F8B0C0",
 31731 => x"C0C0C0B0F9F8B0F9",
 31732 => x"C0C0C0B0F9F8B0A4",
 31733 => x"C0C0C0B0F9F8B0B0",
 31734 => x"C0C0C0B0F9F8B099",
 31735 => x"C0C0C0B0F9F8B092",
 31736 => x"C0C0C0B0F9F8B082",
 31737 => x"C0C0C0B0F9F8B0F8",
 31738 => x"C0C0C0B0F9F8B080",
 31739 => x"C0C0C0B0F9F8B090",
 31740 => x"C0C0C0B0F9F899C0",
 31741 => x"C0C0C0B0F9F899F9",
 31742 => x"C0C0C0B0F9F899A4",
 31743 => x"C0C0C0B0F9F899B0",
 31744 => x"C0C0C0B0F9F89999",
 31745 => x"C0C0C0B0F9F89992",
 31746 => x"C0C0C0B0F9F89982",
 31747 => x"C0C0C0B0F9F899F8",
 31748 => x"C0C0C0B0F9F89980",
 31749 => x"C0C0C0B0F9F89990",
 31750 => x"C0C0C0B0F9F892C0",
 31751 => x"C0C0C0B0F9F892F9",
 31752 => x"C0C0C0B0F9F892A4",
 31753 => x"C0C0C0B0F9F892B0",
 31754 => x"C0C0C0B0F9F89299",
 31755 => x"C0C0C0B0F9F89292",
 31756 => x"C0C0C0B0F9F89282",
 31757 => x"C0C0C0B0F9F892F8",
 31758 => x"C0C0C0B0F9F89280",
 31759 => x"C0C0C0B0F9F89290",
 31760 => x"C0C0C0B0F9F882C0",
 31761 => x"C0C0C0B0F9F882F9",
 31762 => x"C0C0C0B0F9F882A4",
 31763 => x"C0C0C0B0F9F882B0",
 31764 => x"C0C0C0B0F9F88299",
 31765 => x"C0C0C0B0F9F88292",
 31766 => x"C0C0C0B0F9F88282",
 31767 => x"C0C0C0B0F9F882F8",
 31768 => x"C0C0C0B0F9F88280",
 31769 => x"C0C0C0B0F9F88290",
 31770 => x"C0C0C0B0F9F8F8C0",
 31771 => x"C0C0C0B0F9F8F8F9",
 31772 => x"C0C0C0B0F9F8F8A4",
 31773 => x"C0C0C0B0F9F8F8B0",
 31774 => x"C0C0C0B0F9F8F899",
 31775 => x"C0C0C0B0F9F8F892",
 31776 => x"C0C0C0B0F9F8F882",
 31777 => x"C0C0C0B0F9F8F8F8",
 31778 => x"C0C0C0B0F9F8F880",
 31779 => x"C0C0C0B0F9F8F890",
 31780 => x"C0C0C0B0F9F880C0",
 31781 => x"C0C0C0B0F9F880F9",
 31782 => x"C0C0C0B0F9F880A4",
 31783 => x"C0C0C0B0F9F880B0",
 31784 => x"C0C0C0B0F9F88099",
 31785 => x"C0C0C0B0F9F88092",
 31786 => x"C0C0C0B0F9F88082",
 31787 => x"C0C0C0B0F9F880F8",
 31788 => x"C0C0C0B0F9F88080",
 31789 => x"C0C0C0B0F9F88090",
 31790 => x"C0C0C0B0F9F890C0",
 31791 => x"C0C0C0B0F9F890F9",
 31792 => x"C0C0C0B0F9F890A4",
 31793 => x"C0C0C0B0F9F890B0",
 31794 => x"C0C0C0B0F9F89099",
 31795 => x"C0C0C0B0F9F89092",
 31796 => x"C0C0C0B0F9F89082",
 31797 => x"C0C0C0B0F9F890F8",
 31798 => x"C0C0C0B0F9F89080",
 31799 => x"C0C0C0B0F9F89090",
 31800 => x"C0C0C0B0F980C0C0",
 31801 => x"C0C0C0B0F980C0F9",
 31802 => x"C0C0C0B0F980C0A4",
 31803 => x"C0C0C0B0F980C0B0",
 31804 => x"C0C0C0B0F980C099",
 31805 => x"C0C0C0B0F980C092",
 31806 => x"C0C0C0B0F980C082",
 31807 => x"C0C0C0B0F980C0F8",
 31808 => x"C0C0C0B0F980C080",
 31809 => x"C0C0C0B0F980C090",
 31810 => x"C0C0C0B0F980F9C0",
 31811 => x"C0C0C0B0F980F9F9",
 31812 => x"C0C0C0B0F980F9A4",
 31813 => x"C0C0C0B0F980F9B0",
 31814 => x"C0C0C0B0F980F999",
 31815 => x"C0C0C0B0F980F992",
 31816 => x"C0C0C0B0F980F982",
 31817 => x"C0C0C0B0F980F9F8",
 31818 => x"C0C0C0B0F980F980",
 31819 => x"C0C0C0B0F980F990",
 31820 => x"C0C0C0B0F980A4C0",
 31821 => x"C0C0C0B0F980A4F9",
 31822 => x"C0C0C0B0F980A4A4",
 31823 => x"C0C0C0B0F980A4B0",
 31824 => x"C0C0C0B0F980A499",
 31825 => x"C0C0C0B0F980A492",
 31826 => x"C0C0C0B0F980A482",
 31827 => x"C0C0C0B0F980A4F8",
 31828 => x"C0C0C0B0F980A480",
 31829 => x"C0C0C0B0F980A490",
 31830 => x"C0C0C0B0F980B0C0",
 31831 => x"C0C0C0B0F980B0F9",
 31832 => x"C0C0C0B0F980B0A4",
 31833 => x"C0C0C0B0F980B0B0",
 31834 => x"C0C0C0B0F980B099",
 31835 => x"C0C0C0B0F980B092",
 31836 => x"C0C0C0B0F980B082",
 31837 => x"C0C0C0B0F980B0F8",
 31838 => x"C0C0C0B0F980B080",
 31839 => x"C0C0C0B0F980B090",
 31840 => x"C0C0C0B0F98099C0",
 31841 => x"C0C0C0B0F98099F9",
 31842 => x"C0C0C0B0F98099A4",
 31843 => x"C0C0C0B0F98099B0",
 31844 => x"C0C0C0B0F9809999",
 31845 => x"C0C0C0B0F9809992",
 31846 => x"C0C0C0B0F9809982",
 31847 => x"C0C0C0B0F98099F8",
 31848 => x"C0C0C0B0F9809980",
 31849 => x"C0C0C0B0F9809990",
 31850 => x"C0C0C0B0F98092C0",
 31851 => x"C0C0C0B0F98092F9",
 31852 => x"C0C0C0B0F98092A4",
 31853 => x"C0C0C0B0F98092B0",
 31854 => x"C0C0C0B0F9809299",
 31855 => x"C0C0C0B0F9809292",
 31856 => x"C0C0C0B0F9809282",
 31857 => x"C0C0C0B0F98092F8",
 31858 => x"C0C0C0B0F9809280",
 31859 => x"C0C0C0B0F9809290",
 31860 => x"C0C0C0B0F98082C0",
 31861 => x"C0C0C0B0F98082F9",
 31862 => x"C0C0C0B0F98082A4",
 31863 => x"C0C0C0B0F98082B0",
 31864 => x"C0C0C0B0F9808299",
 31865 => x"C0C0C0B0F9808292",
 31866 => x"C0C0C0B0F9808282",
 31867 => x"C0C0C0B0F98082F8",
 31868 => x"C0C0C0B0F9808280",
 31869 => x"C0C0C0B0F9808290",
 31870 => x"C0C0C0B0F980F8C0",
 31871 => x"C0C0C0B0F980F8F9",
 31872 => x"C0C0C0B0F980F8A4",
 31873 => x"C0C0C0B0F980F8B0",
 31874 => x"C0C0C0B0F980F899",
 31875 => x"C0C0C0B0F980F892",
 31876 => x"C0C0C0B0F980F882",
 31877 => x"C0C0C0B0F980F8F8",
 31878 => x"C0C0C0B0F980F880",
 31879 => x"C0C0C0B0F980F890",
 31880 => x"C0C0C0B0F98080C0",
 31881 => x"C0C0C0B0F98080F9",
 31882 => x"C0C0C0B0F98080A4",
 31883 => x"C0C0C0B0F98080B0",
 31884 => x"C0C0C0B0F9808099",
 31885 => x"C0C0C0B0F9808092",
 31886 => x"C0C0C0B0F9808082",
 31887 => x"C0C0C0B0F98080F8",
 31888 => x"C0C0C0B0F9808080",
 31889 => x"C0C0C0B0F9808090",
 31890 => x"C0C0C0B0F98090C0",
 31891 => x"C0C0C0B0F98090F9",
 31892 => x"C0C0C0B0F98090A4",
 31893 => x"C0C0C0B0F98090B0",
 31894 => x"C0C0C0B0F9809099",
 31895 => x"C0C0C0B0F9809092",
 31896 => x"C0C0C0B0F9809082",
 31897 => x"C0C0C0B0F98090F8",
 31898 => x"C0C0C0B0F9809080",
 31899 => x"C0C0C0B0F9809090",
 31900 => x"C0C0C0B0F990C0C0",
 31901 => x"C0C0C0B0F990C0F9",
 31902 => x"C0C0C0B0F990C0A4",
 31903 => x"C0C0C0B0F990C0B0",
 31904 => x"C0C0C0B0F990C099",
 31905 => x"C0C0C0B0F990C092",
 31906 => x"C0C0C0B0F990C082",
 31907 => x"C0C0C0B0F990C0F8",
 31908 => x"C0C0C0B0F990C080",
 31909 => x"C0C0C0B0F990C090",
 31910 => x"C0C0C0B0F990F9C0",
 31911 => x"C0C0C0B0F990F9F9",
 31912 => x"C0C0C0B0F990F9A4",
 31913 => x"C0C0C0B0F990F9B0",
 31914 => x"C0C0C0B0F990F999",
 31915 => x"C0C0C0B0F990F992",
 31916 => x"C0C0C0B0F990F982",
 31917 => x"C0C0C0B0F990F9F8",
 31918 => x"C0C0C0B0F990F980",
 31919 => x"C0C0C0B0F990F990",
 31920 => x"C0C0C0B0F990A4C0",
 31921 => x"C0C0C0B0F990A4F9",
 31922 => x"C0C0C0B0F990A4A4",
 31923 => x"C0C0C0B0F990A4B0",
 31924 => x"C0C0C0B0F990A499",
 31925 => x"C0C0C0B0F990A492",
 31926 => x"C0C0C0B0F990A482",
 31927 => x"C0C0C0B0F990A4F8",
 31928 => x"C0C0C0B0F990A480",
 31929 => x"C0C0C0B0F990A490",
 31930 => x"C0C0C0B0F990B0C0",
 31931 => x"C0C0C0B0F990B0F9",
 31932 => x"C0C0C0B0F990B0A4",
 31933 => x"C0C0C0B0F990B0B0",
 31934 => x"C0C0C0B0F990B099",
 31935 => x"C0C0C0B0F990B092",
 31936 => x"C0C0C0B0F990B082",
 31937 => x"C0C0C0B0F990B0F8",
 31938 => x"C0C0C0B0F990B080",
 31939 => x"C0C0C0B0F990B090",
 31940 => x"C0C0C0B0F99099C0",
 31941 => x"C0C0C0B0F99099F9",
 31942 => x"C0C0C0B0F99099A4",
 31943 => x"C0C0C0B0F99099B0",
 31944 => x"C0C0C0B0F9909999",
 31945 => x"C0C0C0B0F9909992",
 31946 => x"C0C0C0B0F9909982",
 31947 => x"C0C0C0B0F99099F8",
 31948 => x"C0C0C0B0F9909980",
 31949 => x"C0C0C0B0F9909990",
 31950 => x"C0C0C0B0F99092C0",
 31951 => x"C0C0C0B0F99092F9",
 31952 => x"C0C0C0B0F99092A4",
 31953 => x"C0C0C0B0F99092B0",
 31954 => x"C0C0C0B0F9909299",
 31955 => x"C0C0C0B0F9909292",
 31956 => x"C0C0C0B0F9909282",
 31957 => x"C0C0C0B0F99092F8",
 31958 => x"C0C0C0B0F9909280",
 31959 => x"C0C0C0B0F9909290",
 31960 => x"C0C0C0B0F99082C0",
 31961 => x"C0C0C0B0F99082F9",
 31962 => x"C0C0C0B0F99082A4",
 31963 => x"C0C0C0B0F99082B0",
 31964 => x"C0C0C0B0F9908299",
 31965 => x"C0C0C0B0F9908292",
 31966 => x"C0C0C0B0F9908282",
 31967 => x"C0C0C0B0F99082F8",
 31968 => x"C0C0C0B0F9908280",
 31969 => x"C0C0C0B0F9908290",
 31970 => x"C0C0C0B0F990F8C0",
 31971 => x"C0C0C0B0F990F8F9",
 31972 => x"C0C0C0B0F990F8A4",
 31973 => x"C0C0C0B0F990F8B0",
 31974 => x"C0C0C0B0F990F899",
 31975 => x"C0C0C0B0F990F892",
 31976 => x"C0C0C0B0F990F882",
 31977 => x"C0C0C0B0F990F8F8",
 31978 => x"C0C0C0B0F990F880",
 31979 => x"C0C0C0B0F990F890",
 31980 => x"C0C0C0B0F99080C0",
 31981 => x"C0C0C0B0F99080F9",
 31982 => x"C0C0C0B0F99080A4",
 31983 => x"C0C0C0B0F99080B0",
 31984 => x"C0C0C0B0F9908099",
 31985 => x"C0C0C0B0F9908092",
 31986 => x"C0C0C0B0F9908082",
 31987 => x"C0C0C0B0F99080F8",
 31988 => x"C0C0C0B0F9908080",
 31989 => x"C0C0C0B0F9908090",
 31990 => x"C0C0C0B0F99090C0",
 31991 => x"C0C0C0B0F99090F9",
 31992 => x"C0C0C0B0F99090A4",
 31993 => x"C0C0C0B0F99090B0",
 31994 => x"C0C0C0B0F9909099",
 31995 => x"C0C0C0B0F9909092",
 31996 => x"C0C0C0B0F9909082",
 31997 => x"C0C0C0B0F99090F8",
 31998 => x"C0C0C0B0F9909080",
 31999 => x"C0C0C0B0F9909090",
 32000 => x"C0C0C0B0A4C0C0C0",
 32001 => x"C0C0C0B0A4C0C0F9",
 32002 => x"C0C0C0B0A4C0C0A4",
 32003 => x"C0C0C0B0A4C0C0B0",
 32004 => x"C0C0C0B0A4C0C099",
 32005 => x"C0C0C0B0A4C0C092",
 32006 => x"C0C0C0B0A4C0C082",
 32007 => x"C0C0C0B0A4C0C0F8",
 32008 => x"C0C0C0B0A4C0C080",
 32009 => x"C0C0C0B0A4C0C090",
 32010 => x"C0C0C0B0A4C0F9C0",
 32011 => x"C0C0C0B0A4C0F9F9",
 32012 => x"C0C0C0B0A4C0F9A4",
 32013 => x"C0C0C0B0A4C0F9B0",
 32014 => x"C0C0C0B0A4C0F999",
 32015 => x"C0C0C0B0A4C0F992",
 32016 => x"C0C0C0B0A4C0F982",
 32017 => x"C0C0C0B0A4C0F9F8",
 32018 => x"C0C0C0B0A4C0F980",
 32019 => x"C0C0C0B0A4C0F990",
 32020 => x"C0C0C0B0A4C0A4C0",
 32021 => x"C0C0C0B0A4C0A4F9",
 32022 => x"C0C0C0B0A4C0A4A4",
 32023 => x"C0C0C0B0A4C0A4B0",
 32024 => x"C0C0C0B0A4C0A499",
 32025 => x"C0C0C0B0A4C0A492",
 32026 => x"C0C0C0B0A4C0A482",
 32027 => x"C0C0C0B0A4C0A4F8",
 32028 => x"C0C0C0B0A4C0A480",
 32029 => x"C0C0C0B0A4C0A490",
 32030 => x"C0C0C0B0A4C0B0C0",
 32031 => x"C0C0C0B0A4C0B0F9",
 32032 => x"C0C0C0B0A4C0B0A4",
 32033 => x"C0C0C0B0A4C0B0B0",
 32034 => x"C0C0C0B0A4C0B099",
 32035 => x"C0C0C0B0A4C0B092",
 32036 => x"C0C0C0B0A4C0B082",
 32037 => x"C0C0C0B0A4C0B0F8",
 32038 => x"C0C0C0B0A4C0B080",
 32039 => x"C0C0C0B0A4C0B090",
 32040 => x"C0C0C0B0A4C099C0",
 32041 => x"C0C0C0B0A4C099F9",
 32042 => x"C0C0C0B0A4C099A4",
 32043 => x"C0C0C0B0A4C099B0",
 32044 => x"C0C0C0B0A4C09999",
 32045 => x"C0C0C0B0A4C09992",
 32046 => x"C0C0C0B0A4C09982",
 32047 => x"C0C0C0B0A4C099F8",
 32048 => x"C0C0C0B0A4C09980",
 32049 => x"C0C0C0B0A4C09990",
 32050 => x"C0C0C0B0A4C092C0",
 32051 => x"C0C0C0B0A4C092F9",
 32052 => x"C0C0C0B0A4C092A4",
 32053 => x"C0C0C0B0A4C092B0",
 32054 => x"C0C0C0B0A4C09299",
 32055 => x"C0C0C0B0A4C09292",
 32056 => x"C0C0C0B0A4C09282",
 32057 => x"C0C0C0B0A4C092F8",
 32058 => x"C0C0C0B0A4C09280",
 32059 => x"C0C0C0B0A4C09290",
 32060 => x"C0C0C0B0A4C082C0",
 32061 => x"C0C0C0B0A4C082F9",
 32062 => x"C0C0C0B0A4C082A4",
 32063 => x"C0C0C0B0A4C082B0",
 32064 => x"C0C0C0B0A4C08299",
 32065 => x"C0C0C0B0A4C08292",
 32066 => x"C0C0C0B0A4C08282",
 32067 => x"C0C0C0B0A4C082F8",
 32068 => x"C0C0C0B0A4C08280",
 32069 => x"C0C0C0B0A4C08290",
 32070 => x"C0C0C0B0A4C0F8C0",
 32071 => x"C0C0C0B0A4C0F8F9",
 32072 => x"C0C0C0B0A4C0F8A4",
 32073 => x"C0C0C0B0A4C0F8B0",
 32074 => x"C0C0C0B0A4C0F899",
 32075 => x"C0C0C0B0A4C0F892",
 32076 => x"C0C0C0B0A4C0F882",
 32077 => x"C0C0C0B0A4C0F8F8",
 32078 => x"C0C0C0B0A4C0F880",
 32079 => x"C0C0C0B0A4C0F890",
 32080 => x"C0C0C0B0A4C080C0",
 32081 => x"C0C0C0B0A4C080F9",
 32082 => x"C0C0C0B0A4C080A4",
 32083 => x"C0C0C0B0A4C080B0",
 32084 => x"C0C0C0B0A4C08099",
 32085 => x"C0C0C0B0A4C08092",
 32086 => x"C0C0C0B0A4C08082",
 32087 => x"C0C0C0B0A4C080F8",
 32088 => x"C0C0C0B0A4C08080",
 32089 => x"C0C0C0B0A4C08090",
 32090 => x"C0C0C0B0A4C090C0",
 32091 => x"C0C0C0B0A4C090F9",
 32092 => x"C0C0C0B0A4C090A4",
 32093 => x"C0C0C0B0A4C090B0",
 32094 => x"C0C0C0B0A4C09099",
 32095 => x"C0C0C0B0A4C09092",
 32096 => x"C0C0C0B0A4C09082",
 32097 => x"C0C0C0B0A4C090F8",
 32098 => x"C0C0C0B0A4C09080",
 32099 => x"C0C0C0B0A4C09090",
 32100 => x"C0C0C0B0A4F9C0C0",
 32101 => x"C0C0C0B0A4F9C0F9",
 32102 => x"C0C0C0B0A4F9C0A4",
 32103 => x"C0C0C0B0A4F9C0B0",
 32104 => x"C0C0C0B0A4F9C099",
 32105 => x"C0C0C0B0A4F9C092",
 32106 => x"C0C0C0B0A4F9C082",
 32107 => x"C0C0C0B0A4F9C0F8",
 32108 => x"C0C0C0B0A4F9C080",
 32109 => x"C0C0C0B0A4F9C090",
 32110 => x"C0C0C0B0A4F9F9C0",
 32111 => x"C0C0C0B0A4F9F9F9",
 32112 => x"C0C0C0B0A4F9F9A4",
 32113 => x"C0C0C0B0A4F9F9B0",
 32114 => x"C0C0C0B0A4F9F999",
 32115 => x"C0C0C0B0A4F9F992",
 32116 => x"C0C0C0B0A4F9F982",
 32117 => x"C0C0C0B0A4F9F9F8",
 32118 => x"C0C0C0B0A4F9F980",
 32119 => x"C0C0C0B0A4F9F990",
 32120 => x"C0C0C0B0A4F9A4C0",
 32121 => x"C0C0C0B0A4F9A4F9",
 32122 => x"C0C0C0B0A4F9A4A4",
 32123 => x"C0C0C0B0A4F9A4B0",
 32124 => x"C0C0C0B0A4F9A499",
 32125 => x"C0C0C0B0A4F9A492",
 32126 => x"C0C0C0B0A4F9A482",
 32127 => x"C0C0C0B0A4F9A4F8",
 32128 => x"C0C0C0B0A4F9A480",
 32129 => x"C0C0C0B0A4F9A490",
 32130 => x"C0C0C0B0A4F9B0C0",
 32131 => x"C0C0C0B0A4F9B0F9",
 32132 => x"C0C0C0B0A4F9B0A4",
 32133 => x"C0C0C0B0A4F9B0B0",
 32134 => x"C0C0C0B0A4F9B099",
 32135 => x"C0C0C0B0A4F9B092",
 32136 => x"C0C0C0B0A4F9B082",
 32137 => x"C0C0C0B0A4F9B0F8",
 32138 => x"C0C0C0B0A4F9B080",
 32139 => x"C0C0C0B0A4F9B090",
 32140 => x"C0C0C0B0A4F999C0",
 32141 => x"C0C0C0B0A4F999F9",
 32142 => x"C0C0C0B0A4F999A4",
 32143 => x"C0C0C0B0A4F999B0",
 32144 => x"C0C0C0B0A4F99999",
 32145 => x"C0C0C0B0A4F99992",
 32146 => x"C0C0C0B0A4F99982",
 32147 => x"C0C0C0B0A4F999F8",
 32148 => x"C0C0C0B0A4F99980",
 32149 => x"C0C0C0B0A4F99990",
 32150 => x"C0C0C0B0A4F992C0",
 32151 => x"C0C0C0B0A4F992F9",
 32152 => x"C0C0C0B0A4F992A4",
 32153 => x"C0C0C0B0A4F992B0",
 32154 => x"C0C0C0B0A4F99299",
 32155 => x"C0C0C0B0A4F99292",
 32156 => x"C0C0C0B0A4F99282",
 32157 => x"C0C0C0B0A4F992F8",
 32158 => x"C0C0C0B0A4F99280",
 32159 => x"C0C0C0B0A4F99290",
 32160 => x"C0C0C0B0A4F982C0",
 32161 => x"C0C0C0B0A4F982F9",
 32162 => x"C0C0C0B0A4F982A4",
 32163 => x"C0C0C0B0A4F982B0",
 32164 => x"C0C0C0B0A4F98299",
 32165 => x"C0C0C0B0A4F98292",
 32166 => x"C0C0C0B0A4F98282",
 32167 => x"C0C0C0B0A4F982F8",
 32168 => x"C0C0C0B0A4F98280",
 32169 => x"C0C0C0B0A4F98290",
 32170 => x"C0C0C0B0A4F9F8C0",
 32171 => x"C0C0C0B0A4F9F8F9",
 32172 => x"C0C0C0B0A4F9F8A4",
 32173 => x"C0C0C0B0A4F9F8B0",
 32174 => x"C0C0C0B0A4F9F899",
 32175 => x"C0C0C0B0A4F9F892",
 32176 => x"C0C0C0B0A4F9F882",
 32177 => x"C0C0C0B0A4F9F8F8",
 32178 => x"C0C0C0B0A4F9F880",
 32179 => x"C0C0C0B0A4F9F890",
 32180 => x"C0C0C0B0A4F980C0",
 32181 => x"C0C0C0B0A4F980F9",
 32182 => x"C0C0C0B0A4F980A4",
 32183 => x"C0C0C0B0A4F980B0",
 32184 => x"C0C0C0B0A4F98099",
 32185 => x"C0C0C0B0A4F98092",
 32186 => x"C0C0C0B0A4F98082",
 32187 => x"C0C0C0B0A4F980F8",
 32188 => x"C0C0C0B0A4F98080",
 32189 => x"C0C0C0B0A4F98090",
 32190 => x"C0C0C0B0A4F990C0",
 32191 => x"C0C0C0B0A4F990F9",
 32192 => x"C0C0C0B0A4F990A4",
 32193 => x"C0C0C0B0A4F990B0",
 32194 => x"C0C0C0B0A4F99099",
 32195 => x"C0C0C0B0A4F99092",
 32196 => x"C0C0C0B0A4F99082",
 32197 => x"C0C0C0B0A4F990F8",
 32198 => x"C0C0C0B0A4F99080",
 32199 => x"C0C0C0B0A4F99090",
 32200 => x"C0C0C0B0A4A4C0C0",
 32201 => x"C0C0C0B0A4A4C0F9",
 32202 => x"C0C0C0B0A4A4C0A4",
 32203 => x"C0C0C0B0A4A4C0B0",
 32204 => x"C0C0C0B0A4A4C099",
 32205 => x"C0C0C0B0A4A4C092",
 32206 => x"C0C0C0B0A4A4C082",
 32207 => x"C0C0C0B0A4A4C0F8",
 32208 => x"C0C0C0B0A4A4C080",
 32209 => x"C0C0C0B0A4A4C090",
 32210 => x"C0C0C0B0A4A4F9C0",
 32211 => x"C0C0C0B0A4A4F9F9",
 32212 => x"C0C0C0B0A4A4F9A4",
 32213 => x"C0C0C0B0A4A4F9B0",
 32214 => x"C0C0C0B0A4A4F999",
 32215 => x"C0C0C0B0A4A4F992",
 32216 => x"C0C0C0B0A4A4F982",
 32217 => x"C0C0C0B0A4A4F9F8",
 32218 => x"C0C0C0B0A4A4F980",
 32219 => x"C0C0C0B0A4A4F990",
 32220 => x"C0C0C0B0A4A4A4C0",
 32221 => x"C0C0C0B0A4A4A4F9",
 32222 => x"C0C0C0B0A4A4A4A4",
 32223 => x"C0C0C0B0A4A4A4B0",
 32224 => x"C0C0C0B0A4A4A499",
 32225 => x"C0C0C0B0A4A4A492",
 32226 => x"C0C0C0B0A4A4A482",
 32227 => x"C0C0C0B0A4A4A4F8",
 32228 => x"C0C0C0B0A4A4A480",
 32229 => x"C0C0C0B0A4A4A490",
 32230 => x"C0C0C0B0A4A4B0C0",
 32231 => x"C0C0C0B0A4A4B0F9",
 32232 => x"C0C0C0B0A4A4B0A4",
 32233 => x"C0C0C0B0A4A4B0B0",
 32234 => x"C0C0C0B0A4A4B099",
 32235 => x"C0C0C0B0A4A4B092",
 32236 => x"C0C0C0B0A4A4B082",
 32237 => x"C0C0C0B0A4A4B0F8",
 32238 => x"C0C0C0B0A4A4B080",
 32239 => x"C0C0C0B0A4A4B090",
 32240 => x"C0C0C0B0A4A499C0",
 32241 => x"C0C0C0B0A4A499F9",
 32242 => x"C0C0C0B0A4A499A4",
 32243 => x"C0C0C0B0A4A499B0",
 32244 => x"C0C0C0B0A4A49999",
 32245 => x"C0C0C0B0A4A49992",
 32246 => x"C0C0C0B0A4A49982",
 32247 => x"C0C0C0B0A4A499F8",
 32248 => x"C0C0C0B0A4A49980",
 32249 => x"C0C0C0B0A4A49990",
 32250 => x"C0C0C0B0A4A492C0",
 32251 => x"C0C0C0B0A4A492F9",
 32252 => x"C0C0C0B0A4A492A4",
 32253 => x"C0C0C0B0A4A492B0",
 32254 => x"C0C0C0B0A4A49299",
 32255 => x"C0C0C0B0A4A49292",
 32256 => x"C0C0C0B0A4A49282",
 32257 => x"C0C0C0B0A4A492F8",
 32258 => x"C0C0C0B0A4A49280",
 32259 => x"C0C0C0B0A4A49290",
 32260 => x"C0C0C0B0A4A482C0",
 32261 => x"C0C0C0B0A4A482F9",
 32262 => x"C0C0C0B0A4A482A4",
 32263 => x"C0C0C0B0A4A482B0",
 32264 => x"C0C0C0B0A4A48299",
 32265 => x"C0C0C0B0A4A48292",
 32266 => x"C0C0C0B0A4A48282",
 32267 => x"C0C0C0B0A4A482F8",
 32268 => x"C0C0C0B0A4A48280",
 32269 => x"C0C0C0B0A4A48290",
 32270 => x"C0C0C0B0A4A4F8C0",
 32271 => x"C0C0C0B0A4A4F8F9",
 32272 => x"C0C0C0B0A4A4F8A4",
 32273 => x"C0C0C0B0A4A4F8B0",
 32274 => x"C0C0C0B0A4A4F899",
 32275 => x"C0C0C0B0A4A4F892",
 32276 => x"C0C0C0B0A4A4F882",
 32277 => x"C0C0C0B0A4A4F8F8",
 32278 => x"C0C0C0B0A4A4F880",
 32279 => x"C0C0C0B0A4A4F890",
 32280 => x"C0C0C0B0A4A480C0",
 32281 => x"C0C0C0B0A4A480F9",
 32282 => x"C0C0C0B0A4A480A4",
 32283 => x"C0C0C0B0A4A480B0",
 32284 => x"C0C0C0B0A4A48099",
 32285 => x"C0C0C0B0A4A48092",
 32286 => x"C0C0C0B0A4A48082",
 32287 => x"C0C0C0B0A4A480F8",
 32288 => x"C0C0C0B0A4A48080",
 32289 => x"C0C0C0B0A4A48090",
 32290 => x"C0C0C0B0A4A490C0",
 32291 => x"C0C0C0B0A4A490F9",
 32292 => x"C0C0C0B0A4A490A4",
 32293 => x"C0C0C0B0A4A490B0",
 32294 => x"C0C0C0B0A4A49099",
 32295 => x"C0C0C0B0A4A49092",
 32296 => x"C0C0C0B0A4A49082",
 32297 => x"C0C0C0B0A4A490F8",
 32298 => x"C0C0C0B0A4A49080",
 32299 => x"C0C0C0B0A4A49090",
 32300 => x"C0C0C0B0A4B0C0C0",
 32301 => x"C0C0C0B0A4B0C0F9",
 32302 => x"C0C0C0B0A4B0C0A4",
 32303 => x"C0C0C0B0A4B0C0B0",
 32304 => x"C0C0C0B0A4B0C099",
 32305 => x"C0C0C0B0A4B0C092",
 32306 => x"C0C0C0B0A4B0C082",
 32307 => x"C0C0C0B0A4B0C0F8",
 32308 => x"C0C0C0B0A4B0C080",
 32309 => x"C0C0C0B0A4B0C090",
 32310 => x"C0C0C0B0A4B0F9C0",
 32311 => x"C0C0C0B0A4B0F9F9",
 32312 => x"C0C0C0B0A4B0F9A4",
 32313 => x"C0C0C0B0A4B0F9B0",
 32314 => x"C0C0C0B0A4B0F999",
 32315 => x"C0C0C0B0A4B0F992",
 32316 => x"C0C0C0B0A4B0F982",
 32317 => x"C0C0C0B0A4B0F9F8",
 32318 => x"C0C0C0B0A4B0F980",
 32319 => x"C0C0C0B0A4B0F990",
 32320 => x"C0C0C0B0A4B0A4C0",
 32321 => x"C0C0C0B0A4B0A4F9",
 32322 => x"C0C0C0B0A4B0A4A4",
 32323 => x"C0C0C0B0A4B0A4B0",
 32324 => x"C0C0C0B0A4B0A499",
 32325 => x"C0C0C0B0A4B0A492",
 32326 => x"C0C0C0B0A4B0A482",
 32327 => x"C0C0C0B0A4B0A4F8",
 32328 => x"C0C0C0B0A4B0A480",
 32329 => x"C0C0C0B0A4B0A490",
 32330 => x"C0C0C0B0A4B0B0C0",
 32331 => x"C0C0C0B0A4B0B0F9",
 32332 => x"C0C0C0B0A4B0B0A4",
 32333 => x"C0C0C0B0A4B0B0B0",
 32334 => x"C0C0C0B0A4B0B099",
 32335 => x"C0C0C0B0A4B0B092",
 32336 => x"C0C0C0B0A4B0B082",
 32337 => x"C0C0C0B0A4B0B0F8",
 32338 => x"C0C0C0B0A4B0B080",
 32339 => x"C0C0C0B0A4B0B090",
 32340 => x"C0C0C0B0A4B099C0",
 32341 => x"C0C0C0B0A4B099F9",
 32342 => x"C0C0C0B0A4B099A4",
 32343 => x"C0C0C0B0A4B099B0",
 32344 => x"C0C0C0B0A4B09999",
 32345 => x"C0C0C0B0A4B09992",
 32346 => x"C0C0C0B0A4B09982",
 32347 => x"C0C0C0B0A4B099F8",
 32348 => x"C0C0C0B0A4B09980",
 32349 => x"C0C0C0B0A4B09990",
 32350 => x"C0C0C0B0A4B092C0",
 32351 => x"C0C0C0B0A4B092F9",
 32352 => x"C0C0C0B0A4B092A4",
 32353 => x"C0C0C0B0A4B092B0",
 32354 => x"C0C0C0B0A4B09299",
 32355 => x"C0C0C0B0A4B09292",
 32356 => x"C0C0C0B0A4B09282",
 32357 => x"C0C0C0B0A4B092F8",
 32358 => x"C0C0C0B0A4B09280",
 32359 => x"C0C0C0B0A4B09290",
 32360 => x"C0C0C0B0A4B082C0",
 32361 => x"C0C0C0B0A4B082F9",
 32362 => x"C0C0C0B0A4B082A4",
 32363 => x"C0C0C0B0A4B082B0",
 32364 => x"C0C0C0B0A4B08299",
 32365 => x"C0C0C0B0A4B08292",
 32366 => x"C0C0C0B0A4B08282",
 32367 => x"C0C0C0B0A4B082F8",
 32368 => x"C0C0C0B0A4B08280",
 32369 => x"C0C0C0B0A4B08290",
 32370 => x"C0C0C0B0A4B0F8C0",
 32371 => x"C0C0C0B0A4B0F8F9",
 32372 => x"C0C0C0B0A4B0F8A4",
 32373 => x"C0C0C0B0A4B0F8B0",
 32374 => x"C0C0C0B0A4B0F899",
 32375 => x"C0C0C0B0A4B0F892",
 32376 => x"C0C0C0B0A4B0F882",
 32377 => x"C0C0C0B0A4B0F8F8",
 32378 => x"C0C0C0B0A4B0F880",
 32379 => x"C0C0C0B0A4B0F890",
 32380 => x"C0C0C0B0A4B080C0",
 32381 => x"C0C0C0B0A4B080F9",
 32382 => x"C0C0C0B0A4B080A4",
 32383 => x"C0C0C0B0A4B080B0",
 32384 => x"C0C0C0B0A4B08099",
 32385 => x"C0C0C0B0A4B08092",
 32386 => x"C0C0C0B0A4B08082",
 32387 => x"C0C0C0B0A4B080F8",
 32388 => x"C0C0C0B0A4B08080",
 32389 => x"C0C0C0B0A4B08090",
 32390 => x"C0C0C0B0A4B090C0",
 32391 => x"C0C0C0B0A4B090F9",
 32392 => x"C0C0C0B0A4B090A4",
 32393 => x"C0C0C0B0A4B090B0",
 32394 => x"C0C0C0B0A4B09099",
 32395 => x"C0C0C0B0A4B09092",
 32396 => x"C0C0C0B0A4B09082",
 32397 => x"C0C0C0B0A4B090F8",
 32398 => x"C0C0C0B0A4B09080",
 32399 => x"C0C0C0B0A4B09090",
 32400 => x"C0C0C0B0A499C0C0",
 32401 => x"C0C0C0B0A499C0F9",
 32402 => x"C0C0C0B0A499C0A4",
 32403 => x"C0C0C0B0A499C0B0",
 32404 => x"C0C0C0B0A499C099",
 32405 => x"C0C0C0B0A499C092",
 32406 => x"C0C0C0B0A499C082",
 32407 => x"C0C0C0B0A499C0F8",
 32408 => x"C0C0C0B0A499C080",
 32409 => x"C0C0C0B0A499C090",
 32410 => x"C0C0C0B0A499F9C0",
 32411 => x"C0C0C0B0A499F9F9",
 32412 => x"C0C0C0B0A499F9A4",
 32413 => x"C0C0C0B0A499F9B0",
 32414 => x"C0C0C0B0A499F999",
 32415 => x"C0C0C0B0A499F992",
 32416 => x"C0C0C0B0A499F982",
 32417 => x"C0C0C0B0A499F9F8",
 32418 => x"C0C0C0B0A499F980",
 32419 => x"C0C0C0B0A499F990",
 32420 => x"C0C0C0B0A499A4C0",
 32421 => x"C0C0C0B0A499A4F9",
 32422 => x"C0C0C0B0A499A4A4",
 32423 => x"C0C0C0B0A499A4B0",
 32424 => x"C0C0C0B0A499A499",
 32425 => x"C0C0C0B0A499A492",
 32426 => x"C0C0C0B0A499A482",
 32427 => x"C0C0C0B0A499A4F8",
 32428 => x"C0C0C0B0A499A480",
 32429 => x"C0C0C0B0A499A490",
 32430 => x"C0C0C0B0A499B0C0",
 32431 => x"C0C0C0B0A499B0F9",
 32432 => x"C0C0C0B0A499B0A4",
 32433 => x"C0C0C0B0A499B0B0",
 32434 => x"C0C0C0B0A499B099",
 32435 => x"C0C0C0B0A499B092",
 32436 => x"C0C0C0B0A499B082",
 32437 => x"C0C0C0B0A499B0F8",
 32438 => x"C0C0C0B0A499B080",
 32439 => x"C0C0C0B0A499B090",
 32440 => x"C0C0C0B0A49999C0",
 32441 => x"C0C0C0B0A49999F9",
 32442 => x"C0C0C0B0A49999A4",
 32443 => x"C0C0C0B0A49999B0",
 32444 => x"C0C0C0B0A4999999",
 32445 => x"C0C0C0B0A4999992",
 32446 => x"C0C0C0B0A4999982",
 32447 => x"C0C0C0B0A49999F8",
 32448 => x"C0C0C0B0A4999980",
 32449 => x"C0C0C0B0A4999990",
 32450 => x"C0C0C0B0A49992C0",
 32451 => x"C0C0C0B0A49992F9",
 32452 => x"C0C0C0B0A49992A4",
 32453 => x"C0C0C0B0A49992B0",
 32454 => x"C0C0C0B0A4999299",
 32455 => x"C0C0C0B0A4999292",
 32456 => x"C0C0C0B0A4999282",
 32457 => x"C0C0C0B0A49992F8",
 32458 => x"C0C0C0B0A4999280",
 32459 => x"C0C0C0B0A4999290",
 32460 => x"C0C0C0B0A49982C0",
 32461 => x"C0C0C0B0A49982F9",
 32462 => x"C0C0C0B0A49982A4",
 32463 => x"C0C0C0B0A49982B0",
 32464 => x"C0C0C0B0A4998299",
 32465 => x"C0C0C0B0A4998292",
 32466 => x"C0C0C0B0A4998282",
 32467 => x"C0C0C0B0A49982F8",
 32468 => x"C0C0C0B0A4998280",
 32469 => x"C0C0C0B0A4998290",
 32470 => x"C0C0C0B0A499F8C0",
 32471 => x"C0C0C0B0A499F8F9",
 32472 => x"C0C0C0B0A499F8A4",
 32473 => x"C0C0C0B0A499F8B0",
 32474 => x"C0C0C0B0A499F899",
 32475 => x"C0C0C0B0A499F892",
 32476 => x"C0C0C0B0A499F882",
 32477 => x"C0C0C0B0A499F8F8",
 32478 => x"C0C0C0B0A499F880",
 32479 => x"C0C0C0B0A499F890",
 32480 => x"C0C0C0B0A49980C0",
 32481 => x"C0C0C0B0A49980F9",
 32482 => x"C0C0C0B0A49980A4",
 32483 => x"C0C0C0B0A49980B0",
 32484 => x"C0C0C0B0A4998099",
 32485 => x"C0C0C0B0A4998092",
 32486 => x"C0C0C0B0A4998082",
 32487 => x"C0C0C0B0A49980F8",
 32488 => x"C0C0C0B0A4998080",
 32489 => x"C0C0C0B0A4998090",
 32490 => x"C0C0C0B0A49990C0",
 32491 => x"C0C0C0B0A49990F9",
 32492 => x"C0C0C0B0A49990A4",
 32493 => x"C0C0C0B0A49990B0",
 32494 => x"C0C0C0B0A4999099",
 32495 => x"C0C0C0B0A4999092",
 32496 => x"C0C0C0B0A4999082",
 32497 => x"C0C0C0B0A49990F8",
 32498 => x"C0C0C0B0A4999080",
 32499 => x"C0C0C0B0A4999090",
 32500 => x"C0C0C0B0A492C0C0",
 32501 => x"C0C0C0B0A492C0F9",
 32502 => x"C0C0C0B0A492C0A4",
 32503 => x"C0C0C0B0A492C0B0",
 32504 => x"C0C0C0B0A492C099",
 32505 => x"C0C0C0B0A492C092",
 32506 => x"C0C0C0B0A492C082",
 32507 => x"C0C0C0B0A492C0F8",
 32508 => x"C0C0C0B0A492C080",
 32509 => x"C0C0C0B0A492C090",
 32510 => x"C0C0C0B0A492F9C0",
 32511 => x"C0C0C0B0A492F9F9",
 32512 => x"C0C0C0B0A492F9A4",
 32513 => x"C0C0C0B0A492F9B0",
 32514 => x"C0C0C0B0A492F999",
 32515 => x"C0C0C0B0A492F992",
 32516 => x"C0C0C0B0A492F982",
 32517 => x"C0C0C0B0A492F9F8",
 32518 => x"C0C0C0B0A492F980",
 32519 => x"C0C0C0B0A492F990",
 32520 => x"C0C0C0B0A492A4C0",
 32521 => x"C0C0C0B0A492A4F9",
 32522 => x"C0C0C0B0A492A4A4",
 32523 => x"C0C0C0B0A492A4B0",
 32524 => x"C0C0C0B0A492A499",
 32525 => x"C0C0C0B0A492A492",
 32526 => x"C0C0C0B0A492A482",
 32527 => x"C0C0C0B0A492A4F8",
 32528 => x"C0C0C0B0A492A480",
 32529 => x"C0C0C0B0A492A490",
 32530 => x"C0C0C0B0A492B0C0",
 32531 => x"C0C0C0B0A492B0F9",
 32532 => x"C0C0C0B0A492B0A4",
 32533 => x"C0C0C0B0A492B0B0",
 32534 => x"C0C0C0B0A492B099",
 32535 => x"C0C0C0B0A492B092",
 32536 => x"C0C0C0B0A492B082",
 32537 => x"C0C0C0B0A492B0F8",
 32538 => x"C0C0C0B0A492B080",
 32539 => x"C0C0C0B0A492B090",
 32540 => x"C0C0C0B0A49299C0",
 32541 => x"C0C0C0B0A49299F9",
 32542 => x"C0C0C0B0A49299A4",
 32543 => x"C0C0C0B0A49299B0",
 32544 => x"C0C0C0B0A4929999",
 32545 => x"C0C0C0B0A4929992",
 32546 => x"C0C0C0B0A4929982",
 32547 => x"C0C0C0B0A49299F8",
 32548 => x"C0C0C0B0A4929980",
 32549 => x"C0C0C0B0A4929990",
 32550 => x"C0C0C0B0A49292C0",
 32551 => x"C0C0C0B0A49292F9",
 32552 => x"C0C0C0B0A49292A4",
 32553 => x"C0C0C0B0A49292B0",
 32554 => x"C0C0C0B0A4929299",
 32555 => x"C0C0C0B0A4929292",
 32556 => x"C0C0C0B0A4929282",
 32557 => x"C0C0C0B0A49292F8",
 32558 => x"C0C0C0B0A4929280",
 32559 => x"C0C0C0B0A4929290",
 32560 => x"C0C0C0B0A49282C0",
 32561 => x"C0C0C0B0A49282F9",
 32562 => x"C0C0C0B0A49282A4",
 32563 => x"C0C0C0B0A49282B0",
 32564 => x"C0C0C0B0A4928299",
 32565 => x"C0C0C0B0A4928292",
 32566 => x"C0C0C0B0A4928282",
 32567 => x"C0C0C0B0A49282F8",
 32568 => x"C0C0C0B0A4928280",
 32569 => x"C0C0C0B0A4928290",
 32570 => x"C0C0C0B0A492F8C0",
 32571 => x"C0C0C0B0A492F8F9",
 32572 => x"C0C0C0B0A492F8A4",
 32573 => x"C0C0C0B0A492F8B0",
 32574 => x"C0C0C0B0A492F899",
 32575 => x"C0C0C0B0A492F892",
 32576 => x"C0C0C0B0A492F882",
 32577 => x"C0C0C0B0A492F8F8",
 32578 => x"C0C0C0B0A492F880",
 32579 => x"C0C0C0B0A492F890",
 32580 => x"C0C0C0B0A49280C0",
 32581 => x"C0C0C0B0A49280F9",
 32582 => x"C0C0C0B0A49280A4",
 32583 => x"C0C0C0B0A49280B0",
 32584 => x"C0C0C0B0A4928099",
 32585 => x"C0C0C0B0A4928092",
 32586 => x"C0C0C0B0A4928082",
 32587 => x"C0C0C0B0A49280F8",
 32588 => x"C0C0C0B0A4928080",
 32589 => x"C0C0C0B0A4928090",
 32590 => x"C0C0C0B0A49290C0",
 32591 => x"C0C0C0B0A49290F9",
 32592 => x"C0C0C0B0A49290A4",
 32593 => x"C0C0C0B0A49290B0",
 32594 => x"C0C0C0B0A4929099",
 32595 => x"C0C0C0B0A4929092",
 32596 => x"C0C0C0B0A4929082",
 32597 => x"C0C0C0B0A49290F8",
 32598 => x"C0C0C0B0A4929080",
 32599 => x"C0C0C0B0A4929090",
 32600 => x"C0C0C0B0A482C0C0",
 32601 => x"C0C0C0B0A482C0F9",
 32602 => x"C0C0C0B0A482C0A4",
 32603 => x"C0C0C0B0A482C0B0",
 32604 => x"C0C0C0B0A482C099",
 32605 => x"C0C0C0B0A482C092",
 32606 => x"C0C0C0B0A482C082",
 32607 => x"C0C0C0B0A482C0F8",
 32608 => x"C0C0C0B0A482C080",
 32609 => x"C0C0C0B0A482C090",
 32610 => x"C0C0C0B0A482F9C0",
 32611 => x"C0C0C0B0A482F9F9",
 32612 => x"C0C0C0B0A482F9A4",
 32613 => x"C0C0C0B0A482F9B0",
 32614 => x"C0C0C0B0A482F999",
 32615 => x"C0C0C0B0A482F992",
 32616 => x"C0C0C0B0A482F982",
 32617 => x"C0C0C0B0A482F9F8",
 32618 => x"C0C0C0B0A482F980",
 32619 => x"C0C0C0B0A482F990",
 32620 => x"C0C0C0B0A482A4C0",
 32621 => x"C0C0C0B0A482A4F9",
 32622 => x"C0C0C0B0A482A4A4",
 32623 => x"C0C0C0B0A482A4B0",
 32624 => x"C0C0C0B0A482A499",
 32625 => x"C0C0C0B0A482A492",
 32626 => x"C0C0C0B0A482A482",
 32627 => x"C0C0C0B0A482A4F8",
 32628 => x"C0C0C0B0A482A480",
 32629 => x"C0C0C0B0A482A490",
 32630 => x"C0C0C0B0A482B0C0",
 32631 => x"C0C0C0B0A482B0F9",
 32632 => x"C0C0C0B0A482B0A4",
 32633 => x"C0C0C0B0A482B0B0",
 32634 => x"C0C0C0B0A482B099",
 32635 => x"C0C0C0B0A482B092",
 32636 => x"C0C0C0B0A482B082",
 32637 => x"C0C0C0B0A482B0F8",
 32638 => x"C0C0C0B0A482B080",
 32639 => x"C0C0C0B0A482B090",
 32640 => x"C0C0C0B0A48299C0",
 32641 => x"C0C0C0B0A48299F9",
 32642 => x"C0C0C0B0A48299A4",
 32643 => x"C0C0C0B0A48299B0",
 32644 => x"C0C0C0B0A4829999",
 32645 => x"C0C0C0B0A4829992",
 32646 => x"C0C0C0B0A4829982",
 32647 => x"C0C0C0B0A48299F8",
 32648 => x"C0C0C0B0A4829980",
 32649 => x"C0C0C0B0A4829990",
 32650 => x"C0C0C0B0A48292C0",
 32651 => x"C0C0C0B0A48292F9",
 32652 => x"C0C0C0B0A48292A4",
 32653 => x"C0C0C0B0A48292B0",
 32654 => x"C0C0C0B0A4829299",
 32655 => x"C0C0C0B0A4829292",
 32656 => x"C0C0C0B0A4829282",
 32657 => x"C0C0C0B0A48292F8",
 32658 => x"C0C0C0B0A4829280",
 32659 => x"C0C0C0B0A4829290",
 32660 => x"C0C0C0B0A48282C0",
 32661 => x"C0C0C0B0A48282F9",
 32662 => x"C0C0C0B0A48282A4",
 32663 => x"C0C0C0B0A48282B0",
 32664 => x"C0C0C0B0A4828299",
 32665 => x"C0C0C0B0A4828292",
 32666 => x"C0C0C0B0A4828282",
 32667 => x"C0C0C0B0A48282F8",
 32668 => x"C0C0C0B0A4828280",
 32669 => x"C0C0C0B0A4828290",
 32670 => x"C0C0C0B0A482F8C0",
 32671 => x"C0C0C0B0A482F8F9",
 32672 => x"C0C0C0B0A482F8A4",
 32673 => x"C0C0C0B0A482F8B0",
 32674 => x"C0C0C0B0A482F899",
 32675 => x"C0C0C0B0A482F892",
 32676 => x"C0C0C0B0A482F882",
 32677 => x"C0C0C0B0A482F8F8",
 32678 => x"C0C0C0B0A482F880",
 32679 => x"C0C0C0B0A482F890",
 32680 => x"C0C0C0B0A48280C0",
 32681 => x"C0C0C0B0A48280F9",
 32682 => x"C0C0C0B0A48280A4",
 32683 => x"C0C0C0B0A48280B0",
 32684 => x"C0C0C0B0A4828099",
 32685 => x"C0C0C0B0A4828092",
 32686 => x"C0C0C0B0A4828082",
 32687 => x"C0C0C0B0A48280F8",
 32688 => x"C0C0C0B0A4828080",
 32689 => x"C0C0C0B0A4828090",
 32690 => x"C0C0C0B0A48290C0",
 32691 => x"C0C0C0B0A48290F9",
 32692 => x"C0C0C0B0A48290A4",
 32693 => x"C0C0C0B0A48290B0",
 32694 => x"C0C0C0B0A4829099",
 32695 => x"C0C0C0B0A4829092",
 32696 => x"C0C0C0B0A4829082",
 32697 => x"C0C0C0B0A48290F8",
 32698 => x"C0C0C0B0A4829080",
 32699 => x"C0C0C0B0A4829090",
 32700 => x"C0C0C0B0A4F8C0C0",
 32701 => x"C0C0C0B0A4F8C0F9",
 32702 => x"C0C0C0B0A4F8C0A4",
 32703 => x"C0C0C0B0A4F8C0B0",
 32704 => x"C0C0C0B0A4F8C099",
 32705 => x"C0C0C0B0A4F8C092",
 32706 => x"C0C0C0B0A4F8C082",
 32707 => x"C0C0C0B0A4F8C0F8",
 32708 => x"C0C0C0B0A4F8C080",
 32709 => x"C0C0C0B0A4F8C090",
 32710 => x"C0C0C0B0A4F8F9C0",
 32711 => x"C0C0C0B0A4F8F9F9",
 32712 => x"C0C0C0B0A4F8F9A4",
 32713 => x"C0C0C0B0A4F8F9B0",
 32714 => x"C0C0C0B0A4F8F999",
 32715 => x"C0C0C0B0A4F8F992",
 32716 => x"C0C0C0B0A4F8F982",
 32717 => x"C0C0C0B0A4F8F9F8",
 32718 => x"C0C0C0B0A4F8F980",
 32719 => x"C0C0C0B0A4F8F990",
 32720 => x"C0C0C0B0A4F8A4C0",
 32721 => x"C0C0C0B0A4F8A4F9",
 32722 => x"C0C0C0B0A4F8A4A4",
 32723 => x"C0C0C0B0A4F8A4B0",
 32724 => x"C0C0C0B0A4F8A499",
 32725 => x"C0C0C0B0A4F8A492",
 32726 => x"C0C0C0B0A4F8A482",
 32727 => x"C0C0C0B0A4F8A4F8",
 32728 => x"C0C0C0B0A4F8A480",
 32729 => x"C0C0C0B0A4F8A490",
 32730 => x"C0C0C0B0A4F8B0C0",
 32731 => x"C0C0C0B0A4F8B0F9",
 32732 => x"C0C0C0B0A4F8B0A4",
 32733 => x"C0C0C0B0A4F8B0B0",
 32734 => x"C0C0C0B0A4F8B099",
 32735 => x"C0C0C0B0A4F8B092",
 32736 => x"C0C0C0B0A4F8B082",
 32737 => x"C0C0C0B0A4F8B0F8",
 32738 => x"C0C0C0B0A4F8B080",
 32739 => x"C0C0C0B0A4F8B090",
 32740 => x"C0C0C0B0A4F899C0",
 32741 => x"C0C0C0B0A4F899F9",
 32742 => x"C0C0C0B0A4F899A4",
 32743 => x"C0C0C0B0A4F899B0",
 32744 => x"C0C0C0B0A4F89999",
 32745 => x"C0C0C0B0A4F89992",
 32746 => x"C0C0C0B0A4F89982",
 32747 => x"C0C0C0B0A4F899F8",
 32748 => x"C0C0C0B0A4F89980",
 32749 => x"C0C0C0B0A4F89990",
 32750 => x"C0C0C0B0A4F892C0",
 32751 => x"C0C0C0B0A4F892F9",
 32752 => x"C0C0C0B0A4F892A4",
 32753 => x"C0C0C0B0A4F892B0",
 32754 => x"C0C0C0B0A4F89299",
 32755 => x"C0C0C0B0A4F89292",
 32756 => x"C0C0C0B0A4F89282",
 32757 => x"C0C0C0B0A4F892F8",
 32758 => x"C0C0C0B0A4F89280",
 32759 => x"C0C0C0B0A4F89290",
 32760 => x"C0C0C0B0A4F882C0",
 32761 => x"C0C0C0B0A4F882F9",
 32762 => x"C0C0C0B0A4F882A4",
 32763 => x"C0C0C0B0A4F882B0",
 32764 => x"C0C0C0B0A4F88299",
 32765 => x"C0C0C0B0A4F88292",
 32766 => x"C0C0C0B0A4F88282",
 32767 => x"C0C0C0B0A4F882F8"
); 
begin

outp <= ROM(to_integer(signed(inp)));

end Behavioral;
